module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    compressor_CLA162_64 compressor_CLA162_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
        src32 <= 162'h0;
        src33 <= 162'h0;
        src34 <= 162'h0;
        src35 <= 162'h0;
        src36 <= 162'h0;
        src37 <= 162'h0;
        src38 <= 162'h0;
        src39 <= 162'h0;
        src40 <= 162'h0;
        src41 <= 162'h0;
        src42 <= 162'h0;
        src43 <= 162'h0;
        src44 <= 162'h0;
        src45 <= 162'h0;
        src46 <= 162'h0;
        src47 <= 162'h0;
        src48 <= 162'h0;
        src49 <= 162'h0;
        src50 <= 162'h0;
        src51 <= 162'h0;
        src52 <= 162'h0;
        src53 <= 162'h0;
        src54 <= 162'h0;
        src55 <= 162'h0;
        src56 <= 162'h0;
        src57 <= 162'h0;
        src58 <= 162'h0;
        src59 <= 162'h0;
        src60 <= 162'h0;
        src61 <= 162'h0;
        src62 <= 162'h0;
        src63 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA162_64(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    input [161:0]src32,
    input [161:0]src33,
    input [161:0]src34,
    input [161:0]src35,
    input [161:0]src36,
    input [161:0]src37,
    input [161:0]src38,
    input [161:0]src39,
    input [161:0]src40,
    input [161:0]src41,
    input [161:0]src42,
    input [161:0]src43,
    input [161:0]src44,
    input [161:0]src45,
    input [161:0]src46,
    input [161:0]src47,
    input [161:0]src48,
    input [161:0]src49,
    input [161:0]src50,
    input [161:0]src51,
    input [161:0]src52,
    input [161:0]src53,
    input [161:0]src54,
    input [161:0]src55,
    input [161:0]src56,
    input [161:0]src57,
    input [161:0]src58,
    input [161:0]src59,
    input [161:0]src60,
    input [161:0]src61,
    input [161:0]src62,
    input [161:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [0:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [0:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [0:0] comp_out70;
    wire [0:0] comp_out71;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], 1'h0, comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], 1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], 1'h0, comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], 1'h0, 1'h0, 1'h0, comp_out0[1]}),
        .dst({dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      input wire [161:0] src32,
      input wire [161:0] src33,
      input wire [161:0] src34,
      input wire [161:0] src35,
      input wire [161:0] src36,
      input wire [161:0] src37,
      input wire [161:0] src38,
      input wire [161:0] src39,
      input wire [161:0] src40,
      input wire [161:0] src41,
      input wire [161:0] src42,
      input wire [161:0] src43,
      input wire [161:0] src44,
      input wire [161:0] src45,
      input wire [161:0] src46,
      input wire [161:0] src47,
      input wire [161:0] src48,
      input wire [161:0] src49,
      input wire [161:0] src50,
      input wire [161:0] src51,
      input wire [161:0] src52,
      input wire [161:0] src53,
      input wire [161:0] src54,
      input wire [161:0] src55,
      input wire [161:0] src56,
      input wire [161:0] src57,
      input wire [161:0] src58,
      input wire [161:0] src59,
      input wire [161:0] src60,
      input wire [161:0] src61,
      input wire [161:0] src62,
      input wire [161:0] src63,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [0:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [0:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [0:0] dst70,
      output wire [0:0] dst71);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [161:0] stage0_32;
   wire [161:0] stage0_33;
   wire [161:0] stage0_34;
   wire [161:0] stage0_35;
   wire [161:0] stage0_36;
   wire [161:0] stage0_37;
   wire [161:0] stage0_38;
   wire [161:0] stage0_39;
   wire [161:0] stage0_40;
   wire [161:0] stage0_41;
   wire [161:0] stage0_42;
   wire [161:0] stage0_43;
   wire [161:0] stage0_44;
   wire [161:0] stage0_45;
   wire [161:0] stage0_46;
   wire [161:0] stage0_47;
   wire [161:0] stage0_48;
   wire [161:0] stage0_49;
   wire [161:0] stage0_50;
   wire [161:0] stage0_51;
   wire [161:0] stage0_52;
   wire [161:0] stage0_53;
   wire [161:0] stage0_54;
   wire [161:0] stage0_55;
   wire [161:0] stage0_56;
   wire [161:0] stage0_57;
   wire [161:0] stage0_58;
   wire [161:0] stage0_59;
   wire [161:0] stage0_60;
   wire [161:0] stage0_61;
   wire [161:0] stage0_62;
   wire [161:0] stage0_63;
   wire [33:0] stage1_0;
   wire [46:0] stage1_1;
   wire [54:0] stage1_2;
   wire [83:0] stage1_3;
   wire [82:0] stage1_4;
   wire [114:0] stage1_5;
   wire [57:0] stage1_6;
   wire [70:0] stage1_7;
   wire [80:0] stage1_8;
   wire [57:0] stage1_9;
   wire [94:0] stage1_10;
   wire [80:0] stage1_11;
   wire [66:0] stage1_12;
   wire [86:0] stage1_13;
   wire [61:0] stage1_14;
   wire [97:0] stage1_15;
   wire [67:0] stage1_16;
   wire [113:0] stage1_17;
   wire [62:0] stage1_18;
   wire [70:0] stage1_19;
   wire [67:0] stage1_20;
   wire [70:0] stage1_21;
   wire [66:0] stage1_22;
   wire [142:0] stage1_23;
   wire [82:0] stage1_24;
   wire [84:0] stage1_25;
   wire [71:0] stage1_26;
   wire [73:0] stage1_27;
   wire [76:0] stage1_28;
   wire [80:0] stage1_29;
   wire [106:0] stage1_30;
   wire [96:0] stage1_31;
   wire [86:0] stage1_32;
   wire [89:0] stage1_33;
   wire [55:0] stage1_34;
   wire [59:0] stage1_35;
   wire [82:0] stage1_36;
   wire [127:0] stage1_37;
   wire [65:0] stage1_38;
   wire [67:0] stage1_39;
   wire [81:0] stage1_40;
   wire [73:0] stage1_41;
   wire [95:0] stage1_42;
   wire [137:0] stage1_43;
   wire [45:0] stage1_44;
   wire [92:0] stage1_45;
   wire [63:0] stage1_46;
   wire [57:0] stage1_47;
   wire [71:0] stage1_48;
   wire [86:0] stage1_49;
   wire [57:0] stage1_50;
   wire [93:0] stage1_51;
   wire [76:0] stage1_52;
   wire [65:0] stage1_53;
   wire [57:0] stage1_54;
   wire [97:0] stage1_55;
   wire [79:0] stage1_56;
   wire [71:0] stage1_57;
   wire [73:0] stage1_58;
   wire [79:0] stage1_59;
   wire [66:0] stage1_60;
   wire [90:0] stage1_61;
   wire [86:0] stage1_62;
   wire [62:0] stage1_63;
   wire [44:0] stage1_64;
   wire [23:0] stage1_65;
   wire [9:0] stage2_0;
   wire [18:0] stage2_1;
   wire [37:0] stage2_2;
   wire [22:0] stage2_3;
   wire [47:0] stage2_4;
   wire [35:0] stage2_5;
   wire [28:0] stage2_6;
   wire [40:0] stage2_7;
   wire [60:0] stage2_8;
   wire [25:0] stage2_9;
   wire [40:0] stage2_10;
   wire [38:0] stage2_11;
   wire [30:0] stage2_12;
   wire [44:0] stage2_13;
   wire [73:0] stage2_14;
   wire [36:0] stage2_15;
   wire [46:0] stage2_16;
   wire [39:0] stage2_17;
   wire [42:0] stage2_18;
   wire [50:0] stage2_19;
   wire [57:0] stage2_20;
   wire [39:0] stage2_21;
   wire [30:0] stage2_22;
   wire [46:0] stage2_23;
   wire [45:0] stage2_24;
   wire [36:0] stage2_25;
   wire [52:0] stage2_26;
   wire [49:0] stage2_27;
   wire [34:0] stage2_28;
   wire [49:0] stage2_29;
   wire [49:0] stage2_30;
   wire [38:0] stage2_31;
   wire [55:0] stage2_32;
   wire [27:0] stage2_33;
   wire [34:0] stage2_34;
   wire [44:0] stage2_35;
   wire [36:0] stage2_36;
   wire [41:0] stage2_37;
   wire [32:0] stage2_38;
   wire [33:0] stage2_39;
   wire [40:0] stage2_40;
   wire [55:0] stage2_41;
   wire [61:0] stage2_42;
   wire [51:0] stage2_43;
   wire [65:0] stage2_44;
   wire [25:0] stage2_45;
   wire [32:0] stage2_46;
   wire [45:0] stage2_47;
   wire [23:0] stage2_48;
   wire [36:0] stage2_49;
   wire [40:0] stage2_50;
   wire [24:0] stage2_51;
   wire [33:0] stage2_52;
   wire [50:0] stage2_53;
   wire [27:0] stage2_54;
   wire [37:0] stage2_55;
   wire [52:0] stage2_56;
   wire [29:0] stage2_57;
   wire [32:0] stage2_58;
   wire [80:0] stage2_59;
   wire [21:0] stage2_60;
   wire [66:0] stage2_61;
   wire [34:0] stage2_62;
   wire [37:0] stage2_63;
   wire [45:0] stage2_64;
   wire [12:0] stage2_65;
   wire [9:0] stage2_66;
   wire [1:0] stage2_67;
   wire [7:0] stage3_0;
   wire [13:0] stage3_1;
   wire [10:0] stage3_2;
   wire [13:0] stage3_3;
   wire [13:0] stage3_4;
   wire [17:0] stage3_5;
   wire [19:0] stage3_6;
   wire [16:0] stage3_7;
   wire [16:0] stage3_8;
   wire [20:0] stage3_9;
   wire [14:0] stage3_10;
   wire [17:0] stage3_11;
   wire [23:0] stage3_12;
   wire [19:0] stage3_13;
   wire [35:0] stage3_14;
   wire [36:0] stage3_15;
   wire [21:0] stage3_16;
   wire [16:0] stage3_17;
   wire [22:0] stage3_18;
   wire [26:0] stage3_19;
   wire [22:0] stage3_20;
   wire [24:0] stage3_21;
   wire [26:0] stage3_22;
   wire [11:0] stage3_23;
   wire [25:0] stage3_24;
   wire [21:0] stage3_25;
   wire [15:0] stage3_26;
   wire [18:0] stage3_27;
   wire [19:0] stage3_28;
   wire [23:0] stage3_29;
   wire [25:0] stage3_30;
   wire [20:0] stage3_31;
   wire [34:0] stage3_32;
   wire [14:0] stage3_33;
   wire [22:0] stage3_34;
   wire [25:0] stage3_35;
   wire [16:0] stage3_36;
   wire [11:0] stage3_37;
   wire [13:0] stage3_38;
   wire [23:0] stage3_39;
   wire [23:0] stage3_40;
   wire [24:0] stage3_41;
   wire [25:0] stage3_42;
   wire [20:0] stage3_43;
   wire [30:0] stage3_44;
   wire [17:0] stage3_45;
   wire [16:0] stage3_46;
   wire [23:0] stage3_47;
   wire [15:0] stage3_48;
   wire [13:0] stage3_49;
   wire [31:0] stage3_50;
   wire [13:0] stage3_51;
   wire [23:0] stage3_52;
   wire [15:0] stage3_53;
   wire [15:0] stage3_54;
   wire [17:0] stage3_55;
   wire [30:0] stage3_56;
   wire [12:0] stage3_57;
   wire [32:0] stage3_58;
   wire [27:0] stage3_59;
   wire [14:0] stage3_60;
   wire [24:0] stage3_61;
   wire [20:0] stage3_62;
   wire [17:0] stage3_63;
   wire [28:0] stage3_64;
   wire [13:0] stage3_65;
   wire [8:0] stage3_66;
   wire [4:0] stage3_67;
   wire [1:0] stage3_68;
   wire [3:0] stage4_0;
   wire [3:0] stage4_1;
   wire [6:0] stage4_2;
   wire [4:0] stage4_3;
   wire [8:0] stage4_4;
   wire [8:0] stage4_5;
   wire [13:0] stage4_6;
   wire [7:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [8:0] stage4_10;
   wire [6:0] stage4_11;
   wire [8:0] stage4_12;
   wire [9:0] stage4_13;
   wire [10:0] stage4_14;
   wire [16:0] stage4_15;
   wire [12:0] stage4_16;
   wire [16:0] stage4_17;
   wire [5:0] stage4_18;
   wire [15:0] stage4_19;
   wire [10:0] stage4_20;
   wire [7:0] stage4_21;
   wire [13:0] stage4_22;
   wire [9:0] stage4_23;
   wire [17:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [6:0] stage4_27;
   wire [11:0] stage4_28;
   wire [9:0] stage4_29;
   wire [15:0] stage4_30;
   wire [8:0] stage4_31;
   wire [19:0] stage4_32;
   wire [11:0] stage4_33;
   wire [10:0] stage4_34;
   wire [10:0] stage4_35;
   wire [9:0] stage4_36;
   wire [5:0] stage4_37;
   wire [5:0] stage4_38;
   wire [9:0] stage4_39;
   wire [13:0] stage4_40;
   wire [16:0] stage4_41;
   wire [16:0] stage4_42;
   wire [6:0] stage4_43;
   wire [12:0] stage4_44;
   wire [8:0] stage4_45;
   wire [17:0] stage4_46;
   wire [15:0] stage4_47;
   wire [11:0] stage4_48;
   wire [12:0] stage4_49;
   wire [6:0] stage4_50;
   wire [8:0] stage4_51;
   wire [8:0] stage4_52;
   wire [14:0] stage4_53;
   wire [9:0] stage4_54;
   wire [16:0] stage4_55;
   wire [12:0] stage4_56;
   wire [5:0] stage4_57;
   wire [20:0] stage4_58;
   wire [16:0] stage4_59;
   wire [15:0] stage4_60;
   wire [16:0] stage4_61;
   wire [7:0] stage4_62;
   wire [12:0] stage4_63;
   wire [21:0] stage4_64;
   wire [5:0] stage4_65;
   wire [12:0] stage4_66;
   wire [6:0] stage4_67;
   wire [1:0] stage4_68;
   wire [1:0] stage5_0;
   wire [0:0] stage5_1;
   wire [4:0] stage5_2;
   wire [4:0] stage5_3;
   wire [4:0] stage5_4;
   wire [4:0] stage5_5;
   wire [9:0] stage5_6;
   wire [3:0] stage5_7;
   wire [7:0] stage5_8;
   wire [2:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [10:0] stage5_12;
   wire [5:0] stage5_13;
   wire [7:0] stage5_14;
   wire [7:0] stage5_15;
   wire [8:0] stage5_16;
   wire [4:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [3:0] stage5_20;
   wire [5:0] stage5_21;
   wire [10:0] stage5_22;
   wire [6:0] stage5_23;
   wire [9:0] stage5_24;
   wire [2:0] stage5_25;
   wire [2:0] stage5_26;
   wire [3:0] stage5_27;
   wire [4:0] stage5_28;
   wire [3:0] stage5_29;
   wire [4:0] stage5_30;
   wire [5:0] stage5_31;
   wire [11:0] stage5_32;
   wire [4:0] stage5_33;
   wire [7:0] stage5_34;
   wire [3:0] stage5_35;
   wire [4:0] stage5_36;
   wire [3:0] stage5_37;
   wire [1:0] stage5_38;
   wire [5:0] stage5_39;
   wire [5:0] stage5_40;
   wire [12:0] stage5_41;
   wire [4:0] stage5_42;
   wire [3:0] stage5_43;
   wire [5:0] stage5_44;
   wire [4:0] stage5_45;
   wire [5:0] stage5_46;
   wire [12:0] stage5_47;
   wire [3:0] stage5_48;
   wire [6:0] stage5_49;
   wire [4:0] stage5_50;
   wire [3:0] stage5_51;
   wire [5:0] stage5_52;
   wire [6:0] stage5_53;
   wire [8:0] stage5_54;
   wire [6:0] stage5_55;
   wire [4:0] stage5_56;
   wire [5:0] stage5_57;
   wire [5:0] stage5_58;
   wire [5:0] stage5_59;
   wire [8:0] stage5_60;
   wire [10:0] stage5_61;
   wire [5:0] stage5_62;
   wire [11:0] stage5_63;
   wire [10:0] stage5_64;
   wire [3:0] stage5_65;
   wire [4:0] stage5_66;
   wire [3:0] stage5_67;
   wire [4:0] stage5_68;
   wire [0:0] stage5_69;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [4:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [4:0] stage6_7;
   wire [1:0] stage6_8;
   wire [2:0] stage6_9;
   wire [6:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [1:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [6:0] stage6_17;
   wire [0:0] stage6_18;
   wire [3:0] stage6_19;
   wire [2:0] stage6_20;
   wire [5:0] stage6_21;
   wire [3:0] stage6_22;
   wire [2:0] stage6_23;
   wire [2:0] stage6_24;
   wire [2:0] stage6_25;
   wire [2:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [8:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [1:0] stage6_35;
   wire [6:0] stage6_36;
   wire [4:0] stage6_37;
   wire [0:0] stage6_38;
   wire [1:0] stage6_39;
   wire [1:0] stage6_40;
   wire [3:0] stage6_41;
   wire [7:0] stage6_42;
   wire [1:0] stage6_43;
   wire [1:0] stage6_44;
   wire [2:0] stage6_45;
   wire [1:0] stage6_46;
   wire [4:0] stage6_47;
   wire [5:0] stage6_48;
   wire [2:0] stage6_49;
   wire [3:0] stage6_50;
   wire [1:0] stage6_51;
   wire [3:0] stage6_52;
   wire [4:0] stage6_53;
   wire [2:0] stage6_54;
   wire [2:0] stage6_55;
   wire [4:0] stage6_56;
   wire [1:0] stage6_57;
   wire [1:0] stage6_58;
   wire [2:0] stage6_59;
   wire [4:0] stage6_60;
   wire [2:0] stage6_61;
   wire [3:0] stage6_62;
   wire [3:0] stage6_63;
   wire [3:0] stage6_64;
   wire [3:0] stage6_65;
   wire [2:0] stage6_66;
   wire [5:0] stage6_67;
   wire [5:0] stage6_68;
   wire [0:0] stage6_69;
   wire [1:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [0:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [1:0] stage7_25;
   wire [0:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [1:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage7_41;
   wire [1:0] stage7_42;
   wire [1:0] stage7_43;
   wire [1:0] stage7_44;
   wire [1:0] stage7_45;
   wire [1:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [1:0] stage7_49;
   wire [1:0] stage7_50;
   wire [1:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [1:0] stage7_54;
   wire [1:0] stage7_55;
   wire [1:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [1:0] stage7_59;
   wire [1:0] stage7_60;
   wire [0:0] stage7_61;
   wire [1:0] stage7_62;
   wire [1:0] stage7_63;
   wire [1:0] stage7_64;
   wire [1:0] stage7_65;
   wire [1:0] stage7_66;
   wire [1:0] stage7_67;
   wire [1:0] stage7_68;
   wire [1:0] stage7_69;
   wire [0:0] stage7_70;
   wire [0:0] stage7_71;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;
   assign dst40 = stage7_40;
   assign dst41 = stage7_41;
   assign dst42 = stage7_42;
   assign dst43 = stage7_43;
   assign dst44 = stage7_44;
   assign dst45 = stage7_45;
   assign dst46 = stage7_46;
   assign dst47 = stage7_47;
   assign dst48 = stage7_48;
   assign dst49 = stage7_49;
   assign dst50 = stage7_50;
   assign dst51 = stage7_51;
   assign dst52 = stage7_52;
   assign dst53 = stage7_53;
   assign dst54 = stage7_54;
   assign dst55 = stage7_55;
   assign dst56 = stage7_56;
   assign dst57 = stage7_57;
   assign dst58 = stage7_58;
   assign dst59 = stage7_59;
   assign dst60 = stage7_60;
   assign dst61 = stage7_61;
   assign dst62 = stage7_62;
   assign dst63 = stage7_63;
   assign dst64 = stage7_64;
   assign dst65 = stage7_65;
   assign dst66 = stage7_66;
   assign dst67 = stage7_67;
   assign dst68 = stage7_68;
   assign dst69 = stage7_69;
   assign dst70 = stage7_70;
   assign dst71 = stage7_71;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7]},
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[1]},
      {stage0_3[2]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[2]},
      {stage0_3[3]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[3]},
      {stage0_3[4]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[4]},
      {stage0_3[5]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[5]},
      {stage0_3[6]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[6]},
      {stage0_3[7]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[7]},
      {stage0_3[8]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[8]},
      {stage0_3[9]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[9]},
      {stage0_3[10]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[10]},
      {stage0_3[11]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[11]},
      {stage0_3[12]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[12]},
      {stage0_3[13]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[13]},
      {stage0_3[14]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc207_4 gpc14 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[14], stage0_2[15]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[14],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[15],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[16],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc615_5 gpc31 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[81]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc615_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[82]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc615_5 gpc33 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_1[83]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[0],stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[1],stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[2],stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[3],stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[4],stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[5],stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[6],stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[7],stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[8],stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[9],stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[10],stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[11],stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[12],stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage0_3[93]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[13],stage1_4[46],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_3[94]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[14],stage1_4[47],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage0_3[95]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[15],stage1_4[48],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage0_3[96]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[16],stage1_4[49],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154]},
      {stage0_3[97]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[17],stage1_4[50],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159]},
      {stage0_3[98]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[18],stage1_4[51],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage0_4[36]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[6],stage1_5[19],stage1_4[52],stage1_3[53]}
   );
   gpc615_5 gpc54 (
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage0_4[37]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[7],stage1_5[20],stage1_4[53],stage1_3[54]}
   );
   gpc615_5 gpc55 (
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113]},
      {stage0_4[38]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[8],stage1_5[21],stage1_4[54],stage1_3[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage0_4[39]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[9],stage1_5[22],stage1_4[55],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage0_4[40]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[10],stage1_5[23],stage1_4[56],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage0_4[41]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[11],stage1_5[24],stage1_4[57],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage0_4[42]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[12],stage1_5[25],stage1_4[58],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage0_4[43]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[13],stage1_5[26],stage1_4[59],stage1_3[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[14],stage1_5[27],stage1_4[60]}
   );
   gpc606_5 gpc62 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[15],stage1_5[28],stage1_4[61]}
   );
   gpc606_5 gpc63 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[16],stage1_5[29],stage1_4[62]}
   );
   gpc606_5 gpc64 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[17],stage1_5[30],stage1_4[63]}
   );
   gpc606_5 gpc65 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[18],stage1_5[31],stage1_4[64]}
   );
   gpc606_5 gpc66 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[19],stage1_5[32],stage1_4[65]}
   );
   gpc606_5 gpc67 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[20],stage1_5[33],stage1_4[66]}
   );
   gpc606_5 gpc68 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[21],stage1_5[34],stage1_4[67]}
   );
   gpc606_5 gpc69 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[22],stage1_5[35],stage1_4[68]}
   );
   gpc606_5 gpc70 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[23],stage1_5[36],stage1_4[69]}
   );
   gpc606_5 gpc71 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[24],stage1_5[37],stage1_4[70]}
   );
   gpc606_5 gpc72 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[25],stage1_5[38],stage1_4[71]}
   );
   gpc606_5 gpc73 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[26],stage1_5[39],stage1_4[72]}
   );
   gpc606_5 gpc74 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[27],stage1_5[40],stage1_4[73]}
   );
   gpc606_5 gpc75 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[28],stage1_5[41],stage1_4[74]}
   );
   gpc606_5 gpc76 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[29],stage1_5[42],stage1_4[75]}
   );
   gpc606_5 gpc77 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[30],stage1_5[43],stage1_4[76]}
   );
   gpc606_5 gpc78 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[31],stage1_5[44],stage1_4[77]}
   );
   gpc606_5 gpc79 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[32],stage1_5[45],stage1_4[78]}
   );
   gpc606_5 gpc80 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[19],stage1_7[27],stage1_6[33],stage1_5[46]}
   );
   gpc606_5 gpc81 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[20],stage1_7[28],stage1_6[34],stage1_5[47]}
   );
   gpc606_5 gpc82 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[21],stage1_7[29],stage1_6[35],stage1_5[48]}
   );
   gpc606_5 gpc83 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[22],stage1_7[30],stage1_6[36],stage1_5[49]}
   );
   gpc606_5 gpc84 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[23],stage1_7[31],stage1_6[37],stage1_5[50]}
   );
   gpc606_5 gpc85 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[24],stage1_7[32],stage1_6[38],stage1_5[51]}
   );
   gpc606_5 gpc86 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[25],stage1_7[33],stage1_6[39],stage1_5[52]}
   );
   gpc606_5 gpc87 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[26],stage1_7[34],stage1_6[40],stage1_5[53]}
   );
   gpc606_5 gpc88 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[27],stage1_7[35],stage1_6[41],stage1_5[54]}
   );
   gpc615_5 gpc89 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[28],stage1_7[36],stage1_6[42]}
   );
   gpc615_5 gpc90 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[29],stage1_7[37],stage1_6[43]}
   );
   gpc615_5 gpc91 (
      {stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127], stage0_6[128]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[30],stage1_7[38],stage1_6[44]}
   );
   gpc615_5 gpc92 (
      {stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132], stage0_6[133]},
      {stage0_7[57]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[12],stage1_8[31],stage1_7[39],stage1_6[45]}
   );
   gpc615_5 gpc93 (
      {stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage0_7[58]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[13],stage1_8[32],stage1_7[40],stage1_6[46]}
   );
   gpc615_5 gpc94 (
      {stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_7[59]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[14],stage1_8[33],stage1_7[41],stage1_6[47]}
   );
   gpc615_5 gpc95 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148]},
      {stage0_7[60]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[15],stage1_8[34],stage1_7[42],stage1_6[48]}
   );
   gpc615_5 gpc96 (
      {stage0_6[149], stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153]},
      {stage0_7[61]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[16],stage1_8[35],stage1_7[43],stage1_6[49]}
   );
   gpc606_5 gpc97 (
      {stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65], stage0_7[66], stage0_7[67]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[8],stage1_9[17],stage1_8[36],stage1_7[44]}
   );
   gpc615_5 gpc98 (
      {stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71], stage0_7[72]},
      {stage0_8[48]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[9],stage1_9[18],stage1_8[37],stage1_7[45]}
   );
   gpc615_5 gpc99 (
      {stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage0_8[49]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[10],stage1_9[19],stage1_8[38],stage1_7[46]}
   );
   gpc615_5 gpc100 (
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82]},
      {stage0_8[50]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[11],stage1_9[20],stage1_8[39],stage1_7[47]}
   );
   gpc615_5 gpc101 (
      {stage0_7[83], stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87]},
      {stage0_8[51]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[12],stage1_9[21],stage1_8[40],stage1_7[48]}
   );
   gpc615_5 gpc102 (
      {stage0_7[88], stage0_7[89], stage0_7[90], stage0_7[91], stage0_7[92]},
      {stage0_8[52]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[13],stage1_9[22],stage1_8[41],stage1_7[49]}
   );
   gpc615_5 gpc103 (
      {stage0_7[93], stage0_7[94], stage0_7[95], stage0_7[96], stage0_7[97]},
      {stage0_8[53]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[14],stage1_9[23],stage1_8[42],stage1_7[50]}
   );
   gpc615_5 gpc104 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[54]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[15],stage1_9[24],stage1_8[43],stage1_7[51]}
   );
   gpc615_5 gpc105 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[55]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[16],stage1_9[25],stage1_8[44],stage1_7[52]}
   );
   gpc615_5 gpc106 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[56]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[17],stage1_9[26],stage1_8[45],stage1_7[53]}
   );
   gpc615_5 gpc107 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[57]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[18],stage1_9[27],stage1_8[46],stage1_7[54]}
   );
   gpc615_5 gpc108 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[58]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[19],stage1_9[28],stage1_8[47],stage1_7[55]}
   );
   gpc615_5 gpc109 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[59]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[20],stage1_9[29],stage1_8[48],stage1_7[56]}
   );
   gpc615_5 gpc110 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[60]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[21],stage1_9[30],stage1_8[49],stage1_7[57]}
   );
   gpc615_5 gpc111 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[61]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[22],stage1_9[31],stage1_8[50],stage1_7[58]}
   );
   gpc615_5 gpc112 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[62]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[23],stage1_9[32],stage1_8[51],stage1_7[59]}
   );
   gpc615_5 gpc113 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[63]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[24],stage1_9[33],stage1_8[52],stage1_7[60]}
   );
   gpc615_5 gpc114 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[64]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[25],stage1_9[34],stage1_8[53],stage1_7[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[18],stage1_10[26],stage1_9[35],stage1_8[54]}
   );
   gpc606_5 gpc116 (
      {stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[19],stage1_10[27],stage1_9[36],stage1_8[55]}
   );
   gpc606_5 gpc117 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[20],stage1_10[28],stage1_9[37],stage1_8[56]}
   );
   gpc606_5 gpc118 (
      {stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[21],stage1_10[29],stage1_9[38],stage1_8[57]}
   );
   gpc606_5 gpc119 (
      {stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[22],stage1_10[30],stage1_9[39],stage1_8[58]}
   );
   gpc606_5 gpc120 (
      {stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[23],stage1_10[31],stage1_9[40],stage1_8[59]}
   );
   gpc606_5 gpc121 (
      {stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[24],stage1_10[32],stage1_9[41],stage1_8[60]}
   );
   gpc606_5 gpc122 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[25],stage1_10[33],stage1_9[42],stage1_8[61]}
   );
   gpc606_5 gpc123 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[26],stage1_10[34],stage1_9[43],stage1_8[62]}
   );
   gpc606_5 gpc124 (
      {stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[27],stage1_10[35],stage1_9[44],stage1_8[63]}
   );
   gpc606_5 gpc125 (
      {stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[28],stage1_10[36],stage1_9[45],stage1_8[64]}
   );
   gpc606_5 gpc126 (
      {stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[29],stage1_10[37],stage1_9[46],stage1_8[65]}
   );
   gpc606_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[30],stage1_10[38],stage1_9[47],stage1_8[66]}
   );
   gpc606_5 gpc128 (
      {stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[31],stage1_10[39],stage1_9[48],stage1_8[67]}
   );
   gpc606_5 gpc129 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[14],stage1_11[32],stage1_10[40],stage1_9[49]}
   );
   gpc606_5 gpc130 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[15],stage1_11[33],stage1_10[41],stage1_9[50]}
   );
   gpc606_5 gpc131 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[16],stage1_11[34],stage1_10[42],stage1_9[51]}
   );
   gpc606_5 gpc132 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[17],stage1_11[35],stage1_10[43],stage1_9[52]}
   );
   gpc606_5 gpc133 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[18],stage1_11[36],stage1_10[44],stage1_9[53]}
   );
   gpc606_5 gpc134 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[19],stage1_11[37],stage1_10[45],stage1_9[54]}
   );
   gpc606_5 gpc135 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[20],stage1_11[38],stage1_10[46],stage1_9[55]}
   );
   gpc606_5 gpc136 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[21],stage1_11[39],stage1_10[47],stage1_9[56]}
   );
   gpc606_5 gpc137 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[22],stage1_11[40],stage1_10[48],stage1_9[57]}
   );
   gpc615_5 gpc138 (
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88]},
      {stage0_11[54]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[23],stage1_11[41],stage1_10[49]}
   );
   gpc615_5 gpc139 (
      {stage0_10[89], stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93]},
      {stage0_11[55]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[24],stage1_11[42],stage1_10[50]}
   );
   gpc615_5 gpc140 (
      {stage0_10[94], stage0_10[95], stage0_10[96], stage0_10[97], stage0_10[98]},
      {stage0_11[56]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[11],stage1_12[25],stage1_11[43],stage1_10[51]}
   );
   gpc615_5 gpc141 (
      {stage0_10[99], stage0_10[100], stage0_10[101], stage0_10[102], stage0_10[103]},
      {stage0_11[57]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[12],stage1_12[26],stage1_11[44],stage1_10[52]}
   );
   gpc615_5 gpc142 (
      {stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107], stage0_10[108]},
      {stage0_11[58]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[13],stage1_12[27],stage1_11[45],stage1_10[53]}
   );
   gpc615_5 gpc143 (
      {stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage0_11[59]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[14],stage1_12[28],stage1_11[46],stage1_10[54]}
   );
   gpc615_5 gpc144 (
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118]},
      {stage0_11[60]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[15],stage1_12[29],stage1_11[47],stage1_10[55]}
   );
   gpc615_5 gpc145 (
      {stage0_10[119], stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123]},
      {stage0_11[61]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[16],stage1_12[30],stage1_11[48],stage1_10[56]}
   );
   gpc606_5 gpc146 (
      {stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[8],stage1_13[17],stage1_12[31],stage1_11[49]}
   );
   gpc606_5 gpc147 (
      {stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[9],stage1_13[18],stage1_12[32],stage1_11[50]}
   );
   gpc606_5 gpc148 (
      {stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[10],stage1_13[19],stage1_12[33],stage1_11[51]}
   );
   gpc606_5 gpc149 (
      {stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[11],stage1_13[20],stage1_12[34],stage1_11[52]}
   );
   gpc606_5 gpc150 (
      {stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[12],stage1_13[21],stage1_12[35],stage1_11[53]}
   );
   gpc606_5 gpc151 (
      {stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[13],stage1_13[22],stage1_12[36],stage1_11[54]}
   );
   gpc606_5 gpc152 (
      {stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[14],stage1_13[23],stage1_12[37],stage1_11[55]}
   );
   gpc606_5 gpc153 (
      {stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[15],stage1_13[24],stage1_12[38],stage1_11[56]}
   );
   gpc606_5 gpc154 (
      {stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[16],stage1_13[25],stage1_12[39],stage1_11[57]}
   );
   gpc606_5 gpc155 (
      {stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[17],stage1_13[26],stage1_12[40],stage1_11[58]}
   );
   gpc606_5 gpc156 (
      {stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[18],stage1_13[27],stage1_12[41],stage1_11[59]}
   );
   gpc606_5 gpc157 (
      {stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[19],stage1_13[28],stage1_12[42],stage1_11[60]}
   );
   gpc615_5 gpc158 (
      {stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138]},
      {stage0_12[48]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[20],stage1_13[29],stage1_12[43],stage1_11[61]}
   );
   gpc615_5 gpc159 (
      {stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage0_12[49]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[21],stage1_13[30],stage1_12[44],stage1_11[62]}
   );
   gpc606_5 gpc160 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[14],stage1_14[22],stage1_13[31],stage1_12[45]}
   );
   gpc606_5 gpc161 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[15],stage1_14[23],stage1_13[32],stage1_12[46]}
   );
   gpc606_5 gpc162 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[16],stage1_14[24],stage1_13[33],stage1_12[47]}
   );
   gpc606_5 gpc163 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[17],stage1_14[25],stage1_13[34],stage1_12[48]}
   );
   gpc606_5 gpc164 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[18],stage1_14[26],stage1_13[35],stage1_12[49]}
   );
   gpc606_5 gpc165 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[19],stage1_14[27],stage1_13[36],stage1_12[50]}
   );
   gpc606_5 gpc166 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[20],stage1_14[28],stage1_13[37],stage1_12[51]}
   );
   gpc606_5 gpc167 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[21],stage1_14[29],stage1_13[38],stage1_12[52]}
   );
   gpc606_5 gpc168 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[22],stage1_14[30],stage1_13[39],stage1_12[53]}
   );
   gpc606_5 gpc169 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[23],stage1_14[31],stage1_13[40],stage1_12[54]}
   );
   gpc606_5 gpc170 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[24],stage1_14[32],stage1_13[41],stage1_12[55]}
   );
   gpc606_5 gpc171 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[25],stage1_14[33],stage1_13[42],stage1_12[56]}
   );
   gpc606_5 gpc172 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[26],stage1_14[34],stage1_13[43],stage1_12[57]}
   );
   gpc606_5 gpc173 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[27],stage1_14[35],stage1_13[44],stage1_12[58]}
   );
   gpc606_5 gpc174 (
      {stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[28],stage1_14[36],stage1_13[45],stage1_12[59]}
   );
   gpc606_5 gpc175 (
      {stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[29],stage1_14[37],stage1_13[46],stage1_12[60]}
   );
   gpc606_5 gpc176 (
      {stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[30],stage1_14[38],stage1_13[47],stage1_12[61]}
   );
   gpc606_5 gpc177 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[31],stage1_14[39],stage1_13[48],stage1_12[62]}
   );
   gpc606_5 gpc178 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[18],stage1_15[32],stage1_14[40],stage1_13[49]}
   );
   gpc606_5 gpc179 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[19],stage1_15[33],stage1_14[41],stage1_13[50]}
   );
   gpc606_5 gpc180 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[20],stage1_15[34],stage1_14[42],stage1_13[51]}
   );
   gpc606_5 gpc181 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[21],stage1_15[35],stage1_14[43],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[22],stage1_15[36],stage1_14[44],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[23],stage1_15[37],stage1_14[45],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[24],stage1_15[38],stage1_14[46],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[25],stage1_15[39],stage1_14[47],stage1_13[56]}
   );
   gpc615_5 gpc186 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112]},
      {stage0_15[48]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[8],stage1_16[26],stage1_15[40],stage1_14[48]}
   );
   gpc615_5 gpc187 (
      {stage0_14[113], stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117]},
      {stage0_15[49]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[9],stage1_16[27],stage1_15[41],stage1_14[49]}
   );
   gpc615_5 gpc188 (
      {stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121], stage0_14[122]},
      {stage0_15[50]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[10],stage1_16[28],stage1_15[42],stage1_14[50]}
   );
   gpc615_5 gpc189 (
      {stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage0_15[51]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[11],stage1_16[29],stage1_15[43],stage1_14[51]}
   );
   gpc615_5 gpc190 (
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[52]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[12],stage1_16[30],stage1_15[44],stage1_14[52]}
   );
   gpc615_5 gpc191 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_15[53]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[13],stage1_16[31],stage1_15[45],stage1_14[53]}
   );
   gpc615_5 gpc192 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142]},
      {stage0_15[54]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[14],stage1_16[32],stage1_15[46],stage1_14[54]}
   );
   gpc615_5 gpc193 (
      {stage0_14[143], stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147]},
      {stage0_15[55]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[15],stage1_16[33],stage1_15[47],stage1_14[55]}
   );
   gpc615_5 gpc194 (
      {stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151], stage0_14[152]},
      {stage0_15[56]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[16],stage1_16[34],stage1_15[48],stage1_14[56]}
   );
   gpc615_5 gpc195 (
      {stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage0_15[57]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[17],stage1_16[35],stage1_15[49],stage1_14[57]}
   );
   gpc615_5 gpc196 (
      {stage0_15[58], stage0_15[59], stage0_15[60], stage0_15[61], stage0_15[62]},
      {stage0_16[60]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[10],stage1_17[18],stage1_16[36],stage1_15[50]}
   );
   gpc615_5 gpc197 (
      {stage0_15[63], stage0_15[64], stage0_15[65], stage0_15[66], stage0_15[67]},
      {stage0_16[61]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[11],stage1_17[19],stage1_16[37],stage1_15[51]}
   );
   gpc615_5 gpc198 (
      {stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71], stage0_15[72]},
      {stage0_16[62]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[12],stage1_17[20],stage1_16[38],stage1_15[52]}
   );
   gpc615_5 gpc199 (
      {stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage0_16[63]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[13],stage1_17[21],stage1_16[39],stage1_15[53]}
   );
   gpc615_5 gpc200 (
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82]},
      {stage0_16[64]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[14],stage1_17[22],stage1_16[40],stage1_15[54]}
   );
   gpc615_5 gpc201 (
      {stage0_15[83], stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87]},
      {stage0_16[65]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[15],stage1_17[23],stage1_16[41],stage1_15[55]}
   );
   gpc615_5 gpc202 (
      {stage0_15[88], stage0_15[89], stage0_15[90], stage0_15[91], stage0_15[92]},
      {stage0_16[66]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[16],stage1_17[24],stage1_16[42],stage1_15[56]}
   );
   gpc615_5 gpc203 (
      {stage0_15[93], stage0_15[94], stage0_15[95], stage0_15[96], stage0_15[97]},
      {stage0_16[67]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[17],stage1_17[25],stage1_16[43],stage1_15[57]}
   );
   gpc615_5 gpc204 (
      {stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101], stage0_15[102]},
      {stage0_16[68]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[18],stage1_17[26],stage1_16[44],stage1_15[58]}
   );
   gpc615_5 gpc205 (
      {stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage0_16[69]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[19],stage1_17[27],stage1_16[45],stage1_15[59]}
   );
   gpc615_5 gpc206 (
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112]},
      {stage0_16[70]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[20],stage1_17[28],stage1_16[46],stage1_15[60]}
   );
   gpc615_5 gpc207 (
      {stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117]},
      {stage0_16[71]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[21],stage1_17[29],stage1_16[47],stage1_15[61]}
   );
   gpc615_5 gpc208 (
      {stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121], stage0_15[122]},
      {stage0_16[72]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[22],stage1_17[30],stage1_16[48],stage1_15[62]}
   );
   gpc615_5 gpc209 (
      {stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126], stage0_15[127]},
      {stage0_16[73]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[23],stage1_17[31],stage1_16[49],stage1_15[63]}
   );
   gpc606_5 gpc210 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[14],stage1_18[24],stage1_17[32],stage1_16[50]}
   );
   gpc606_5 gpc211 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[15],stage1_18[25],stage1_17[33],stage1_16[51]}
   );
   gpc606_5 gpc212 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[16],stage1_18[26],stage1_17[34],stage1_16[52]}
   );
   gpc606_5 gpc213 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[17],stage1_18[27],stage1_17[35],stage1_16[53]}
   );
   gpc606_5 gpc214 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[18],stage1_18[28],stage1_17[36],stage1_16[54]}
   );
   gpc606_5 gpc215 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[19],stage1_18[29],stage1_17[37],stage1_16[55]}
   );
   gpc606_5 gpc216 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[20],stage1_18[30],stage1_17[38],stage1_16[56]}
   );
   gpc606_5 gpc217 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[21],stage1_18[31],stage1_17[39],stage1_16[57]}
   );
   gpc606_5 gpc218 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[22],stage1_18[32],stage1_17[40],stage1_16[58]}
   );
   gpc606_5 gpc219 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[23],stage1_18[33],stage1_17[41],stage1_16[59]}
   );
   gpc606_5 gpc220 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[24],stage1_18[34],stage1_17[42],stage1_16[60]}
   );
   gpc606_5 gpc221 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[25],stage1_18[35],stage1_17[43],stage1_16[61]}
   );
   gpc606_5 gpc222 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[26],stage1_18[36],stage1_17[44],stage1_16[62]}
   );
   gpc606_5 gpc223 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[27],stage1_18[37],stage1_17[45],stage1_16[63]}
   );
   gpc606_5 gpc224 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[14],stage1_19[28],stage1_18[38],stage1_17[46]}
   );
   gpc606_5 gpc225 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[15],stage1_19[29],stage1_18[39],stage1_17[47]}
   );
   gpc606_5 gpc226 (
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[2],stage1_20[16],stage1_19[30],stage1_18[40]}
   );
   gpc606_5 gpc227 (
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[3],stage1_20[17],stage1_19[31],stage1_18[41]}
   );
   gpc606_5 gpc228 (
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[4],stage1_20[18],stage1_19[32],stage1_18[42]}
   );
   gpc606_5 gpc229 (
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[5],stage1_20[19],stage1_19[33],stage1_18[43]}
   );
   gpc606_5 gpc230 (
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[6],stage1_20[20],stage1_19[34],stage1_18[44]}
   );
   gpc606_5 gpc231 (
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[7],stage1_20[21],stage1_19[35],stage1_18[45]}
   );
   gpc606_5 gpc232 (
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[8],stage1_20[22],stage1_19[36],stage1_18[46]}
   );
   gpc615_5 gpc233 (
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130]},
      {stage0_19[12]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[9],stage1_20[23],stage1_19[37],stage1_18[47]}
   );
   gpc615_5 gpc234 (
      {stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_19[13]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[10],stage1_20[24],stage1_19[38],stage1_18[48]}
   );
   gpc615_5 gpc235 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140]},
      {stage0_19[14]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[11],stage1_20[25],stage1_19[39],stage1_18[49]}
   );
   gpc615_5 gpc236 (
      {stage0_18[141], stage0_18[142], stage0_18[143], stage0_18[144], stage0_18[145]},
      {stage0_19[15]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[12],stage1_20[26],stage1_19[40],stage1_18[50]}
   );
   gpc615_5 gpc237 (
      {stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149], stage0_18[150]},
      {stage0_19[16]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[13],stage1_20[27],stage1_19[41],stage1_18[51]}
   );
   gpc207_4 gpc238 (
      {stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage0_21[0], stage0_21[1]},
      {stage1_22[12],stage1_21[14],stage1_20[28],stage1_19[42]}
   );
   gpc207_4 gpc239 (
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29], stage0_19[30]},
      {stage0_21[2], stage0_21[3]},
      {stage1_22[13],stage1_21[15],stage1_20[29],stage1_19[43]}
   );
   gpc207_4 gpc240 (
      {stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35], stage0_19[36], stage0_19[37]},
      {stage0_21[4], stage0_21[5]},
      {stage1_22[14],stage1_21[16],stage1_20[30],stage1_19[44]}
   );
   gpc207_4 gpc241 (
      {stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41], stage0_19[42], stage0_19[43], stage0_19[44]},
      {stage0_21[6], stage0_21[7]},
      {stage1_22[15],stage1_21[17],stage1_20[31],stage1_19[45]}
   );
   gpc606_5 gpc242 (
      {stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50]},
      {stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13]},
      {stage1_23[0],stage1_22[16],stage1_21[18],stage1_20[32],stage1_19[46]}
   );
   gpc606_5 gpc243 (
      {stage0_19[51], stage0_19[52], stage0_19[53], stage0_19[54], stage0_19[55], stage0_19[56]},
      {stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19]},
      {stage1_23[1],stage1_22[17],stage1_21[19],stage1_20[33],stage1_19[47]}
   );
   gpc606_5 gpc244 (
      {stage0_19[57], stage0_19[58], stage0_19[59], stage0_19[60], stage0_19[61], stage0_19[62]},
      {stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25]},
      {stage1_23[2],stage1_22[18],stage1_21[20],stage1_20[34],stage1_19[48]}
   );
   gpc606_5 gpc245 (
      {stage0_19[63], stage0_19[64], stage0_19[65], stage0_19[66], stage0_19[67], stage0_19[68]},
      {stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage1_23[3],stage1_22[19],stage1_21[21],stage1_20[35],stage1_19[49]}
   );
   gpc606_5 gpc246 (
      {stage0_19[69], stage0_19[70], stage0_19[71], stage0_19[72], stage0_19[73], stage0_19[74]},
      {stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37]},
      {stage1_23[4],stage1_22[20],stage1_21[22],stage1_20[36],stage1_19[50]}
   );
   gpc606_5 gpc247 (
      {stage0_19[75], stage0_19[76], stage0_19[77], stage0_19[78], stage0_19[79], stage0_19[80]},
      {stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43]},
      {stage1_23[5],stage1_22[21],stage1_21[23],stage1_20[37],stage1_19[51]}
   );
   gpc606_5 gpc248 (
      {stage0_19[81], stage0_19[82], stage0_19[83], stage0_19[84], stage0_19[85], stage0_19[86]},
      {stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49]},
      {stage1_23[6],stage1_22[22],stage1_21[24],stage1_20[38],stage1_19[52]}
   );
   gpc606_5 gpc249 (
      {stage0_19[87], stage0_19[88], stage0_19[89], stage0_19[90], stage0_19[91], stage0_19[92]},
      {stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54], stage0_21[55]},
      {stage1_23[7],stage1_22[23],stage1_21[25],stage1_20[39],stage1_19[53]}
   );
   gpc606_5 gpc250 (
      {stage0_19[93], stage0_19[94], stage0_19[95], stage0_19[96], stage0_19[97], stage0_19[98]},
      {stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60], stage0_21[61]},
      {stage1_23[8],stage1_22[24],stage1_21[26],stage1_20[40],stage1_19[54]}
   );
   gpc606_5 gpc251 (
      {stage0_19[99], stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104]},
      {stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66], stage0_21[67]},
      {stage1_23[9],stage1_22[25],stage1_21[27],stage1_20[41],stage1_19[55]}
   );
   gpc606_5 gpc252 (
      {stage0_19[105], stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110]},
      {stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72], stage0_21[73]},
      {stage1_23[10],stage1_22[26],stage1_21[28],stage1_20[42],stage1_19[56]}
   );
   gpc606_5 gpc253 (
      {stage0_19[111], stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116]},
      {stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78], stage0_21[79]},
      {stage1_23[11],stage1_22[27],stage1_21[29],stage1_20[43],stage1_19[57]}
   );
   gpc606_5 gpc254 (
      {stage0_19[117], stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122]},
      {stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84], stage0_21[85]},
      {stage1_23[12],stage1_22[28],stage1_21[30],stage1_20[44],stage1_19[58]}
   );
   gpc606_5 gpc255 (
      {stage0_19[123], stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128]},
      {stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90], stage0_21[91]},
      {stage1_23[13],stage1_22[29],stage1_21[31],stage1_20[45],stage1_19[59]}
   );
   gpc606_5 gpc256 (
      {stage0_19[129], stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134]},
      {stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97]},
      {stage1_23[14],stage1_22[30],stage1_21[32],stage1_20[46],stage1_19[60]}
   );
   gpc606_5 gpc257 (
      {stage0_19[135], stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140]},
      {stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103]},
      {stage1_23[15],stage1_22[31],stage1_21[33],stage1_20[47],stage1_19[61]}
   );
   gpc615_5 gpc258 (
      {stage0_19[141], stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145]},
      {stage0_20[72]},
      {stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109]},
      {stage1_23[16],stage1_22[32],stage1_21[34],stage1_20[48],stage1_19[62]}
   );
   gpc615_5 gpc259 (
      {stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149], stage0_19[150]},
      {stage0_20[73]},
      {stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage1_23[17],stage1_22[33],stage1_21[35],stage1_20[49],stage1_19[63]}
   );
   gpc615_5 gpc260 (
      {stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage0_20[74]},
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121]},
      {stage1_23[18],stage1_22[34],stage1_21[36],stage1_20[50],stage1_19[64]}
   );
   gpc606_5 gpc261 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[19],stage1_22[35],stage1_21[37],stage1_20[51]}
   );
   gpc606_5 gpc262 (
      {stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[20],stage1_22[36],stage1_21[38],stage1_20[52]}
   );
   gpc606_5 gpc263 (
      {stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[21],stage1_22[37],stage1_21[39],stage1_20[53]}
   );
   gpc606_5 gpc264 (
      {stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[22],stage1_22[38],stage1_21[40],stage1_20[54]}
   );
   gpc606_5 gpc265 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[23],stage1_22[39],stage1_21[41],stage1_20[55]}
   );
   gpc606_5 gpc266 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[24],stage1_22[40],stage1_21[42],stage1_20[56]}
   );
   gpc606_5 gpc267 (
      {stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[25],stage1_22[41],stage1_21[43],stage1_20[57]}
   );
   gpc606_5 gpc268 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121], stage0_20[122]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[26],stage1_22[42],stage1_21[44],stage1_20[58]}
   );
   gpc606_5 gpc269 (
      {stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[27],stage1_22[43],stage1_21[45],stage1_20[59]}
   );
   gpc606_5 gpc270 (
      {stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[28],stage1_22[44],stage1_21[46],stage1_20[60]}
   );
   gpc606_5 gpc271 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[29],stage1_22[45],stage1_21[47],stage1_20[61]}
   );
   gpc606_5 gpc272 (
      {stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[30],stage1_22[46],stage1_21[48],stage1_20[62]}
   );
   gpc606_5 gpc273 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151], stage0_20[152]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[31],stage1_22[47],stage1_21[49],stage1_20[63]}
   );
   gpc606_5 gpc274 (
      {stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[32],stage1_22[48],stage1_21[50],stage1_20[64]}
   );
   gpc615_5 gpc275 (
      {stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_22[84]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[14],stage1_23[33],stage1_22[49],stage1_21[51]}
   );
   gpc615_5 gpc276 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_22[85]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[15],stage1_23[34],stage1_22[50],stage1_21[52]}
   );
   gpc615_5 gpc277 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136]},
      {stage0_22[86]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[16],stage1_23[35],stage1_22[51],stage1_21[53]}
   );
   gpc615_5 gpc278 (
      {stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_22[87]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[17],stage1_23[36],stage1_22[52],stage1_21[54]}
   );
   gpc615_5 gpc279 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146]},
      {stage0_22[88]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[18],stage1_23[37],stage1_22[53],stage1_21[55]}
   );
   gpc606_5 gpc280 (
      {stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[19],stage1_23[38],stage1_22[54]}
   );
   gpc606_5 gpc281 (
      {stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[20],stage1_23[39],stage1_22[55]}
   );
   gpc606_5 gpc282 (
      {stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[21],stage1_23[40],stage1_22[56]}
   );
   gpc606_5 gpc283 (
      {stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[22],stage1_23[41],stage1_22[57]}
   );
   gpc606_5 gpc284 (
      {stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[23],stage1_23[42],stage1_22[58]}
   );
   gpc606_5 gpc285 (
      {stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[24],stage1_23[43],stage1_22[59]}
   );
   gpc606_5 gpc286 (
      {stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[11],stage1_24[25],stage1_23[44],stage1_22[60]}
   );
   gpc606_5 gpc287 (
      {stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[12],stage1_24[26],stage1_23[45],stage1_22[61]}
   );
   gpc615_5 gpc288 (
      {stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141]},
      {stage0_23[30]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[13],stage1_24[27],stage1_23[46],stage1_22[62]}
   );
   gpc615_5 gpc289 (
      {stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage0_23[31]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[14],stage1_24[28],stage1_23[47],stage1_22[63]}
   );
   gpc615_5 gpc290 (
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151]},
      {stage0_23[32]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[15],stage1_24[29],stage1_23[48],stage1_22[64]}
   );
   gpc615_5 gpc291 (
      {stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156]},
      {stage0_23[33]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[16],stage1_24[30],stage1_23[49],stage1_22[65]}
   );
   gpc615_5 gpc292 (
      {stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage0_23[34]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[17],stage1_24[31],stage1_23[50],stage1_22[66]}
   );
   gpc606_5 gpc293 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[13],stage1_25[18],stage1_24[32],stage1_23[51]}
   );
   gpc606_5 gpc294 (
      {stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[14],stage1_25[19],stage1_24[33],stage1_23[52]}
   );
   gpc606_5 gpc295 (
      {stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[15],stage1_25[20],stage1_24[34],stage1_23[53]}
   );
   gpc606_5 gpc296 (
      {stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[16],stage1_25[21],stage1_24[35],stage1_23[54]}
   );
   gpc606_5 gpc297 (
      {stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[17],stage1_25[22],stage1_24[36],stage1_23[55]}
   );
   gpc606_5 gpc298 (
      {stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[18],stage1_25[23],stage1_24[37],stage1_23[56]}
   );
   gpc606_5 gpc299 (
      {stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[19],stage1_25[24],stage1_24[38],stage1_23[57]}
   );
   gpc606_5 gpc300 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[7],stage1_26[20],stage1_25[25],stage1_24[39]}
   );
   gpc606_5 gpc301 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[8],stage1_26[21],stage1_25[26],stage1_24[40]}
   );
   gpc606_5 gpc302 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[9],stage1_26[22],stage1_25[27],stage1_24[41]}
   );
   gpc606_5 gpc303 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[10],stage1_26[23],stage1_25[28],stage1_24[42]}
   );
   gpc606_5 gpc304 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[11],stage1_26[24],stage1_25[29],stage1_24[43]}
   );
   gpc606_5 gpc305 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[12],stage1_26[25],stage1_25[30],stage1_24[44]}
   );
   gpc606_5 gpc306 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[13],stage1_26[26],stage1_25[31],stage1_24[45]}
   );
   gpc606_5 gpc307 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[14],stage1_26[27],stage1_25[32],stage1_24[46]}
   );
   gpc615_5 gpc308 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46]},
      {stage0_26[48]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[15],stage1_26[28],stage1_25[33]}
   );
   gpc615_5 gpc309 (
      {stage0_25[47], stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51]},
      {stage0_26[49]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[16],stage1_26[29],stage1_25[34]}
   );
   gpc615_5 gpc310 (
      {stage0_25[52], stage0_25[53], stage0_25[54], stage0_25[55], stage0_25[56]},
      {stage0_26[50]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[17],stage1_26[30],stage1_25[35]}
   );
   gpc615_5 gpc311 (
      {stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_26[51]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[18],stage1_26[31],stage1_25[36]}
   );
   gpc615_5 gpc312 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66]},
      {stage0_26[52]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[19],stage1_26[32],stage1_25[37]}
   );
   gpc615_5 gpc313 (
      {stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_26[53]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[13],stage1_27[20],stage1_26[33],stage1_25[38]}
   );
   gpc615_5 gpc314 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76]},
      {stage0_26[54]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[14],stage1_27[21],stage1_26[34],stage1_25[39]}
   );
   gpc615_5 gpc315 (
      {stage0_25[77], stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81]},
      {stage0_26[55]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[15],stage1_27[22],stage1_26[35],stage1_25[40]}
   );
   gpc615_5 gpc316 (
      {stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85], stage0_25[86]},
      {stage0_26[56]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[16],stage1_27[23],stage1_26[36],stage1_25[41]}
   );
   gpc615_5 gpc317 (
      {stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_26[57]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[17],stage1_27[24],stage1_26[37],stage1_25[42]}
   );
   gpc615_5 gpc318 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96]},
      {stage0_26[58]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[18],stage1_27[25],stage1_26[38],stage1_25[43]}
   );
   gpc615_5 gpc319 (
      {stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_26[59]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[19],stage1_27[26],stage1_26[39],stage1_25[44]}
   );
   gpc615_5 gpc320 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106]},
      {stage0_26[60]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[20],stage1_27[27],stage1_26[40],stage1_25[45]}
   );
   gpc615_5 gpc321 (
      {stage0_25[107], stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111]},
      {stage0_26[61]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[21],stage1_27[28],stage1_26[41],stage1_25[46]}
   );
   gpc615_5 gpc322 (
      {stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116]},
      {stage0_26[62]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[22],stage1_27[29],stage1_26[42],stage1_25[47]}
   );
   gpc615_5 gpc323 (
      {stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_26[63]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[23],stage1_27[30],stage1_26[43],stage1_25[48]}
   );
   gpc615_5 gpc324 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126]},
      {stage0_26[64]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[24],stage1_27[31],stage1_26[44],stage1_25[49]}
   );
   gpc606_5 gpc325 (
      {stage0_26[65], stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[17],stage1_28[25],stage1_27[32],stage1_26[45]}
   );
   gpc606_5 gpc326 (
      {stage0_26[71], stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[18],stage1_28[26],stage1_27[33],stage1_26[46]}
   );
   gpc606_5 gpc327 (
      {stage0_26[77], stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[19],stage1_28[27],stage1_27[34],stage1_26[47]}
   );
   gpc606_5 gpc328 (
      {stage0_26[83], stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[20],stage1_28[28],stage1_27[35],stage1_26[48]}
   );
   gpc606_5 gpc329 (
      {stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[21],stage1_28[29],stage1_27[36],stage1_26[49]}
   );
   gpc606_5 gpc330 (
      {stage0_26[95], stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[22],stage1_28[30],stage1_27[37],stage1_26[50]}
   );
   gpc606_5 gpc331 (
      {stage0_26[101], stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[23],stage1_28[31],stage1_27[38],stage1_26[51]}
   );
   gpc606_5 gpc332 (
      {stage0_26[107], stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[24],stage1_28[32],stage1_27[39],stage1_26[52]}
   );
   gpc606_5 gpc333 (
      {stage0_26[113], stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[25],stage1_28[33],stage1_27[40],stage1_26[53]}
   );
   gpc606_5 gpc334 (
      {stage0_26[119], stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[26],stage1_28[34],stage1_27[41],stage1_26[54]}
   );
   gpc606_5 gpc335 (
      {stage0_26[125], stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[27],stage1_28[35],stage1_27[42],stage1_26[55]}
   );
   gpc606_5 gpc336 (
      {stage0_26[131], stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[28],stage1_28[36],stage1_27[43],stage1_26[56]}
   );
   gpc606_5 gpc337 (
      {stage0_26[137], stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142]},
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage1_30[12],stage1_29[29],stage1_28[37],stage1_27[44],stage1_26[57]}
   );
   gpc606_5 gpc338 (
      {stage0_26[143], stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148]},
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage1_30[13],stage1_29[30],stage1_28[38],stage1_27[45],stage1_26[58]}
   );
   gpc615_5 gpc339 (
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106]},
      {stage0_28[84]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[14],stage1_29[31],stage1_28[39],stage1_27[46]}
   );
   gpc615_5 gpc340 (
      {stage0_27[107], stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111]},
      {stage0_28[85]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[15],stage1_29[32],stage1_28[40],stage1_27[47]}
   );
   gpc615_5 gpc341 (
      {stage0_27[112], stage0_27[113], stage0_27[114], stage0_27[115], stage0_27[116]},
      {stage0_28[86]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[16],stage1_29[33],stage1_28[41],stage1_27[48]}
   );
   gpc615_5 gpc342 (
      {stage0_27[117], stage0_27[118], stage0_27[119], stage0_27[120], stage0_27[121]},
      {stage0_28[87]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[17],stage1_29[34],stage1_28[42],stage1_27[49]}
   );
   gpc615_5 gpc343 (
      {stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125], stage0_27[126]},
      {stage0_28[88]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[18],stage1_29[35],stage1_28[43],stage1_27[50]}
   );
   gpc615_5 gpc344 (
      {stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage0_28[89]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[19],stage1_29[36],stage1_28[44],stage1_27[51]}
   );
   gpc615_5 gpc345 (
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136]},
      {stage0_28[90]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[20],stage1_29[37],stage1_28[45],stage1_27[52]}
   );
   gpc615_5 gpc346 (
      {stage0_27[137], stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141]},
      {stage0_28[91]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[21],stage1_29[38],stage1_28[46],stage1_27[53]}
   );
   gpc606_5 gpc347 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[8],stage1_30[22],stage1_29[39],stage1_28[47]}
   );
   gpc606_5 gpc348 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[9],stage1_30[23],stage1_29[40],stage1_28[48]}
   );
   gpc606_5 gpc349 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[10],stage1_30[24],stage1_29[41],stage1_28[49]}
   );
   gpc606_5 gpc350 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[11],stage1_30[25],stage1_29[42],stage1_28[50]}
   );
   gpc606_5 gpc351 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[12],stage1_30[26],stage1_29[43],stage1_28[51]}
   );
   gpc606_5 gpc352 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[13],stage1_30[27],stage1_29[44],stage1_28[52]}
   );
   gpc606_5 gpc353 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[14],stage1_30[28],stage1_29[45],stage1_28[53]}
   );
   gpc606_5 gpc354 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[15],stage1_30[29],stage1_29[46],stage1_28[54]}
   );
   gpc606_5 gpc355 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[8],stage1_31[16],stage1_30[30],stage1_29[47]}
   );
   gpc606_5 gpc356 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[9],stage1_31[17],stage1_30[31],stage1_29[48]}
   );
   gpc606_5 gpc357 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[10],stage1_31[18],stage1_30[32],stage1_29[49]}
   );
   gpc606_5 gpc358 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[11],stage1_31[19],stage1_30[33],stage1_29[50]}
   );
   gpc606_5 gpc359 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[12],stage1_31[20],stage1_30[34],stage1_29[51]}
   );
   gpc606_5 gpc360 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[13],stage1_31[21],stage1_30[35],stage1_29[52]}
   );
   gpc606_5 gpc361 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[14],stage1_31[22],stage1_30[36],stage1_29[53]}
   );
   gpc606_5 gpc362 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[15],stage1_31[23],stage1_30[37],stage1_29[54]}
   );
   gpc606_5 gpc363 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[16],stage1_31[24],stage1_30[38],stage1_29[55]}
   );
   gpc606_5 gpc364 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[17],stage1_31[25],stage1_30[39],stage1_29[56]}
   );
   gpc606_5 gpc365 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[18],stage1_31[26],stage1_30[40],stage1_29[57]}
   );
   gpc606_5 gpc366 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[19],stage1_31[27],stage1_30[41],stage1_29[58]}
   );
   gpc606_5 gpc367 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[20],stage1_31[28],stage1_30[42],stage1_29[59]}
   );
   gpc606_5 gpc368 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[21],stage1_31[29],stage1_30[43],stage1_29[60]}
   );
   gpc606_5 gpc369 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[22],stage1_31[30],stage1_30[44],stage1_29[61]}
   );
   gpc606_5 gpc370 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[23],stage1_31[31],stage1_30[45],stage1_29[62]}
   );
   gpc1406_5 gpc371 (
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[16],stage1_32[24],stage1_31[32],stage1_30[46]}
   );
   gpc207_4 gpc372 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage0_32[4], stage0_32[5]},
      {stage1_33[17],stage1_32[25],stage1_31[33],stage1_30[47]}
   );
   gpc207_4 gpc373 (
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66], stage0_30[67]},
      {stage0_32[6], stage0_32[7]},
      {stage1_33[18],stage1_32[26],stage1_31[34],stage1_30[48]}
   );
   gpc207_4 gpc374 (
      {stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72], stage0_30[73], stage0_30[74]},
      {stage0_32[8], stage0_32[9]},
      {stage1_33[19],stage1_32[27],stage1_31[35],stage1_30[49]}
   );
   gpc207_4 gpc375 (
      {stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81]},
      {stage0_32[10], stage0_32[11]},
      {stage1_33[20],stage1_32[28],stage1_31[36],stage1_30[50]}
   );
   gpc207_4 gpc376 (
      {stage0_30[82], stage0_30[83], stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88]},
      {stage0_32[12], stage0_32[13]},
      {stage1_33[21],stage1_32[29],stage1_31[37],stage1_30[51]}
   );
   gpc207_4 gpc377 (
      {stage0_30[89], stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage0_32[14], stage0_32[15]},
      {stage1_33[22],stage1_32[30],stage1_31[38],stage1_30[52]}
   );
   gpc615_5 gpc378 (
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100]},
      {stage0_31[96]},
      {stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21]},
      {stage1_34[1],stage1_33[23],stage1_32[31],stage1_31[39],stage1_30[53]}
   );
   gpc615_5 gpc379 (
      {stage0_30[101], stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105]},
      {stage0_31[97]},
      {stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27]},
      {stage1_34[2],stage1_33[24],stage1_32[32],stage1_31[40],stage1_30[54]}
   );
   gpc615_5 gpc380 (
      {stage0_30[106], stage0_30[107], stage0_30[108], stage0_30[109], stage0_30[110]},
      {stage0_31[98]},
      {stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33]},
      {stage1_34[3],stage1_33[25],stage1_32[33],stage1_31[41],stage1_30[55]}
   );
   gpc615_5 gpc381 (
      {stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage0_32[34]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[4],stage1_33[26],stage1_32[34],stage1_31[42]}
   );
   gpc615_5 gpc382 (
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108]},
      {stage0_32[35]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[5],stage1_33[27],stage1_32[35],stage1_31[43]}
   );
   gpc606_5 gpc383 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[28],stage1_32[36]}
   );
   gpc606_5 gpc384 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[29],stage1_32[37]}
   );
   gpc606_5 gpc385 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[30],stage1_32[38]}
   );
   gpc615_5 gpc386 (
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58]},
      {stage0_33[13]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[31],stage1_32[39]}
   );
   gpc615_5 gpc387 (
      {stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63]},
      {stage0_33[14]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[32],stage1_32[40]}
   );
   gpc615_5 gpc388 (
      {stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_33[15]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[33],stage1_32[41]}
   );
   gpc615_5 gpc389 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73]},
      {stage0_33[16]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[34],stage1_32[42]}
   );
   gpc615_5 gpc390 (
      {stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78]},
      {stage0_33[17]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[9],stage1_34[13],stage1_33[35],stage1_32[43]}
   );
   gpc615_5 gpc391 (
      {stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage0_33[18]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[10],stage1_34[14],stage1_33[36],stage1_32[44]}
   );
   gpc615_5 gpc392 (
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88]},
      {stage0_33[19]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[11],stage1_34[15],stage1_33[37],stage1_32[45]}
   );
   gpc615_5 gpc393 (
      {stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93]},
      {stage0_33[20]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[12],stage1_34[16],stage1_33[38],stage1_32[46]}
   );
   gpc615_5 gpc394 (
      {stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_33[21]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[13],stage1_34[17],stage1_33[39],stage1_32[47]}
   );
   gpc615_5 gpc395 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103]},
      {stage0_33[22]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[14],stage1_34[18],stage1_33[40],stage1_32[48]}
   );
   gpc615_5 gpc396 (
      {stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108]},
      {stage0_33[23]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[15],stage1_34[19],stage1_33[41],stage1_32[49]}
   );
   gpc615_5 gpc397 (
      {stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage0_33[24]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[16],stage1_34[20],stage1_33[42],stage1_32[50]}
   );
   gpc615_5 gpc398 (
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118]},
      {stage0_33[25]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[17],stage1_34[21],stage1_33[43],stage1_32[51]}
   );
   gpc615_5 gpc399 (
      {stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122], stage0_32[123]},
      {stage0_33[26]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[18],stage1_34[22],stage1_33[44],stage1_32[52]}
   );
   gpc615_5 gpc400 (
      {stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_33[27]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[19],stage1_34[23],stage1_33[45],stage1_32[53]}
   );
   gpc606_5 gpc401 (
      {stage0_33[28], stage0_33[29], stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[18],stage1_35[20],stage1_34[24],stage1_33[46]}
   );
   gpc606_5 gpc402 (
      {stage0_33[34], stage0_33[35], stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[19],stage1_35[21],stage1_34[25],stage1_33[47]}
   );
   gpc606_5 gpc403 (
      {stage0_33[40], stage0_33[41], stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[20],stage1_35[22],stage1_34[26],stage1_33[48]}
   );
   gpc606_5 gpc404 (
      {stage0_33[46], stage0_33[47], stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[21],stage1_35[23],stage1_34[27],stage1_33[49]}
   );
   gpc606_5 gpc405 (
      {stage0_33[52], stage0_33[53], stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[22],stage1_35[24],stage1_34[28],stage1_33[50]}
   );
   gpc606_5 gpc406 (
      {stage0_33[58], stage0_33[59], stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[23],stage1_35[25],stage1_34[29],stage1_33[51]}
   );
   gpc606_5 gpc407 (
      {stage0_33[64], stage0_33[65], stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[24],stage1_35[26],stage1_34[30],stage1_33[52]}
   );
   gpc606_5 gpc408 (
      {stage0_33[70], stage0_33[71], stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[25],stage1_35[27],stage1_34[31],stage1_33[53]}
   );
   gpc606_5 gpc409 (
      {stage0_33[76], stage0_33[77], stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[26],stage1_35[28],stage1_34[32],stage1_33[54]}
   );
   gpc606_5 gpc410 (
      {stage0_33[82], stage0_33[83], stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[27],stage1_35[29],stage1_34[33],stage1_33[55]}
   );
   gpc606_5 gpc411 (
      {stage0_33[88], stage0_33[89], stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[28],stage1_35[30],stage1_34[34],stage1_33[56]}
   );
   gpc606_5 gpc412 (
      {stage0_33[94], stage0_33[95], stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[29],stage1_35[31],stage1_34[35],stage1_33[57]}
   );
   gpc606_5 gpc413 (
      {stage0_33[100], stage0_33[101], stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[30],stage1_35[32],stage1_34[36],stage1_33[58]}
   );
   gpc606_5 gpc414 (
      {stage0_33[106], stage0_33[107], stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[31],stage1_35[33],stage1_34[37],stage1_33[59]}
   );
   gpc606_5 gpc415 (
      {stage0_33[112], stage0_33[113], stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[32],stage1_35[34],stage1_34[38],stage1_33[60]}
   );
   gpc606_5 gpc416 (
      {stage0_33[118], stage0_33[119], stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[33],stage1_35[35],stage1_34[39],stage1_33[61]}
   );
   gpc606_5 gpc417 (
      {stage0_33[124], stage0_33[125], stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[34],stage1_35[36],stage1_34[40],stage1_33[62]}
   );
   gpc606_5 gpc418 (
      {stage0_33[130], stage0_33[131], stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[35],stage1_35[37],stage1_34[41],stage1_33[63]}
   );
   gpc615_5 gpc419 (
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112]},
      {stage0_35[108]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[18],stage1_36[36],stage1_35[38],stage1_34[42]}
   );
   gpc615_5 gpc420 (
      {stage0_34[113], stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117]},
      {stage0_35[109]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[19],stage1_36[37],stage1_35[39],stage1_34[43]}
   );
   gpc615_5 gpc421 (
      {stage0_34[118], stage0_34[119], stage0_34[120], stage0_34[121], stage0_34[122]},
      {stage0_35[110]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[20],stage1_36[38],stage1_35[40],stage1_34[44]}
   );
   gpc615_5 gpc422 (
      {stage0_34[123], stage0_34[124], stage0_34[125], stage0_34[126], stage0_34[127]},
      {stage0_35[111]},
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage1_38[3],stage1_37[21],stage1_36[39],stage1_35[41],stage1_34[45]}
   );
   gpc615_5 gpc423 (
      {stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131], stage0_34[132]},
      {stage0_35[112]},
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage1_38[4],stage1_37[22],stage1_36[40],stage1_35[42],stage1_34[46]}
   );
   gpc615_5 gpc424 (
      {stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage0_35[113]},
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage1_38[5],stage1_37[23],stage1_36[41],stage1_35[43],stage1_34[47]}
   );
   gpc615_5 gpc425 (
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142]},
      {stage0_35[114]},
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage1_38[6],stage1_37[24],stage1_36[42],stage1_35[44],stage1_34[48]}
   );
   gpc615_5 gpc426 (
      {stage0_34[143], stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147]},
      {stage0_35[115]},
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage1_38[7],stage1_37[25],stage1_36[43],stage1_35[45],stage1_34[49]}
   );
   gpc615_5 gpc427 (
      {stage0_34[148], stage0_34[149], stage0_34[150], stage0_34[151], stage0_34[152]},
      {stage0_35[116]},
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage1_38[8],stage1_37[26],stage1_36[44],stage1_35[46],stage1_34[50]}
   );
   gpc615_5 gpc428 (
      {stage0_34[153], stage0_34[154], stage0_34[155], stage0_34[156], stage0_34[157]},
      {stage0_35[117]},
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage1_38[9],stage1_37[27],stage1_36[45],stage1_35[47],stage1_34[51]}
   );
   gpc615_5 gpc429 (
      {stage0_35[118], stage0_35[119], stage0_35[120], stage0_35[121], stage0_35[122]},
      {stage0_36[60]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[10],stage1_37[28],stage1_36[46],stage1_35[48]}
   );
   gpc615_5 gpc430 (
      {stage0_35[123], stage0_35[124], stage0_35[125], stage0_35[126], stage0_35[127]},
      {stage0_36[61]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[11],stage1_37[29],stage1_36[47],stage1_35[49]}
   );
   gpc615_5 gpc431 (
      {stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131], stage0_35[132]},
      {stage0_36[62]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[12],stage1_37[30],stage1_36[48],stage1_35[50]}
   );
   gpc615_5 gpc432 (
      {stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[63]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[13],stage1_37[31],stage1_36[49],stage1_35[51]}
   );
   gpc615_5 gpc433 (
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142]},
      {stage0_36[64]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[14],stage1_37[32],stage1_36[50],stage1_35[52]}
   );
   gpc615_5 gpc434 (
      {stage0_35[143], stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147]},
      {stage0_36[65]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[15],stage1_37[33],stage1_36[51],stage1_35[53]}
   );
   gpc615_5 gpc435 (
      {stage0_35[148], stage0_35[149], stage0_35[150], stage0_35[151], stage0_35[152]},
      {stage0_36[66]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[16],stage1_37[34],stage1_36[52],stage1_35[54]}
   );
   gpc615_5 gpc436 (
      {stage0_35[153], stage0_35[154], stage0_35[155], stage0_35[156], stage0_35[157]},
      {stage0_36[67]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[17],stage1_37[35],stage1_36[53],stage1_35[55]}
   );
   gpc606_5 gpc437 (
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[8],stage1_38[18],stage1_37[36],stage1_36[54]}
   );
   gpc606_5 gpc438 (
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[9],stage1_38[19],stage1_37[37],stage1_36[55]}
   );
   gpc606_5 gpc439 (
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[10],stage1_38[20],stage1_37[38],stage1_36[56]}
   );
   gpc606_5 gpc440 (
      {stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90], stage0_36[91]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[11],stage1_38[21],stage1_37[39],stage1_36[57]}
   );
   gpc606_5 gpc441 (
      {stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96], stage0_36[97]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[12],stage1_38[22],stage1_37[40],stage1_36[58]}
   );
   gpc606_5 gpc442 (
      {stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102], stage0_36[103]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[13],stage1_38[23],stage1_37[41],stage1_36[59]}
   );
   gpc606_5 gpc443 (
      {stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108], stage0_36[109]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[14],stage1_38[24],stage1_37[42],stage1_36[60]}
   );
   gpc606_5 gpc444 (
      {stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114], stage0_36[115]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[15],stage1_38[25],stage1_37[43],stage1_36[61]}
   );
   gpc606_5 gpc445 (
      {stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120], stage0_36[121]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[16],stage1_38[26],stage1_37[44],stage1_36[62]}
   );
   gpc606_5 gpc446 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[17],stage1_38[27],stage1_37[45],stage1_36[63]}
   );
   gpc606_5 gpc447 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[18],stage1_38[28],stage1_37[46],stage1_36[64]}
   );
   gpc606_5 gpc448 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[19],stage1_38[29],stage1_37[47],stage1_36[65]}
   );
   gpc606_5 gpc449 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[20],stage1_38[30],stage1_37[48],stage1_36[66]}
   );
   gpc606_5 gpc450 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[13],stage1_39[21],stage1_38[31],stage1_37[49]}
   );
   gpc606_5 gpc451 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[14],stage1_39[22],stage1_38[32],stage1_37[50]}
   );
   gpc606_5 gpc452 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[15],stage1_39[23],stage1_38[33],stage1_37[51]}
   );
   gpc606_5 gpc453 (
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[16],stage1_39[24],stage1_38[34],stage1_37[52]}
   );
   gpc606_5 gpc454 (
      {stage0_37[72], stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[17],stage1_39[25],stage1_38[35],stage1_37[53]}
   );
   gpc606_5 gpc455 (
      {stage0_37[78], stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[18],stage1_39[26],stage1_38[36],stage1_37[54]}
   );
   gpc606_5 gpc456 (
      {stage0_37[84], stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[19],stage1_39[27],stage1_38[37],stage1_37[55]}
   );
   gpc615_5 gpc457 (
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[20],stage1_39[28],stage1_38[38]}
   );
   gpc615_5 gpc458 (
      {stage0_38[83], stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87]},
      {stage0_39[43]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[8],stage1_40[21],stage1_39[29],stage1_38[39]}
   );
   gpc615_5 gpc459 (
      {stage0_38[88], stage0_38[89], stage0_38[90], stage0_38[91], stage0_38[92]},
      {stage0_39[44]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[9],stage1_40[22],stage1_39[30],stage1_38[40]}
   );
   gpc615_5 gpc460 (
      {stage0_38[93], stage0_38[94], stage0_38[95], stage0_38[96], stage0_38[97]},
      {stage0_39[45]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[10],stage1_40[23],stage1_39[31],stage1_38[41]}
   );
   gpc615_5 gpc461 (
      {stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101], stage0_38[102]},
      {stage0_39[46]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[11],stage1_40[24],stage1_39[32],stage1_38[42]}
   );
   gpc615_5 gpc462 (
      {stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage0_39[47]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[12],stage1_40[25],stage1_39[33],stage1_38[43]}
   );
   gpc615_5 gpc463 (
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112]},
      {stage0_39[48]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[13],stage1_40[26],stage1_39[34],stage1_38[44]}
   );
   gpc615_5 gpc464 (
      {stage0_38[113], stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117]},
      {stage0_39[49]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[14],stage1_40[27],stage1_39[35],stage1_38[45]}
   );
   gpc615_5 gpc465 (
      {stage0_38[118], stage0_38[119], stage0_38[120], stage0_38[121], stage0_38[122]},
      {stage0_39[50]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[15],stage1_40[28],stage1_39[36],stage1_38[46]}
   );
   gpc615_5 gpc466 (
      {stage0_38[123], stage0_38[124], stage0_38[125], stage0_38[126], stage0_38[127]},
      {stage0_39[51]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[16],stage1_40[29],stage1_39[37],stage1_38[47]}
   );
   gpc615_5 gpc467 (
      {stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131], stage0_38[132]},
      {stage0_39[52]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[17],stage1_40[30],stage1_39[38],stage1_38[48]}
   );
   gpc615_5 gpc468 (
      {stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage0_39[53]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[18],stage1_40[31],stage1_39[39],stage1_38[49]}
   );
   gpc615_5 gpc469 (
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142]},
      {stage0_39[54]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[19],stage1_40[32],stage1_39[40],stage1_38[50]}
   );
   gpc615_5 gpc470 (
      {stage0_38[143], stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147]},
      {stage0_39[55]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[20],stage1_40[33],stage1_39[41],stage1_38[51]}
   );
   gpc615_5 gpc471 (
      {stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59], stage0_39[60]},
      {stage0_40[84]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[14],stage1_41[21],stage1_40[34],stage1_39[42]}
   );
   gpc615_5 gpc472 (
      {stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage0_40[85]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[15],stage1_41[22],stage1_40[35],stage1_39[43]}
   );
   gpc615_5 gpc473 (
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70]},
      {stage0_40[86]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[16],stage1_41[23],stage1_40[36],stage1_39[44]}
   );
   gpc615_5 gpc474 (
      {stage0_39[71], stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75]},
      {stage0_40[87]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[17],stage1_41[24],stage1_40[37],stage1_39[45]}
   );
   gpc615_5 gpc475 (
      {stage0_39[76], stage0_39[77], stage0_39[78], stage0_39[79], stage0_39[80]},
      {stage0_40[88]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[18],stage1_41[25],stage1_40[38],stage1_39[46]}
   );
   gpc615_5 gpc476 (
      {stage0_39[81], stage0_39[82], stage0_39[83], stage0_39[84], stage0_39[85]},
      {stage0_40[89]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[19],stage1_41[26],stage1_40[39],stage1_39[47]}
   );
   gpc615_5 gpc477 (
      {stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89], stage0_39[90]},
      {stage0_40[90]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[20],stage1_41[27],stage1_40[40],stage1_39[48]}
   );
   gpc615_5 gpc478 (
      {stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage0_40[91]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[21],stage1_41[28],stage1_40[41],stage1_39[49]}
   );
   gpc615_5 gpc479 (
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100]},
      {stage0_40[92]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[22],stage1_41[29],stage1_40[42],stage1_39[50]}
   );
   gpc615_5 gpc480 (
      {stage0_39[101], stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105]},
      {stage0_40[93]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[23],stage1_41[30],stage1_40[43],stage1_39[51]}
   );
   gpc615_5 gpc481 (
      {stage0_39[106], stage0_39[107], stage0_39[108], stage0_39[109], stage0_39[110]},
      {stage0_40[94]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[24],stage1_41[31],stage1_40[44],stage1_39[52]}
   );
   gpc615_5 gpc482 (
      {stage0_39[111], stage0_39[112], stage0_39[113], stage0_39[114], stage0_39[115]},
      {stage0_40[95]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[25],stage1_41[32],stage1_40[45],stage1_39[53]}
   );
   gpc615_5 gpc483 (
      {stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119], stage0_39[120]},
      {stage0_40[96]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[26],stage1_41[33],stage1_40[46],stage1_39[54]}
   );
   gpc615_5 gpc484 (
      {stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage0_40[97]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[27],stage1_41[34],stage1_40[47],stage1_39[55]}
   );
   gpc615_5 gpc485 (
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130]},
      {stage0_40[98]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[28],stage1_41[35],stage1_40[48],stage1_39[56]}
   );
   gpc615_5 gpc486 (
      {stage0_39[131], stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135]},
      {stage0_40[99]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[29],stage1_41[36],stage1_40[49],stage1_39[57]}
   );
   gpc615_5 gpc487 (
      {stage0_39[136], stage0_39[137], stage0_39[138], stage0_39[139], stage0_39[140]},
      {stage0_40[100]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[30],stage1_41[37],stage1_40[50],stage1_39[58]}
   );
   gpc615_5 gpc488 (
      {stage0_39[141], stage0_39[142], stage0_39[143], stage0_39[144], stage0_39[145]},
      {stage0_40[101]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[31],stage1_41[38],stage1_40[51],stage1_39[59]}
   );
   gpc615_5 gpc489 (
      {stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149], stage0_39[150]},
      {stage0_40[102]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[32],stage1_41[39],stage1_40[52],stage1_39[60]}
   );
   gpc615_5 gpc490 (
      {stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage0_40[103]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[33],stage1_41[40],stage1_40[53],stage1_39[61]}
   );
   gpc606_5 gpc491 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[20],stage1_42[34],stage1_41[41],stage1_40[54]}
   );
   gpc606_5 gpc492 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[21],stage1_42[35],stage1_41[42],stage1_40[55]}
   );
   gpc606_5 gpc493 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[22],stage1_42[36],stage1_41[43],stage1_40[56]}
   );
   gpc606_5 gpc494 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[23],stage1_42[37],stage1_41[44],stage1_40[57]}
   );
   gpc606_5 gpc495 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[24],stage1_42[38],stage1_41[45],stage1_40[58]}
   );
   gpc606_5 gpc496 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[25],stage1_42[39],stage1_41[46],stage1_40[59]}
   );
   gpc606_5 gpc497 (
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[6],stage1_43[26],stage1_42[40],stage1_41[47]}
   );
   gpc606_5 gpc498 (
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[7],stage1_43[27],stage1_42[41],stage1_41[48]}
   );
   gpc606_5 gpc499 (
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[8],stage1_43[28],stage1_42[42],stage1_41[49]}
   );
   gpc606_5 gpc500 (
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[3],stage1_44[9],stage1_43[29],stage1_42[43]}
   );
   gpc606_5 gpc501 (
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[4],stage1_44[10],stage1_43[30],stage1_42[44]}
   );
   gpc606_5 gpc502 (
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[5],stage1_44[11],stage1_43[31],stage1_42[45]}
   );
   gpc606_5 gpc503 (
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[6],stage1_44[12],stage1_43[32],stage1_42[46]}
   );
   gpc606_5 gpc504 (
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[7],stage1_44[13],stage1_43[33],stage1_42[47]}
   );
   gpc615_5 gpc505 (
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70]},
      {stage0_43[18]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[8],stage1_44[14],stage1_43[34],stage1_42[48]}
   );
   gpc615_5 gpc506 (
      {stage0_42[71], stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75]},
      {stage0_43[19]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[9],stage1_44[15],stage1_43[35],stage1_42[49]}
   );
   gpc615_5 gpc507 (
      {stage0_42[76], stage0_42[77], stage0_42[78], stage0_42[79], stage0_42[80]},
      {stage0_43[20]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[10],stage1_44[16],stage1_43[36],stage1_42[50]}
   );
   gpc615_5 gpc508 (
      {stage0_42[81], stage0_42[82], stage0_42[83], stage0_42[84], stage0_42[85]},
      {stage0_43[21]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[11],stage1_44[17],stage1_43[37],stage1_42[51]}
   );
   gpc615_5 gpc509 (
      {stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89], stage0_42[90]},
      {stage0_43[22]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[12],stage1_44[18],stage1_43[38],stage1_42[52]}
   );
   gpc615_5 gpc510 (
      {stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage0_43[23]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[13],stage1_44[19],stage1_43[39],stage1_42[53]}
   );
   gpc615_5 gpc511 (
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100]},
      {stage0_43[24]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[14],stage1_44[20],stage1_43[40],stage1_42[54]}
   );
   gpc615_5 gpc512 (
      {stage0_42[101], stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105]},
      {stage0_43[25]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[15],stage1_44[21],stage1_43[41],stage1_42[55]}
   );
   gpc615_5 gpc513 (
      {stage0_42[106], stage0_42[107], stage0_42[108], stage0_42[109], stage0_42[110]},
      {stage0_43[26]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[16],stage1_44[22],stage1_43[42],stage1_42[56]}
   );
   gpc615_5 gpc514 (
      {stage0_42[111], stage0_42[112], stage0_42[113], stage0_42[114], stage0_42[115]},
      {stage0_43[27]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[17],stage1_44[23],stage1_43[43],stage1_42[57]}
   );
   gpc615_5 gpc515 (
      {stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119], stage0_42[120]},
      {stage0_43[28]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[18],stage1_44[24],stage1_43[44],stage1_42[58]}
   );
   gpc615_5 gpc516 (
      {stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage0_43[29]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[19],stage1_44[25],stage1_43[45],stage1_42[59]}
   );
   gpc606_5 gpc517 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[17],stage1_45[20],stage1_44[26],stage1_43[46]}
   );
   gpc606_5 gpc518 (
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[18],stage1_45[21],stage1_44[27],stage1_43[47]}
   );
   gpc606_5 gpc519 (
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[19],stage1_45[22],stage1_44[28],stage1_43[48]}
   );
   gpc606_5 gpc520 (
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[20],stage1_45[23],stage1_44[29],stage1_43[49]}
   );
   gpc606_5 gpc521 (
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[21],stage1_45[24],stage1_44[30],stage1_43[50]}
   );
   gpc606_5 gpc522 (
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[22],stage1_45[25],stage1_44[31],stage1_43[51]}
   );
   gpc606_5 gpc523 (
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[23],stage1_45[26],stage1_44[32],stage1_43[52]}
   );
   gpc606_5 gpc524 (
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[24],stage1_45[27],stage1_44[33],stage1_43[53]}
   );
   gpc606_5 gpc525 (
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[8],stage1_46[25],stage1_45[28],stage1_44[34]}
   );
   gpc606_5 gpc526 (
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[9],stage1_46[26],stage1_45[29],stage1_44[35]}
   );
   gpc606_5 gpc527 (
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[10],stage1_46[27],stage1_45[30],stage1_44[36]}
   );
   gpc606_5 gpc528 (
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[11],stage1_46[28],stage1_45[31],stage1_44[37]}
   );
   gpc606_5 gpc529 (
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[12],stage1_46[29],stage1_45[32],stage1_44[38]}
   );
   gpc606_5 gpc530 (
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[13],stage1_46[30],stage1_45[33],stage1_44[39]}
   );
   gpc606_5 gpc531 (
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[14],stage1_46[31],stage1_45[34],stage1_44[40]}
   );
   gpc606_5 gpc532 (
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[15],stage1_46[32],stage1_45[35],stage1_44[41]}
   );
   gpc615_5 gpc533 (
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154]},
      {stage0_45[48]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[16],stage1_46[33],stage1_45[36],stage1_44[42]}
   );
   gpc615_5 gpc534 (
      {stage0_44[155], stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159]},
      {stage0_45[49]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[17],stage1_46[34],stage1_45[37],stage1_44[43]}
   );
   gpc606_5 gpc535 (
      {stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53], stage0_45[54], stage0_45[55]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[10],stage1_47[18],stage1_46[35],stage1_45[38]}
   );
   gpc615_5 gpc536 (
      {stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59], stage0_45[60]},
      {stage0_46[60]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[11],stage1_47[19],stage1_46[36],stage1_45[39]}
   );
   gpc615_5 gpc537 (
      {stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage0_46[61]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[12],stage1_47[20],stage1_46[37],stage1_45[40]}
   );
   gpc615_5 gpc538 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70]},
      {stage0_46[62]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[13],stage1_47[21],stage1_46[38],stage1_45[41]}
   );
   gpc615_5 gpc539 (
      {stage0_45[71], stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75]},
      {stage0_46[63]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[14],stage1_47[22],stage1_46[39],stage1_45[42]}
   );
   gpc615_5 gpc540 (
      {stage0_45[76], stage0_45[77], stage0_45[78], stage0_45[79], stage0_45[80]},
      {stage0_46[64]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[15],stage1_47[23],stage1_46[40],stage1_45[43]}
   );
   gpc615_5 gpc541 (
      {stage0_45[81], stage0_45[82], stage0_45[83], stage0_45[84], stage0_45[85]},
      {stage0_46[65]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[16],stage1_47[24],stage1_46[41],stage1_45[44]}
   );
   gpc615_5 gpc542 (
      {stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89], stage0_45[90]},
      {stage0_46[66]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[17],stage1_47[25],stage1_46[42],stage1_45[45]}
   );
   gpc615_5 gpc543 (
      {stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_46[67]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[18],stage1_47[26],stage1_46[43],stage1_45[46]}
   );
   gpc615_5 gpc544 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100]},
      {stage0_46[68]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[19],stage1_47[27],stage1_46[44],stage1_45[47]}
   );
   gpc615_5 gpc545 (
      {stage0_45[101], stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105]},
      {stage0_46[69]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[20],stage1_47[28],stage1_46[45],stage1_45[48]}
   );
   gpc615_5 gpc546 (
      {stage0_45[106], stage0_45[107], stage0_45[108], stage0_45[109], stage0_45[110]},
      {stage0_46[70]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[21],stage1_47[29],stage1_46[46],stage1_45[49]}
   );
   gpc615_5 gpc547 (
      {stage0_45[111], stage0_45[112], stage0_45[113], stage0_45[114], stage0_45[115]},
      {stage0_46[71]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[22],stage1_47[30],stage1_46[47],stage1_45[50]}
   );
   gpc615_5 gpc548 (
      {stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119], stage0_45[120]},
      {stage0_46[72]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[23],stage1_47[31],stage1_46[48],stage1_45[51]}
   );
   gpc117_4 gpc549 (
      {stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77], stage0_46[78], stage0_46[79]},
      {stage0_47[84]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[24],stage1_47[32],stage1_46[49]}
   );
   gpc117_4 gpc550 (
      {stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83], stage0_46[84], stage0_46[85], stage0_46[86]},
      {stage0_47[85]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[25],stage1_47[33],stage1_46[50]}
   );
   gpc117_4 gpc551 (
      {stage0_46[87], stage0_46[88], stage0_46[89], stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93]},
      {stage0_47[86]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[26],stage1_47[34],stage1_46[51]}
   );
   gpc117_4 gpc552 (
      {stage0_46[94], stage0_46[95], stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100]},
      {stage0_47[87]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[27],stage1_47[35],stage1_46[52]}
   );
   gpc117_4 gpc553 (
      {stage0_46[101], stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage0_47[88]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[28],stage1_47[36],stage1_46[53]}
   );
   gpc117_4 gpc554 (
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113], stage0_46[114]},
      {stage0_47[89]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[29],stage1_47[37],stage1_46[54]}
   );
   gpc117_4 gpc555 (
      {stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119], stage0_46[120], stage0_46[121]},
      {stage0_47[90]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[30],stage1_47[38],stage1_46[55]}
   );
   gpc606_5 gpc556 (
      {stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125], stage0_46[126], stage0_46[127]},
      {stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11], stage0_48[12]},
      {stage1_50[0],stage1_49[21],stage1_48[31],stage1_47[39],stage1_46[56]}
   );
   gpc606_5 gpc557 (
      {stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131], stage0_46[132], stage0_46[133]},
      {stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17], stage0_48[18]},
      {stage1_50[1],stage1_49[22],stage1_48[32],stage1_47[40],stage1_46[57]}
   );
   gpc606_5 gpc558 (
      {stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137], stage0_46[138], stage0_46[139]},
      {stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23], stage0_48[24]},
      {stage1_50[2],stage1_49[23],stage1_48[33],stage1_47[41],stage1_46[58]}
   );
   gpc606_5 gpc559 (
      {stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143], stage0_46[144], stage0_46[145]},
      {stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29], stage0_48[30]},
      {stage1_50[3],stage1_49[24],stage1_48[34],stage1_47[42],stage1_46[59]}
   );
   gpc615_5 gpc560 (
      {stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149], stage0_46[150]},
      {stage0_47[91]},
      {stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35], stage0_48[36]},
      {stage1_50[4],stage1_49[25],stage1_48[35],stage1_47[43],stage1_46[60]}
   );
   gpc615_5 gpc561 (
      {stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage0_47[92]},
      {stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41], stage0_48[42]},
      {stage1_50[5],stage1_49[26],stage1_48[36],stage1_47[44],stage1_46[61]}
   );
   gpc615_5 gpc562 (
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160]},
      {stage0_47[93]},
      {stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47], stage0_48[48]},
      {stage1_50[6],stage1_49[27],stage1_48[37],stage1_47[45],stage1_46[62]}
   );
   gpc606_5 gpc563 (
      {stage0_47[94], stage0_47[95], stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[7],stage1_49[28],stage1_48[38],stage1_47[46]}
   );
   gpc606_5 gpc564 (
      {stage0_47[100], stage0_47[101], stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[8],stage1_49[29],stage1_48[39],stage1_47[47]}
   );
   gpc606_5 gpc565 (
      {stage0_47[106], stage0_47[107], stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[9],stage1_49[30],stage1_48[40],stage1_47[48]}
   );
   gpc606_5 gpc566 (
      {stage0_47[112], stage0_47[113], stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[10],stage1_49[31],stage1_48[41],stage1_47[49]}
   );
   gpc606_5 gpc567 (
      {stage0_47[118], stage0_47[119], stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[11],stage1_49[32],stage1_48[42],stage1_47[50]}
   );
   gpc606_5 gpc568 (
      {stage0_47[124], stage0_47[125], stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[12],stage1_49[33],stage1_48[43],stage1_47[51]}
   );
   gpc606_5 gpc569 (
      {stage0_47[130], stage0_47[131], stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[13],stage1_49[34],stage1_48[44],stage1_47[52]}
   );
   gpc606_5 gpc570 (
      {stage0_47[136], stage0_47[137], stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[14],stage1_49[35],stage1_48[45],stage1_47[53]}
   );
   gpc615_5 gpc571 (
      {stage0_47[142], stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146]},
      {stage0_48[49]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[15],stage1_49[36],stage1_48[46],stage1_47[54]}
   );
   gpc615_5 gpc572 (
      {stage0_47[147], stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151]},
      {stage0_48[50]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[16],stage1_49[37],stage1_48[47],stage1_47[55]}
   );
   gpc615_5 gpc573 (
      {stage0_47[152], stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156]},
      {stage0_48[51]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[17],stage1_49[38],stage1_48[48],stage1_47[56]}
   );
   gpc615_5 gpc574 (
      {stage0_47[157], stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161]},
      {stage0_48[52]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[18],stage1_49[39],stage1_48[49],stage1_47[57]}
   );
   gpc606_5 gpc575 (
      {stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[12],stage1_50[19],stage1_49[40],stage1_48[50]}
   );
   gpc606_5 gpc576 (
      {stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[13],stage1_50[20],stage1_49[41],stage1_48[51]}
   );
   gpc606_5 gpc577 (
      {stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[14],stage1_50[21],stage1_49[42],stage1_48[52]}
   );
   gpc615_5 gpc578 (
      {stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage0_49[72]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[15],stage1_50[22],stage1_49[43],stage1_48[53]}
   );
   gpc615_5 gpc579 (
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80]},
      {stage0_49[73]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[16],stage1_50[23],stage1_49[44],stage1_48[54]}
   );
   gpc615_5 gpc580 (
      {stage0_48[81], stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85]},
      {stage0_49[74]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[17],stage1_50[24],stage1_49[45],stage1_48[55]}
   );
   gpc615_5 gpc581 (
      {stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89], stage0_48[90]},
      {stage0_49[75]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[18],stage1_50[25],stage1_49[46],stage1_48[56]}
   );
   gpc615_5 gpc582 (
      {stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage0_49[76]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[19],stage1_50[26],stage1_49[47],stage1_48[57]}
   );
   gpc615_5 gpc583 (
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100]},
      {stage0_49[77]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[20],stage1_50[27],stage1_49[48],stage1_48[58]}
   );
   gpc615_5 gpc584 (
      {stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage0_49[78]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[21],stage1_50[28],stage1_49[49],stage1_48[59]}
   );
   gpc615_5 gpc585 (
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110]},
      {stage0_49[79]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[22],stage1_50[29],stage1_49[50],stage1_48[60]}
   );
   gpc615_5 gpc586 (
      {stage0_48[111], stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115]},
      {stage0_49[80]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[23],stage1_50[30],stage1_49[51],stage1_48[61]}
   );
   gpc615_5 gpc587 (
      {stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119], stage0_48[120]},
      {stage0_49[81]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[24],stage1_50[31],stage1_49[52],stage1_48[62]}
   );
   gpc615_5 gpc588 (
      {stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage0_49[82]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[25],stage1_50[32],stage1_49[53],stage1_48[63]}
   );
   gpc615_5 gpc589 (
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130]},
      {stage0_49[83]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[26],stage1_50[33],stage1_49[54],stage1_48[64]}
   );
   gpc615_5 gpc590 (
      {stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage0_49[84]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[27],stage1_50[34],stage1_49[55],stage1_48[65]}
   );
   gpc615_5 gpc591 (
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140]},
      {stage0_49[85]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[28],stage1_50[35],stage1_49[56],stage1_48[66]}
   );
   gpc615_5 gpc592 (
      {stage0_48[141], stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145]},
      {stage0_49[86]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[29],stage1_50[36],stage1_49[57],stage1_48[67]}
   );
   gpc615_5 gpc593 (
      {stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149], stage0_48[150]},
      {stage0_49[87]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[30],stage1_50[37],stage1_49[58],stage1_48[68]}
   );
   gpc615_5 gpc594 (
      {stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage0_49[88]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[31],stage1_50[38],stage1_49[59],stage1_48[69]}
   );
   gpc615_5 gpc595 (
      {stage0_48[156], stage0_48[157], stage0_48[158], stage0_48[159], stage0_48[160]},
      {stage0_49[89]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[32],stage1_50[39],stage1_49[60],stage1_48[70]}
   );
   gpc606_5 gpc596 (
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[21],stage1_51[33],stage1_50[40],stage1_49[61]}
   );
   gpc606_5 gpc597 (
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[22],stage1_51[34],stage1_50[41],stage1_49[62]}
   );
   gpc615_5 gpc598 (
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_50[126]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[23],stage1_51[35],stage1_50[42],stage1_49[63]}
   );
   gpc615_5 gpc599 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111]},
      {stage0_50[127]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[24],stage1_51[36],stage1_50[43],stage1_49[64]}
   );
   gpc615_5 gpc600 (
      {stage0_49[112], stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116]},
      {stage0_50[128]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[25],stage1_51[37],stage1_50[44],stage1_49[65]}
   );
   gpc615_5 gpc601 (
      {stage0_49[117], stage0_49[118], stage0_49[119], stage0_49[120], stage0_49[121]},
      {stage0_50[129]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[26],stage1_51[38],stage1_50[45],stage1_49[66]}
   );
   gpc615_5 gpc602 (
      {stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125], stage0_49[126]},
      {stage0_50[130]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[27],stage1_51[39],stage1_50[46],stage1_49[67]}
   );
   gpc615_5 gpc603 (
      {stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage0_50[131]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[28],stage1_51[40],stage1_50[47],stage1_49[68]}
   );
   gpc615_5 gpc604 (
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136]},
      {stage0_50[132]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[29],stage1_51[41],stage1_50[48],stage1_49[69]}
   );
   gpc615_5 gpc605 (
      {stage0_49[137], stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141]},
      {stage0_50[133]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[30],stage1_51[42],stage1_50[49],stage1_49[70]}
   );
   gpc615_5 gpc606 (
      {stage0_49[142], stage0_49[143], stage0_49[144], stage0_49[145], stage0_49[146]},
      {stage0_50[134]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[31],stage1_51[43],stage1_50[50],stage1_49[71]}
   );
   gpc606_5 gpc607 (
      {stage0_50[135], stage0_50[136], stage0_50[137], stage0_50[138], stage0_50[139], stage0_50[140]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[11],stage1_52[32],stage1_51[44],stage1_50[51]}
   );
   gpc606_5 gpc608 (
      {stage0_50[141], stage0_50[142], stage0_50[143], stage0_50[144], stage0_50[145], stage0_50[146]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[12],stage1_52[33],stage1_51[45],stage1_50[52]}
   );
   gpc606_5 gpc609 (
      {stage0_50[147], stage0_50[148], stage0_50[149], stage0_50[150], stage0_50[151], stage0_50[152]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[13],stage1_52[34],stage1_51[46],stage1_50[53]}
   );
   gpc606_5 gpc610 (
      {stage0_50[153], stage0_50[154], stage0_50[155], stage0_50[156], stage0_50[157], stage0_50[158]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[14],stage1_52[35],stage1_51[47],stage1_50[54]}
   );
   gpc606_5 gpc611 (
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[15],stage1_52[36],stage1_51[48]}
   );
   gpc606_5 gpc612 (
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[16],stage1_52[37],stage1_51[49]}
   );
   gpc606_5 gpc613 (
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[17],stage1_52[38],stage1_51[50]}
   );
   gpc606_5 gpc614 (
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[18],stage1_52[39],stage1_51[51]}
   );
   gpc606_5 gpc615 (
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[19],stage1_52[40],stage1_51[52]}
   );
   gpc606_5 gpc616 (
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[20],stage1_52[41],stage1_51[53]}
   );
   gpc606_5 gpc617 (
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[10],stage1_53[21],stage1_52[42],stage1_51[54]}
   );
   gpc606_5 gpc618 (
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[11],stage1_53[22],stage1_52[43],stage1_51[55]}
   );
   gpc606_5 gpc619 (
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[12],stage1_53[23],stage1_52[44],stage1_51[56]}
   );
   gpc606_5 gpc620 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[13],stage1_53[24],stage1_52[45],stage1_51[57]}
   );
   gpc606_5 gpc621 (
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[10],stage1_54[14],stage1_53[25],stage1_52[46]}
   );
   gpc606_5 gpc622 (
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[11],stage1_54[15],stage1_53[26],stage1_52[47]}
   );
   gpc606_5 gpc623 (
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[12],stage1_54[16],stage1_53[27],stage1_52[48]}
   );
   gpc606_5 gpc624 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[13],stage1_54[17],stage1_53[28],stage1_52[49]}
   );
   gpc606_5 gpc625 (
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[14],stage1_54[18],stage1_53[29],stage1_52[50]}
   );
   gpc606_5 gpc626 (
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[15],stage1_54[19],stage1_53[30],stage1_52[51]}
   );
   gpc606_5 gpc627 (
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[16],stage1_54[20],stage1_53[31],stage1_52[52]}
   );
   gpc606_5 gpc628 (
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[17],stage1_54[21],stage1_53[32],stage1_52[53]}
   );
   gpc606_5 gpc629 (
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[18],stage1_54[22],stage1_53[33],stage1_52[54]}
   );
   gpc606_5 gpc630 (
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[19],stage1_54[23],stage1_53[34],stage1_52[55]}
   );
   gpc606_5 gpc631 (
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[20],stage1_54[24],stage1_53[35],stage1_52[56]}
   );
   gpc606_5 gpc632 (
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[21],stage1_54[25],stage1_53[36],stage1_52[57]}
   );
   gpc606_5 gpc633 (
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[22],stage1_54[26],stage1_53[37],stage1_52[58]}
   );
   gpc606_5 gpc634 (
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[23],stage1_54[27],stage1_53[38],stage1_52[59]}
   );
   gpc606_5 gpc635 (
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[24],stage1_54[28],stage1_53[39],stage1_52[60]}
   );
   gpc606_5 gpc636 (
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[25],stage1_54[29],stage1_53[40],stage1_52[61]}
   );
   gpc606_5 gpc637 (
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[26],stage1_54[30],stage1_53[41],stage1_52[62]}
   );
   gpc606_5 gpc638 (
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[27],stage1_54[31],stage1_53[42],stage1_52[63]}
   );
   gpc606_5 gpc639 (
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[28],stage1_54[32],stage1_53[43],stage1_52[64]}
   );
   gpc615_5 gpc640 (
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142]},
      {stage0_53[60]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[29],stage1_54[33],stage1_53[44],stage1_52[65]}
   );
   gpc615_5 gpc641 (
      {stage0_52[143], stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147]},
      {stage0_53[61]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[30],stage1_54[34],stage1_53[45],stage1_52[66]}
   );
   gpc615_5 gpc642 (
      {stage0_52[148], stage0_52[149], stage0_52[150], stage0_52[151], stage0_52[152]},
      {stage0_53[62]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[31],stage1_54[35],stage1_53[46],stage1_52[67]}
   );
   gpc606_5 gpc643 (
      {stage0_53[63], stage0_53[64], stage0_53[65], stage0_53[66], stage0_53[67], stage0_53[68]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[22],stage1_55[32],stage1_54[36],stage1_53[47]}
   );
   gpc606_5 gpc644 (
      {stage0_53[69], stage0_53[70], stage0_53[71], stage0_53[72], stage0_53[73], stage0_53[74]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[23],stage1_55[33],stage1_54[37],stage1_53[48]}
   );
   gpc606_5 gpc645 (
      {stage0_53[75], stage0_53[76], stage0_53[77], stage0_53[78], stage0_53[79], stage0_53[80]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[24],stage1_55[34],stage1_54[38],stage1_53[49]}
   );
   gpc606_5 gpc646 (
      {stage0_53[81], stage0_53[82], stage0_53[83], stage0_53[84], stage0_53[85], stage0_53[86]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[25],stage1_55[35],stage1_54[39],stage1_53[50]}
   );
   gpc606_5 gpc647 (
      {stage0_53[87], stage0_53[88], stage0_53[89], stage0_53[90], stage0_53[91], stage0_53[92]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[26],stage1_55[36],stage1_54[40],stage1_53[51]}
   );
   gpc606_5 gpc648 (
      {stage0_53[93], stage0_53[94], stage0_53[95], stage0_53[96], stage0_53[97], stage0_53[98]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[27],stage1_55[37],stage1_54[41],stage1_53[52]}
   );
   gpc606_5 gpc649 (
      {stage0_53[99], stage0_53[100], stage0_53[101], stage0_53[102], stage0_53[103], stage0_53[104]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[28],stage1_55[38],stage1_54[42],stage1_53[53]}
   );
   gpc606_5 gpc650 (
      {stage0_53[105], stage0_53[106], stage0_53[107], stage0_53[108], stage0_53[109], stage0_53[110]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[29],stage1_55[39],stage1_54[43],stage1_53[54]}
   );
   gpc606_5 gpc651 (
      {stage0_53[111], stage0_53[112], stage0_53[113], stage0_53[114], stage0_53[115], stage0_53[116]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[30],stage1_55[40],stage1_54[44],stage1_53[55]}
   );
   gpc606_5 gpc652 (
      {stage0_53[117], stage0_53[118], stage0_53[119], stage0_53[120], stage0_53[121], stage0_53[122]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[31],stage1_55[41],stage1_54[45],stage1_53[56]}
   );
   gpc606_5 gpc653 (
      {stage0_53[123], stage0_53[124], stage0_53[125], stage0_53[126], stage0_53[127], stage0_53[128]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[32],stage1_55[42],stage1_54[46],stage1_53[57]}
   );
   gpc606_5 gpc654 (
      {stage0_53[129], stage0_53[130], stage0_53[131], stage0_53[132], stage0_53[133], stage0_53[134]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[33],stage1_55[43],stage1_54[47],stage1_53[58]}
   );
   gpc606_5 gpc655 (
      {stage0_53[135], stage0_53[136], stage0_53[137], stage0_53[138], stage0_53[139], stage0_53[140]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[34],stage1_55[44],stage1_54[48],stage1_53[59]}
   );
   gpc606_5 gpc656 (
      {stage0_53[141], stage0_53[142], stage0_53[143], stage0_53[144], stage0_53[145], stage0_53[146]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[35],stage1_55[45],stage1_54[49],stage1_53[60]}
   );
   gpc606_5 gpc657 (
      {stage0_53[147], stage0_53[148], stage0_53[149], stage0_53[150], stage0_53[151], stage0_53[152]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[36],stage1_55[46],stage1_54[50],stage1_53[61]}
   );
   gpc606_5 gpc658 (
      {stage0_53[153], stage0_53[154], stage0_53[155], stage0_53[156], stage0_53[157], stage0_53[158]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[37],stage1_55[47],stage1_54[51],stage1_53[62]}
   );
   gpc615_5 gpc659 (
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136]},
      {stage0_55[96]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[16],stage1_56[38],stage1_55[48],stage1_54[52]}
   );
   gpc615_5 gpc660 (
      {stage0_54[137], stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141]},
      {stage0_55[97]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[17],stage1_56[39],stage1_55[49],stage1_54[53]}
   );
   gpc615_5 gpc661 (
      {stage0_54[142], stage0_54[143], stage0_54[144], stage0_54[145], stage0_54[146]},
      {stage0_55[98]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[18],stage1_56[40],stage1_55[50],stage1_54[54]}
   );
   gpc615_5 gpc662 (
      {stage0_54[147], stage0_54[148], stage0_54[149], stage0_54[150], stage0_54[151]},
      {stage0_55[99]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[19],stage1_56[41],stage1_55[51],stage1_54[55]}
   );
   gpc615_5 gpc663 (
      {stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155], stage0_54[156]},
      {stage0_55[100]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[20],stage1_56[42],stage1_55[52],stage1_54[56]}
   );
   gpc615_5 gpc664 (
      {stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage0_55[101]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[21],stage1_56[43],stage1_55[53],stage1_54[57]}
   );
   gpc615_5 gpc665 (
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106]},
      {stage0_56[36]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[22],stage1_56[44],stage1_55[54]}
   );
   gpc615_5 gpc666 (
      {stage0_55[107], stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111]},
      {stage0_56[37]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[23],stage1_56[45],stage1_55[55]}
   );
   gpc615_5 gpc667 (
      {stage0_55[112], stage0_55[113], stage0_55[114], stage0_55[115], stage0_55[116]},
      {stage0_56[38]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[24],stage1_56[46],stage1_55[56]}
   );
   gpc615_5 gpc668 (
      {stage0_55[117], stage0_55[118], stage0_55[119], stage0_55[120], stage0_55[121]},
      {stage0_56[39]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[25],stage1_56[47],stage1_55[57]}
   );
   gpc606_5 gpc669 (
      {stage0_56[40], stage0_56[41], stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[4],stage1_58[10],stage1_57[26],stage1_56[48]}
   );
   gpc606_5 gpc670 (
      {stage0_56[46], stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[5],stage1_58[11],stage1_57[27],stage1_56[49]}
   );
   gpc606_5 gpc671 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[6],stage1_58[12],stage1_57[28],stage1_56[50]}
   );
   gpc606_5 gpc672 (
      {stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[7],stage1_58[13],stage1_57[29],stage1_56[51]}
   );
   gpc606_5 gpc673 (
      {stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[8],stage1_58[14],stage1_57[30],stage1_56[52]}
   );
   gpc606_5 gpc674 (
      {stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[9],stage1_58[15],stage1_57[31],stage1_56[53]}
   );
   gpc606_5 gpc675 (
      {stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[10],stage1_58[16],stage1_57[32],stage1_56[54]}
   );
   gpc606_5 gpc676 (
      {stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[11],stage1_58[17],stage1_57[33],stage1_56[55]}
   );
   gpc606_5 gpc677 (
      {stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[12],stage1_58[18],stage1_57[34],stage1_56[56]}
   );
   gpc606_5 gpc678 (
      {stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[13],stage1_58[19],stage1_57[35],stage1_56[57]}
   );
   gpc606_5 gpc679 (
      {stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[14],stage1_58[20],stage1_57[36],stage1_56[58]}
   );
   gpc606_5 gpc680 (
      {stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[15],stage1_58[21],stage1_57[37],stage1_56[59]}
   );
   gpc606_5 gpc681 (
      {stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[16],stage1_58[22],stage1_57[38],stage1_56[60]}
   );
   gpc606_5 gpc682 (
      {stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[17],stage1_58[23],stage1_57[39],stage1_56[61]}
   );
   gpc606_5 gpc683 (
      {stage0_56[124], stage0_56[125], stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[18],stage1_58[24],stage1_57[40],stage1_56[62]}
   );
   gpc606_5 gpc684 (
      {stage0_56[130], stage0_56[131], stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[19],stage1_58[25],stage1_57[41],stage1_56[63]}
   );
   gpc606_5 gpc685 (
      {stage0_56[136], stage0_56[137], stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[20],stage1_58[26],stage1_57[42],stage1_56[64]}
   );
   gpc606_5 gpc686 (
      {stage0_56[142], stage0_56[143], stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[21],stage1_58[27],stage1_57[43],stage1_56[65]}
   );
   gpc606_5 gpc687 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[18],stage1_59[22],stage1_58[28],stage1_57[44]}
   );
   gpc606_5 gpc688 (
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[19],stage1_59[23],stage1_58[29],stage1_57[45]}
   );
   gpc606_5 gpc689 (
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[20],stage1_59[24],stage1_58[30],stage1_57[46]}
   );
   gpc606_5 gpc690 (
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[21],stage1_59[25],stage1_58[31],stage1_57[47]}
   );
   gpc606_5 gpc691 (
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[22],stage1_59[26],stage1_58[32],stage1_57[48]}
   );
   gpc606_5 gpc692 (
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[23],stage1_59[27],stage1_58[33],stage1_57[49]}
   );
   gpc606_5 gpc693 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[24],stage1_59[28],stage1_58[34],stage1_57[50]}
   );
   gpc606_5 gpc694 (
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[25],stage1_59[29],stage1_58[35],stage1_57[51]}
   );
   gpc606_5 gpc695 (
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[26],stage1_59[30],stage1_58[36],stage1_57[52]}
   );
   gpc606_5 gpc696 (
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[27],stage1_59[31],stage1_58[37],stage1_57[53]}
   );
   gpc606_5 gpc697 (
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[28],stage1_59[32],stage1_58[38],stage1_57[54]}
   );
   gpc606_5 gpc698 (
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[29],stage1_59[33],stage1_58[39],stage1_57[55]}
   );
   gpc606_5 gpc699 (
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[30],stage1_59[34],stage1_58[40],stage1_57[56]}
   );
   gpc606_5 gpc700 (
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[31],stage1_59[35],stage1_58[41],stage1_57[57]}
   );
   gpc606_5 gpc701 (
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[32],stage1_59[36],stage1_58[42],stage1_57[58]}
   );
   gpc606_5 gpc702 (
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[33],stage1_59[37],stage1_58[43],stage1_57[59]}
   );
   gpc606_5 gpc703 (
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[34],stage1_59[38],stage1_58[44],stage1_57[60]}
   );
   gpc606_5 gpc704 (
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[35],stage1_59[39],stage1_58[45],stage1_57[61]}
   );
   gpc606_5 gpc705 (
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[36],stage1_59[40],stage1_58[46],stage1_57[62]}
   );
   gpc606_5 gpc706 (
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[37],stage1_59[41],stage1_58[47],stage1_57[63]}
   );
   gpc606_5 gpc707 (
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[38],stage1_59[42],stage1_58[48],stage1_57[64]}
   );
   gpc606_5 gpc708 (
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[39],stage1_59[43],stage1_58[49],stage1_57[65]}
   );
   gpc606_5 gpc709 (
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[22],stage1_60[40],stage1_59[44],stage1_58[50]}
   );
   gpc606_5 gpc710 (
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[23],stage1_60[41],stage1_59[45],stage1_58[51]}
   );
   gpc606_5 gpc711 (
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[24],stage1_60[42],stage1_59[46],stage1_58[52]}
   );
   gpc606_5 gpc712 (
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[25],stage1_60[43],stage1_59[47],stage1_58[53]}
   );
   gpc606_5 gpc713 (
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[26],stage1_60[44],stage1_59[48],stage1_58[54]}
   );
   gpc606_5 gpc714 (
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[27],stage1_60[45],stage1_59[49],stage1_58[55]}
   );
   gpc606_5 gpc715 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[0],stage1_62[6],stage1_61[28],stage1_60[46]}
   );
   gpc606_5 gpc716 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[1],stage1_62[7],stage1_61[29],stage1_60[47]}
   );
   gpc606_5 gpc717 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[2],stage1_62[8],stage1_61[30],stage1_60[48]}
   );
   gpc606_5 gpc718 (
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[3],stage1_62[9],stage1_61[31],stage1_60[49]}
   );
   gpc606_5 gpc719 (
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[4],stage1_62[10],stage1_61[32],stage1_60[50]}
   );
   gpc606_5 gpc720 (
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[5],stage1_62[11],stage1_61[33],stage1_60[51]}
   );
   gpc606_5 gpc721 (
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[6],stage1_62[12],stage1_61[34],stage1_60[52]}
   );
   gpc606_5 gpc722 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[7],stage1_62[13],stage1_61[35],stage1_60[53]}
   );
   gpc606_5 gpc723 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[8],stage1_62[14],stage1_61[36],stage1_60[54]}
   );
   gpc606_5 gpc724 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[9],stage1_62[15],stage1_61[37],stage1_60[55]}
   );
   gpc606_5 gpc725 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[10],stage1_62[16],stage1_61[38],stage1_60[56]}
   );
   gpc606_5 gpc726 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[11],stage1_62[17],stage1_61[39],stage1_60[57]}
   );
   gpc606_5 gpc727 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[12],stage1_62[18],stage1_61[40],stage1_60[58]}
   );
   gpc606_5 gpc728 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[13],stage1_62[19],stage1_61[41],stage1_60[59]}
   );
   gpc606_5 gpc729 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[14],stage1_62[20],stage1_61[42],stage1_60[60]}
   );
   gpc606_5 gpc730 (
      {stage0_60[126], stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[15],stage1_62[21],stage1_61[43],stage1_60[61]}
   );
   gpc606_5 gpc731 (
      {stage0_60[132], stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[16],stage1_62[22],stage1_61[44],stage1_60[62]}
   );
   gpc606_5 gpc732 (
      {stage0_60[138], stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[17],stage1_62[23],stage1_61[45],stage1_60[63]}
   );
   gpc606_5 gpc733 (
      {stage0_60[144], stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[18],stage1_62[24],stage1_61[46],stage1_60[64]}
   );
   gpc606_5 gpc734 (
      {stage0_60[150], stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[19],stage1_62[25],stage1_61[47],stage1_60[65]}
   );
   gpc606_5 gpc735 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[20],stage1_62[26],stage1_61[48],stage1_60[66]}
   );
   gpc606_5 gpc736 (
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[21],stage1_63[21],stage1_62[27],stage1_61[49]}
   );
   gpc606_5 gpc737 (
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[22],stage1_63[22],stage1_62[28],stage1_61[50]}
   );
   gpc606_5 gpc738 (
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[23],stage1_63[23],stage1_62[29],stage1_61[51]}
   );
   gpc606_5 gpc739 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[24],stage1_63[24],stage1_62[30],stage1_61[52]}
   );
   gpc606_5 gpc740 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[25],stage1_63[25],stage1_62[31],stage1_61[53]}
   );
   gpc606_5 gpc741 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[26],stage1_63[26],stage1_62[32],stage1_61[54]}
   );
   gpc606_5 gpc742 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[27],stage1_63[27],stage1_62[33],stage1_61[55]}
   );
   gpc606_5 gpc743 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[28],stage1_63[28],stage1_62[34],stage1_61[56]}
   );
   gpc606_5 gpc744 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[29],stage1_63[29],stage1_62[35],stage1_61[57]}
   );
   gpc606_5 gpc745 (
      {stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58], stage0_61[59]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[30],stage1_63[30],stage1_62[36],stage1_61[58]}
   );
   gpc606_5 gpc746 (
      {stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64], stage0_61[65]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[31],stage1_63[31],stage1_62[37],stage1_61[59]}
   );
   gpc606_5 gpc747 (
      {stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70], stage0_61[71]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[32],stage1_63[32],stage1_62[38],stage1_61[60]}
   );
   gpc606_5 gpc748 (
      {stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76], stage0_61[77]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[33],stage1_63[33],stage1_62[39],stage1_61[61]}
   );
   gpc606_5 gpc749 (
      {stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82], stage0_61[83]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[34],stage1_63[34],stage1_62[40],stage1_61[62]}
   );
   gpc606_5 gpc750 (
      {stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88], stage0_61[89]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[35],stage1_63[35],stage1_62[41],stage1_61[63]}
   );
   gpc606_5 gpc751 (
      {stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94], stage0_61[95]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[36],stage1_63[36],stage1_62[42],stage1_61[64]}
   );
   gpc606_5 gpc752 (
      {stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100], stage0_61[101]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[37],stage1_63[37],stage1_62[43],stage1_61[65]}
   );
   gpc606_5 gpc753 (
      {stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106], stage0_61[107]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[38],stage1_63[38],stage1_62[44],stage1_61[66]}
   );
   gpc606_5 gpc754 (
      {stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112], stage0_61[113]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[39],stage1_63[39],stage1_62[45],stage1_61[67]}
   );
   gpc606_5 gpc755 (
      {stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118], stage0_61[119]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[40],stage1_63[40],stage1_62[46],stage1_61[68]}
   );
   gpc606_5 gpc756 (
      {stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124], stage0_61[125]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[41],stage1_63[41],stage1_62[47],stage1_61[69]}
   );
   gpc606_5 gpc757 (
      {stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130], stage0_61[131]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[42],stage1_63[42],stage1_62[48],stage1_61[70]}
   );
   gpc606_5 gpc758 (
      {stage0_61[132], stage0_61[133], stage0_61[134], stage0_61[135], stage0_61[136], stage0_61[137]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[43],stage1_63[43],stage1_62[49],stage1_61[71]}
   );
   gpc606_5 gpc759 (
      {stage0_61[138], stage0_61[139], stage0_61[140], stage0_61[141], stage0_61[142], stage0_61[143]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[44],stage1_63[44],stage1_62[50],stage1_61[72]}
   );
   gpc1_1 gpc760 (
      {stage0_2[160]},
      {stage1_2[53]}
   );
   gpc1_1 gpc761 (
      {stage0_2[161]},
      {stage1_2[54]}
   );
   gpc1_1 gpc762 (
      {stage0_3[139]},
      {stage1_3[61]}
   );
   gpc1_1 gpc763 (
      {stage0_3[140]},
      {stage1_3[62]}
   );
   gpc1_1 gpc764 (
      {stage0_3[141]},
      {stage1_3[63]}
   );
   gpc1_1 gpc765 (
      {stage0_3[142]},
      {stage1_3[64]}
   );
   gpc1_1 gpc766 (
      {stage0_3[143]},
      {stage1_3[65]}
   );
   gpc1_1 gpc767 (
      {stage0_3[144]},
      {stage1_3[66]}
   );
   gpc1_1 gpc768 (
      {stage0_3[145]},
      {stage1_3[67]}
   );
   gpc1_1 gpc769 (
      {stage0_3[146]},
      {stage1_3[68]}
   );
   gpc1_1 gpc770 (
      {stage0_3[147]},
      {stage1_3[69]}
   );
   gpc1_1 gpc771 (
      {stage0_3[148]},
      {stage1_3[70]}
   );
   gpc1_1 gpc772 (
      {stage0_3[149]},
      {stage1_3[71]}
   );
   gpc1_1 gpc773 (
      {stage0_3[150]},
      {stage1_3[72]}
   );
   gpc1_1 gpc774 (
      {stage0_3[151]},
      {stage1_3[73]}
   );
   gpc1_1 gpc775 (
      {stage0_3[152]},
      {stage1_3[74]}
   );
   gpc1_1 gpc776 (
      {stage0_3[153]},
      {stage1_3[75]}
   );
   gpc1_1 gpc777 (
      {stage0_3[154]},
      {stage1_3[76]}
   );
   gpc1_1 gpc778 (
      {stage0_3[155]},
      {stage1_3[77]}
   );
   gpc1_1 gpc779 (
      {stage0_3[156]},
      {stage1_3[78]}
   );
   gpc1_1 gpc780 (
      {stage0_3[157]},
      {stage1_3[79]}
   );
   gpc1_1 gpc781 (
      {stage0_3[158]},
      {stage1_3[80]}
   );
   gpc1_1 gpc782 (
      {stage0_3[159]},
      {stage1_3[81]}
   );
   gpc1_1 gpc783 (
      {stage0_3[160]},
      {stage1_3[82]}
   );
   gpc1_1 gpc784 (
      {stage0_3[161]},
      {stage1_3[83]}
   );
   gpc1_1 gpc785 (
      {stage0_4[158]},
      {stage1_4[79]}
   );
   gpc1_1 gpc786 (
      {stage0_4[159]},
      {stage1_4[80]}
   );
   gpc1_1 gpc787 (
      {stage0_4[160]},
      {stage1_4[81]}
   );
   gpc1_1 gpc788 (
      {stage0_4[161]},
      {stage1_4[82]}
   );
   gpc1_1 gpc789 (
      {stage0_5[102]},
      {stage1_5[55]}
   );
   gpc1_1 gpc790 (
      {stage0_5[103]},
      {stage1_5[56]}
   );
   gpc1_1 gpc791 (
      {stage0_5[104]},
      {stage1_5[57]}
   );
   gpc1_1 gpc792 (
      {stage0_5[105]},
      {stage1_5[58]}
   );
   gpc1_1 gpc793 (
      {stage0_5[106]},
      {stage1_5[59]}
   );
   gpc1_1 gpc794 (
      {stage0_5[107]},
      {stage1_5[60]}
   );
   gpc1_1 gpc795 (
      {stage0_5[108]},
      {stage1_5[61]}
   );
   gpc1_1 gpc796 (
      {stage0_5[109]},
      {stage1_5[62]}
   );
   gpc1_1 gpc797 (
      {stage0_5[110]},
      {stage1_5[63]}
   );
   gpc1_1 gpc798 (
      {stage0_5[111]},
      {stage1_5[64]}
   );
   gpc1_1 gpc799 (
      {stage0_5[112]},
      {stage1_5[65]}
   );
   gpc1_1 gpc800 (
      {stage0_5[113]},
      {stage1_5[66]}
   );
   gpc1_1 gpc801 (
      {stage0_5[114]},
      {stage1_5[67]}
   );
   gpc1_1 gpc802 (
      {stage0_5[115]},
      {stage1_5[68]}
   );
   gpc1_1 gpc803 (
      {stage0_5[116]},
      {stage1_5[69]}
   );
   gpc1_1 gpc804 (
      {stage0_5[117]},
      {stage1_5[70]}
   );
   gpc1_1 gpc805 (
      {stage0_5[118]},
      {stage1_5[71]}
   );
   gpc1_1 gpc806 (
      {stage0_5[119]},
      {stage1_5[72]}
   );
   gpc1_1 gpc807 (
      {stage0_5[120]},
      {stage1_5[73]}
   );
   gpc1_1 gpc808 (
      {stage0_5[121]},
      {stage1_5[74]}
   );
   gpc1_1 gpc809 (
      {stage0_5[122]},
      {stage1_5[75]}
   );
   gpc1_1 gpc810 (
      {stage0_5[123]},
      {stage1_5[76]}
   );
   gpc1_1 gpc811 (
      {stage0_5[124]},
      {stage1_5[77]}
   );
   gpc1_1 gpc812 (
      {stage0_5[125]},
      {stage1_5[78]}
   );
   gpc1_1 gpc813 (
      {stage0_5[126]},
      {stage1_5[79]}
   );
   gpc1_1 gpc814 (
      {stage0_5[127]},
      {stage1_5[80]}
   );
   gpc1_1 gpc815 (
      {stage0_5[128]},
      {stage1_5[81]}
   );
   gpc1_1 gpc816 (
      {stage0_5[129]},
      {stage1_5[82]}
   );
   gpc1_1 gpc817 (
      {stage0_5[130]},
      {stage1_5[83]}
   );
   gpc1_1 gpc818 (
      {stage0_5[131]},
      {stage1_5[84]}
   );
   gpc1_1 gpc819 (
      {stage0_5[132]},
      {stage1_5[85]}
   );
   gpc1_1 gpc820 (
      {stage0_5[133]},
      {stage1_5[86]}
   );
   gpc1_1 gpc821 (
      {stage0_5[134]},
      {stage1_5[87]}
   );
   gpc1_1 gpc822 (
      {stage0_5[135]},
      {stage1_5[88]}
   );
   gpc1_1 gpc823 (
      {stage0_5[136]},
      {stage1_5[89]}
   );
   gpc1_1 gpc824 (
      {stage0_5[137]},
      {stage1_5[90]}
   );
   gpc1_1 gpc825 (
      {stage0_5[138]},
      {stage1_5[91]}
   );
   gpc1_1 gpc826 (
      {stage0_5[139]},
      {stage1_5[92]}
   );
   gpc1_1 gpc827 (
      {stage0_5[140]},
      {stage1_5[93]}
   );
   gpc1_1 gpc828 (
      {stage0_5[141]},
      {stage1_5[94]}
   );
   gpc1_1 gpc829 (
      {stage0_5[142]},
      {stage1_5[95]}
   );
   gpc1_1 gpc830 (
      {stage0_5[143]},
      {stage1_5[96]}
   );
   gpc1_1 gpc831 (
      {stage0_5[144]},
      {stage1_5[97]}
   );
   gpc1_1 gpc832 (
      {stage0_5[145]},
      {stage1_5[98]}
   );
   gpc1_1 gpc833 (
      {stage0_5[146]},
      {stage1_5[99]}
   );
   gpc1_1 gpc834 (
      {stage0_5[147]},
      {stage1_5[100]}
   );
   gpc1_1 gpc835 (
      {stage0_5[148]},
      {stage1_5[101]}
   );
   gpc1_1 gpc836 (
      {stage0_5[149]},
      {stage1_5[102]}
   );
   gpc1_1 gpc837 (
      {stage0_5[150]},
      {stage1_5[103]}
   );
   gpc1_1 gpc838 (
      {stage0_5[151]},
      {stage1_5[104]}
   );
   gpc1_1 gpc839 (
      {stage0_5[152]},
      {stage1_5[105]}
   );
   gpc1_1 gpc840 (
      {stage0_5[153]},
      {stage1_5[106]}
   );
   gpc1_1 gpc841 (
      {stage0_5[154]},
      {stage1_5[107]}
   );
   gpc1_1 gpc842 (
      {stage0_5[155]},
      {stage1_5[108]}
   );
   gpc1_1 gpc843 (
      {stage0_5[156]},
      {stage1_5[109]}
   );
   gpc1_1 gpc844 (
      {stage0_5[157]},
      {stage1_5[110]}
   );
   gpc1_1 gpc845 (
      {stage0_5[158]},
      {stage1_5[111]}
   );
   gpc1_1 gpc846 (
      {stage0_5[159]},
      {stage1_5[112]}
   );
   gpc1_1 gpc847 (
      {stage0_5[160]},
      {stage1_5[113]}
   );
   gpc1_1 gpc848 (
      {stage0_5[161]},
      {stage1_5[114]}
   );
   gpc1_1 gpc849 (
      {stage0_6[154]},
      {stage1_6[50]}
   );
   gpc1_1 gpc850 (
      {stage0_6[155]},
      {stage1_6[51]}
   );
   gpc1_1 gpc851 (
      {stage0_6[156]},
      {stage1_6[52]}
   );
   gpc1_1 gpc852 (
      {stage0_6[157]},
      {stage1_6[53]}
   );
   gpc1_1 gpc853 (
      {stage0_6[158]},
      {stage1_6[54]}
   );
   gpc1_1 gpc854 (
      {stage0_6[159]},
      {stage1_6[55]}
   );
   gpc1_1 gpc855 (
      {stage0_6[160]},
      {stage1_6[56]}
   );
   gpc1_1 gpc856 (
      {stage0_6[161]},
      {stage1_6[57]}
   );
   gpc1_1 gpc857 (
      {stage0_7[153]},
      {stage1_7[62]}
   );
   gpc1_1 gpc858 (
      {stage0_7[154]},
      {stage1_7[63]}
   );
   gpc1_1 gpc859 (
      {stage0_7[155]},
      {stage1_7[64]}
   );
   gpc1_1 gpc860 (
      {stage0_7[156]},
      {stage1_7[65]}
   );
   gpc1_1 gpc861 (
      {stage0_7[157]},
      {stage1_7[66]}
   );
   gpc1_1 gpc862 (
      {stage0_7[158]},
      {stage1_7[67]}
   );
   gpc1_1 gpc863 (
      {stage0_7[159]},
      {stage1_7[68]}
   );
   gpc1_1 gpc864 (
      {stage0_7[160]},
      {stage1_7[69]}
   );
   gpc1_1 gpc865 (
      {stage0_7[161]},
      {stage1_7[70]}
   );
   gpc1_1 gpc866 (
      {stage0_8[149]},
      {stage1_8[68]}
   );
   gpc1_1 gpc867 (
      {stage0_8[150]},
      {stage1_8[69]}
   );
   gpc1_1 gpc868 (
      {stage0_8[151]},
      {stage1_8[70]}
   );
   gpc1_1 gpc869 (
      {stage0_8[152]},
      {stage1_8[71]}
   );
   gpc1_1 gpc870 (
      {stage0_8[153]},
      {stage1_8[72]}
   );
   gpc1_1 gpc871 (
      {stage0_8[154]},
      {stage1_8[73]}
   );
   gpc1_1 gpc872 (
      {stage0_8[155]},
      {stage1_8[74]}
   );
   gpc1_1 gpc873 (
      {stage0_8[156]},
      {stage1_8[75]}
   );
   gpc1_1 gpc874 (
      {stage0_8[157]},
      {stage1_8[76]}
   );
   gpc1_1 gpc875 (
      {stage0_8[158]},
      {stage1_8[77]}
   );
   gpc1_1 gpc876 (
      {stage0_8[159]},
      {stage1_8[78]}
   );
   gpc1_1 gpc877 (
      {stage0_8[160]},
      {stage1_8[79]}
   );
   gpc1_1 gpc878 (
      {stage0_8[161]},
      {stage1_8[80]}
   );
   gpc1_1 gpc879 (
      {stage0_10[124]},
      {stage1_10[57]}
   );
   gpc1_1 gpc880 (
      {stage0_10[125]},
      {stage1_10[58]}
   );
   gpc1_1 gpc881 (
      {stage0_10[126]},
      {stage1_10[59]}
   );
   gpc1_1 gpc882 (
      {stage0_10[127]},
      {stage1_10[60]}
   );
   gpc1_1 gpc883 (
      {stage0_10[128]},
      {stage1_10[61]}
   );
   gpc1_1 gpc884 (
      {stage0_10[129]},
      {stage1_10[62]}
   );
   gpc1_1 gpc885 (
      {stage0_10[130]},
      {stage1_10[63]}
   );
   gpc1_1 gpc886 (
      {stage0_10[131]},
      {stage1_10[64]}
   );
   gpc1_1 gpc887 (
      {stage0_10[132]},
      {stage1_10[65]}
   );
   gpc1_1 gpc888 (
      {stage0_10[133]},
      {stage1_10[66]}
   );
   gpc1_1 gpc889 (
      {stage0_10[134]},
      {stage1_10[67]}
   );
   gpc1_1 gpc890 (
      {stage0_10[135]},
      {stage1_10[68]}
   );
   gpc1_1 gpc891 (
      {stage0_10[136]},
      {stage1_10[69]}
   );
   gpc1_1 gpc892 (
      {stage0_10[137]},
      {stage1_10[70]}
   );
   gpc1_1 gpc893 (
      {stage0_10[138]},
      {stage1_10[71]}
   );
   gpc1_1 gpc894 (
      {stage0_10[139]},
      {stage1_10[72]}
   );
   gpc1_1 gpc895 (
      {stage0_10[140]},
      {stage1_10[73]}
   );
   gpc1_1 gpc896 (
      {stage0_10[141]},
      {stage1_10[74]}
   );
   gpc1_1 gpc897 (
      {stage0_10[142]},
      {stage1_10[75]}
   );
   gpc1_1 gpc898 (
      {stage0_10[143]},
      {stage1_10[76]}
   );
   gpc1_1 gpc899 (
      {stage0_10[144]},
      {stage1_10[77]}
   );
   gpc1_1 gpc900 (
      {stage0_10[145]},
      {stage1_10[78]}
   );
   gpc1_1 gpc901 (
      {stage0_10[146]},
      {stage1_10[79]}
   );
   gpc1_1 gpc902 (
      {stage0_10[147]},
      {stage1_10[80]}
   );
   gpc1_1 gpc903 (
      {stage0_10[148]},
      {stage1_10[81]}
   );
   gpc1_1 gpc904 (
      {stage0_10[149]},
      {stage1_10[82]}
   );
   gpc1_1 gpc905 (
      {stage0_10[150]},
      {stage1_10[83]}
   );
   gpc1_1 gpc906 (
      {stage0_10[151]},
      {stage1_10[84]}
   );
   gpc1_1 gpc907 (
      {stage0_10[152]},
      {stage1_10[85]}
   );
   gpc1_1 gpc908 (
      {stage0_10[153]},
      {stage1_10[86]}
   );
   gpc1_1 gpc909 (
      {stage0_10[154]},
      {stage1_10[87]}
   );
   gpc1_1 gpc910 (
      {stage0_10[155]},
      {stage1_10[88]}
   );
   gpc1_1 gpc911 (
      {stage0_10[156]},
      {stage1_10[89]}
   );
   gpc1_1 gpc912 (
      {stage0_10[157]},
      {stage1_10[90]}
   );
   gpc1_1 gpc913 (
      {stage0_10[158]},
      {stage1_10[91]}
   );
   gpc1_1 gpc914 (
      {stage0_10[159]},
      {stage1_10[92]}
   );
   gpc1_1 gpc915 (
      {stage0_10[160]},
      {stage1_10[93]}
   );
   gpc1_1 gpc916 (
      {stage0_10[161]},
      {stage1_10[94]}
   );
   gpc1_1 gpc917 (
      {stage0_11[144]},
      {stage1_11[63]}
   );
   gpc1_1 gpc918 (
      {stage0_11[145]},
      {stage1_11[64]}
   );
   gpc1_1 gpc919 (
      {stage0_11[146]},
      {stage1_11[65]}
   );
   gpc1_1 gpc920 (
      {stage0_11[147]},
      {stage1_11[66]}
   );
   gpc1_1 gpc921 (
      {stage0_11[148]},
      {stage1_11[67]}
   );
   gpc1_1 gpc922 (
      {stage0_11[149]},
      {stage1_11[68]}
   );
   gpc1_1 gpc923 (
      {stage0_11[150]},
      {stage1_11[69]}
   );
   gpc1_1 gpc924 (
      {stage0_11[151]},
      {stage1_11[70]}
   );
   gpc1_1 gpc925 (
      {stage0_11[152]},
      {stage1_11[71]}
   );
   gpc1_1 gpc926 (
      {stage0_11[153]},
      {stage1_11[72]}
   );
   gpc1_1 gpc927 (
      {stage0_11[154]},
      {stage1_11[73]}
   );
   gpc1_1 gpc928 (
      {stage0_11[155]},
      {stage1_11[74]}
   );
   gpc1_1 gpc929 (
      {stage0_11[156]},
      {stage1_11[75]}
   );
   gpc1_1 gpc930 (
      {stage0_11[157]},
      {stage1_11[76]}
   );
   gpc1_1 gpc931 (
      {stage0_11[158]},
      {stage1_11[77]}
   );
   gpc1_1 gpc932 (
      {stage0_11[159]},
      {stage1_11[78]}
   );
   gpc1_1 gpc933 (
      {stage0_11[160]},
      {stage1_11[79]}
   );
   gpc1_1 gpc934 (
      {stage0_11[161]},
      {stage1_11[80]}
   );
   gpc1_1 gpc935 (
      {stage0_12[158]},
      {stage1_12[63]}
   );
   gpc1_1 gpc936 (
      {stage0_12[159]},
      {stage1_12[64]}
   );
   gpc1_1 gpc937 (
      {stage0_12[160]},
      {stage1_12[65]}
   );
   gpc1_1 gpc938 (
      {stage0_12[161]},
      {stage1_12[66]}
   );
   gpc1_1 gpc939 (
      {stage0_13[132]},
      {stage1_13[57]}
   );
   gpc1_1 gpc940 (
      {stage0_13[133]},
      {stage1_13[58]}
   );
   gpc1_1 gpc941 (
      {stage0_13[134]},
      {stage1_13[59]}
   );
   gpc1_1 gpc942 (
      {stage0_13[135]},
      {stage1_13[60]}
   );
   gpc1_1 gpc943 (
      {stage0_13[136]},
      {stage1_13[61]}
   );
   gpc1_1 gpc944 (
      {stage0_13[137]},
      {stage1_13[62]}
   );
   gpc1_1 gpc945 (
      {stage0_13[138]},
      {stage1_13[63]}
   );
   gpc1_1 gpc946 (
      {stage0_13[139]},
      {stage1_13[64]}
   );
   gpc1_1 gpc947 (
      {stage0_13[140]},
      {stage1_13[65]}
   );
   gpc1_1 gpc948 (
      {stage0_13[141]},
      {stage1_13[66]}
   );
   gpc1_1 gpc949 (
      {stage0_13[142]},
      {stage1_13[67]}
   );
   gpc1_1 gpc950 (
      {stage0_13[143]},
      {stage1_13[68]}
   );
   gpc1_1 gpc951 (
      {stage0_13[144]},
      {stage1_13[69]}
   );
   gpc1_1 gpc952 (
      {stage0_13[145]},
      {stage1_13[70]}
   );
   gpc1_1 gpc953 (
      {stage0_13[146]},
      {stage1_13[71]}
   );
   gpc1_1 gpc954 (
      {stage0_13[147]},
      {stage1_13[72]}
   );
   gpc1_1 gpc955 (
      {stage0_13[148]},
      {stage1_13[73]}
   );
   gpc1_1 gpc956 (
      {stage0_13[149]},
      {stage1_13[74]}
   );
   gpc1_1 gpc957 (
      {stage0_13[150]},
      {stage1_13[75]}
   );
   gpc1_1 gpc958 (
      {stage0_13[151]},
      {stage1_13[76]}
   );
   gpc1_1 gpc959 (
      {stage0_13[152]},
      {stage1_13[77]}
   );
   gpc1_1 gpc960 (
      {stage0_13[153]},
      {stage1_13[78]}
   );
   gpc1_1 gpc961 (
      {stage0_13[154]},
      {stage1_13[79]}
   );
   gpc1_1 gpc962 (
      {stage0_13[155]},
      {stage1_13[80]}
   );
   gpc1_1 gpc963 (
      {stage0_13[156]},
      {stage1_13[81]}
   );
   gpc1_1 gpc964 (
      {stage0_13[157]},
      {stage1_13[82]}
   );
   gpc1_1 gpc965 (
      {stage0_13[158]},
      {stage1_13[83]}
   );
   gpc1_1 gpc966 (
      {stage0_13[159]},
      {stage1_13[84]}
   );
   gpc1_1 gpc967 (
      {stage0_13[160]},
      {stage1_13[85]}
   );
   gpc1_1 gpc968 (
      {stage0_13[161]},
      {stage1_13[86]}
   );
   gpc1_1 gpc969 (
      {stage0_14[158]},
      {stage1_14[58]}
   );
   gpc1_1 gpc970 (
      {stage0_14[159]},
      {stage1_14[59]}
   );
   gpc1_1 gpc971 (
      {stage0_14[160]},
      {stage1_14[60]}
   );
   gpc1_1 gpc972 (
      {stage0_14[161]},
      {stage1_14[61]}
   );
   gpc1_1 gpc973 (
      {stage0_15[128]},
      {stage1_15[64]}
   );
   gpc1_1 gpc974 (
      {stage0_15[129]},
      {stage1_15[65]}
   );
   gpc1_1 gpc975 (
      {stage0_15[130]},
      {stage1_15[66]}
   );
   gpc1_1 gpc976 (
      {stage0_15[131]},
      {stage1_15[67]}
   );
   gpc1_1 gpc977 (
      {stage0_15[132]},
      {stage1_15[68]}
   );
   gpc1_1 gpc978 (
      {stage0_15[133]},
      {stage1_15[69]}
   );
   gpc1_1 gpc979 (
      {stage0_15[134]},
      {stage1_15[70]}
   );
   gpc1_1 gpc980 (
      {stage0_15[135]},
      {stage1_15[71]}
   );
   gpc1_1 gpc981 (
      {stage0_15[136]},
      {stage1_15[72]}
   );
   gpc1_1 gpc982 (
      {stage0_15[137]},
      {stage1_15[73]}
   );
   gpc1_1 gpc983 (
      {stage0_15[138]},
      {stage1_15[74]}
   );
   gpc1_1 gpc984 (
      {stage0_15[139]},
      {stage1_15[75]}
   );
   gpc1_1 gpc985 (
      {stage0_15[140]},
      {stage1_15[76]}
   );
   gpc1_1 gpc986 (
      {stage0_15[141]},
      {stage1_15[77]}
   );
   gpc1_1 gpc987 (
      {stage0_15[142]},
      {stage1_15[78]}
   );
   gpc1_1 gpc988 (
      {stage0_15[143]},
      {stage1_15[79]}
   );
   gpc1_1 gpc989 (
      {stage0_15[144]},
      {stage1_15[80]}
   );
   gpc1_1 gpc990 (
      {stage0_15[145]},
      {stage1_15[81]}
   );
   gpc1_1 gpc991 (
      {stage0_15[146]},
      {stage1_15[82]}
   );
   gpc1_1 gpc992 (
      {stage0_15[147]},
      {stage1_15[83]}
   );
   gpc1_1 gpc993 (
      {stage0_15[148]},
      {stage1_15[84]}
   );
   gpc1_1 gpc994 (
      {stage0_15[149]},
      {stage1_15[85]}
   );
   gpc1_1 gpc995 (
      {stage0_15[150]},
      {stage1_15[86]}
   );
   gpc1_1 gpc996 (
      {stage0_15[151]},
      {stage1_15[87]}
   );
   gpc1_1 gpc997 (
      {stage0_15[152]},
      {stage1_15[88]}
   );
   gpc1_1 gpc998 (
      {stage0_15[153]},
      {stage1_15[89]}
   );
   gpc1_1 gpc999 (
      {stage0_15[154]},
      {stage1_15[90]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[155]},
      {stage1_15[91]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[156]},
      {stage1_15[92]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[157]},
      {stage1_15[93]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[158]},
      {stage1_15[94]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[159]},
      {stage1_15[95]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[160]},
      {stage1_15[96]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[161]},
      {stage1_15[97]}
   );
   gpc1_1 gpc1007 (
      {stage0_16[158]},
      {stage1_16[64]}
   );
   gpc1_1 gpc1008 (
      {stage0_16[159]},
      {stage1_16[65]}
   );
   gpc1_1 gpc1009 (
      {stage0_16[160]},
      {stage1_16[66]}
   );
   gpc1_1 gpc1010 (
      {stage0_16[161]},
      {stage1_16[67]}
   );
   gpc1_1 gpc1011 (
      {stage0_17[96]},
      {stage1_17[48]}
   );
   gpc1_1 gpc1012 (
      {stage0_17[97]},
      {stage1_17[49]}
   );
   gpc1_1 gpc1013 (
      {stage0_17[98]},
      {stage1_17[50]}
   );
   gpc1_1 gpc1014 (
      {stage0_17[99]},
      {stage1_17[51]}
   );
   gpc1_1 gpc1015 (
      {stage0_17[100]},
      {stage1_17[52]}
   );
   gpc1_1 gpc1016 (
      {stage0_17[101]},
      {stage1_17[53]}
   );
   gpc1_1 gpc1017 (
      {stage0_17[102]},
      {stage1_17[54]}
   );
   gpc1_1 gpc1018 (
      {stage0_17[103]},
      {stage1_17[55]}
   );
   gpc1_1 gpc1019 (
      {stage0_17[104]},
      {stage1_17[56]}
   );
   gpc1_1 gpc1020 (
      {stage0_17[105]},
      {stage1_17[57]}
   );
   gpc1_1 gpc1021 (
      {stage0_17[106]},
      {stage1_17[58]}
   );
   gpc1_1 gpc1022 (
      {stage0_17[107]},
      {stage1_17[59]}
   );
   gpc1_1 gpc1023 (
      {stage0_17[108]},
      {stage1_17[60]}
   );
   gpc1_1 gpc1024 (
      {stage0_17[109]},
      {stage1_17[61]}
   );
   gpc1_1 gpc1025 (
      {stage0_17[110]},
      {stage1_17[62]}
   );
   gpc1_1 gpc1026 (
      {stage0_17[111]},
      {stage1_17[63]}
   );
   gpc1_1 gpc1027 (
      {stage0_17[112]},
      {stage1_17[64]}
   );
   gpc1_1 gpc1028 (
      {stage0_17[113]},
      {stage1_17[65]}
   );
   gpc1_1 gpc1029 (
      {stage0_17[114]},
      {stage1_17[66]}
   );
   gpc1_1 gpc1030 (
      {stage0_17[115]},
      {stage1_17[67]}
   );
   gpc1_1 gpc1031 (
      {stage0_17[116]},
      {stage1_17[68]}
   );
   gpc1_1 gpc1032 (
      {stage0_17[117]},
      {stage1_17[69]}
   );
   gpc1_1 gpc1033 (
      {stage0_17[118]},
      {stage1_17[70]}
   );
   gpc1_1 gpc1034 (
      {stage0_17[119]},
      {stage1_17[71]}
   );
   gpc1_1 gpc1035 (
      {stage0_17[120]},
      {stage1_17[72]}
   );
   gpc1_1 gpc1036 (
      {stage0_17[121]},
      {stage1_17[73]}
   );
   gpc1_1 gpc1037 (
      {stage0_17[122]},
      {stage1_17[74]}
   );
   gpc1_1 gpc1038 (
      {stage0_17[123]},
      {stage1_17[75]}
   );
   gpc1_1 gpc1039 (
      {stage0_17[124]},
      {stage1_17[76]}
   );
   gpc1_1 gpc1040 (
      {stage0_17[125]},
      {stage1_17[77]}
   );
   gpc1_1 gpc1041 (
      {stage0_17[126]},
      {stage1_17[78]}
   );
   gpc1_1 gpc1042 (
      {stage0_17[127]},
      {stage1_17[79]}
   );
   gpc1_1 gpc1043 (
      {stage0_17[128]},
      {stage1_17[80]}
   );
   gpc1_1 gpc1044 (
      {stage0_17[129]},
      {stage1_17[81]}
   );
   gpc1_1 gpc1045 (
      {stage0_17[130]},
      {stage1_17[82]}
   );
   gpc1_1 gpc1046 (
      {stage0_17[131]},
      {stage1_17[83]}
   );
   gpc1_1 gpc1047 (
      {stage0_17[132]},
      {stage1_17[84]}
   );
   gpc1_1 gpc1048 (
      {stage0_17[133]},
      {stage1_17[85]}
   );
   gpc1_1 gpc1049 (
      {stage0_17[134]},
      {stage1_17[86]}
   );
   gpc1_1 gpc1050 (
      {stage0_17[135]},
      {stage1_17[87]}
   );
   gpc1_1 gpc1051 (
      {stage0_17[136]},
      {stage1_17[88]}
   );
   gpc1_1 gpc1052 (
      {stage0_17[137]},
      {stage1_17[89]}
   );
   gpc1_1 gpc1053 (
      {stage0_17[138]},
      {stage1_17[90]}
   );
   gpc1_1 gpc1054 (
      {stage0_17[139]},
      {stage1_17[91]}
   );
   gpc1_1 gpc1055 (
      {stage0_17[140]},
      {stage1_17[92]}
   );
   gpc1_1 gpc1056 (
      {stage0_17[141]},
      {stage1_17[93]}
   );
   gpc1_1 gpc1057 (
      {stage0_17[142]},
      {stage1_17[94]}
   );
   gpc1_1 gpc1058 (
      {stage0_17[143]},
      {stage1_17[95]}
   );
   gpc1_1 gpc1059 (
      {stage0_17[144]},
      {stage1_17[96]}
   );
   gpc1_1 gpc1060 (
      {stage0_17[145]},
      {stage1_17[97]}
   );
   gpc1_1 gpc1061 (
      {stage0_17[146]},
      {stage1_17[98]}
   );
   gpc1_1 gpc1062 (
      {stage0_17[147]},
      {stage1_17[99]}
   );
   gpc1_1 gpc1063 (
      {stage0_17[148]},
      {stage1_17[100]}
   );
   gpc1_1 gpc1064 (
      {stage0_17[149]},
      {stage1_17[101]}
   );
   gpc1_1 gpc1065 (
      {stage0_17[150]},
      {stage1_17[102]}
   );
   gpc1_1 gpc1066 (
      {stage0_17[151]},
      {stage1_17[103]}
   );
   gpc1_1 gpc1067 (
      {stage0_17[152]},
      {stage1_17[104]}
   );
   gpc1_1 gpc1068 (
      {stage0_17[153]},
      {stage1_17[105]}
   );
   gpc1_1 gpc1069 (
      {stage0_17[154]},
      {stage1_17[106]}
   );
   gpc1_1 gpc1070 (
      {stage0_17[155]},
      {stage1_17[107]}
   );
   gpc1_1 gpc1071 (
      {stage0_17[156]},
      {stage1_17[108]}
   );
   gpc1_1 gpc1072 (
      {stage0_17[157]},
      {stage1_17[109]}
   );
   gpc1_1 gpc1073 (
      {stage0_17[158]},
      {stage1_17[110]}
   );
   gpc1_1 gpc1074 (
      {stage0_17[159]},
      {stage1_17[111]}
   );
   gpc1_1 gpc1075 (
      {stage0_17[160]},
      {stage1_17[112]}
   );
   gpc1_1 gpc1076 (
      {stage0_17[161]},
      {stage1_17[113]}
   );
   gpc1_1 gpc1077 (
      {stage0_18[151]},
      {stage1_18[52]}
   );
   gpc1_1 gpc1078 (
      {stage0_18[152]},
      {stage1_18[53]}
   );
   gpc1_1 gpc1079 (
      {stage0_18[153]},
      {stage1_18[54]}
   );
   gpc1_1 gpc1080 (
      {stage0_18[154]},
      {stage1_18[55]}
   );
   gpc1_1 gpc1081 (
      {stage0_18[155]},
      {stage1_18[56]}
   );
   gpc1_1 gpc1082 (
      {stage0_18[156]},
      {stage1_18[57]}
   );
   gpc1_1 gpc1083 (
      {stage0_18[157]},
      {stage1_18[58]}
   );
   gpc1_1 gpc1084 (
      {stage0_18[158]},
      {stage1_18[59]}
   );
   gpc1_1 gpc1085 (
      {stage0_18[159]},
      {stage1_18[60]}
   );
   gpc1_1 gpc1086 (
      {stage0_18[160]},
      {stage1_18[61]}
   );
   gpc1_1 gpc1087 (
      {stage0_18[161]},
      {stage1_18[62]}
   );
   gpc1_1 gpc1088 (
      {stage0_19[156]},
      {stage1_19[65]}
   );
   gpc1_1 gpc1089 (
      {stage0_19[157]},
      {stage1_19[66]}
   );
   gpc1_1 gpc1090 (
      {stage0_19[158]},
      {stage1_19[67]}
   );
   gpc1_1 gpc1091 (
      {stage0_19[159]},
      {stage1_19[68]}
   );
   gpc1_1 gpc1092 (
      {stage0_19[160]},
      {stage1_19[69]}
   );
   gpc1_1 gpc1093 (
      {stage0_19[161]},
      {stage1_19[70]}
   );
   gpc1_1 gpc1094 (
      {stage0_20[159]},
      {stage1_20[65]}
   );
   gpc1_1 gpc1095 (
      {stage0_20[160]},
      {stage1_20[66]}
   );
   gpc1_1 gpc1096 (
      {stage0_20[161]},
      {stage1_20[67]}
   );
   gpc1_1 gpc1097 (
      {stage0_21[147]},
      {stage1_21[56]}
   );
   gpc1_1 gpc1098 (
      {stage0_21[148]},
      {stage1_21[57]}
   );
   gpc1_1 gpc1099 (
      {stage0_21[149]},
      {stage1_21[58]}
   );
   gpc1_1 gpc1100 (
      {stage0_21[150]},
      {stage1_21[59]}
   );
   gpc1_1 gpc1101 (
      {stage0_21[151]},
      {stage1_21[60]}
   );
   gpc1_1 gpc1102 (
      {stage0_21[152]},
      {stage1_21[61]}
   );
   gpc1_1 gpc1103 (
      {stage0_21[153]},
      {stage1_21[62]}
   );
   gpc1_1 gpc1104 (
      {stage0_21[154]},
      {stage1_21[63]}
   );
   gpc1_1 gpc1105 (
      {stage0_21[155]},
      {stage1_21[64]}
   );
   gpc1_1 gpc1106 (
      {stage0_21[156]},
      {stage1_21[65]}
   );
   gpc1_1 gpc1107 (
      {stage0_21[157]},
      {stage1_21[66]}
   );
   gpc1_1 gpc1108 (
      {stage0_21[158]},
      {stage1_21[67]}
   );
   gpc1_1 gpc1109 (
      {stage0_21[159]},
      {stage1_21[68]}
   );
   gpc1_1 gpc1110 (
      {stage0_21[160]},
      {stage1_21[69]}
   );
   gpc1_1 gpc1111 (
      {stage0_21[161]},
      {stage1_21[70]}
   );
   gpc1_1 gpc1112 (
      {stage0_23[77]},
      {stage1_23[58]}
   );
   gpc1_1 gpc1113 (
      {stage0_23[78]},
      {stage1_23[59]}
   );
   gpc1_1 gpc1114 (
      {stage0_23[79]},
      {stage1_23[60]}
   );
   gpc1_1 gpc1115 (
      {stage0_23[80]},
      {stage1_23[61]}
   );
   gpc1_1 gpc1116 (
      {stage0_23[81]},
      {stage1_23[62]}
   );
   gpc1_1 gpc1117 (
      {stage0_23[82]},
      {stage1_23[63]}
   );
   gpc1_1 gpc1118 (
      {stage0_23[83]},
      {stage1_23[64]}
   );
   gpc1_1 gpc1119 (
      {stage0_23[84]},
      {stage1_23[65]}
   );
   gpc1_1 gpc1120 (
      {stage0_23[85]},
      {stage1_23[66]}
   );
   gpc1_1 gpc1121 (
      {stage0_23[86]},
      {stage1_23[67]}
   );
   gpc1_1 gpc1122 (
      {stage0_23[87]},
      {stage1_23[68]}
   );
   gpc1_1 gpc1123 (
      {stage0_23[88]},
      {stage1_23[69]}
   );
   gpc1_1 gpc1124 (
      {stage0_23[89]},
      {stage1_23[70]}
   );
   gpc1_1 gpc1125 (
      {stage0_23[90]},
      {stage1_23[71]}
   );
   gpc1_1 gpc1126 (
      {stage0_23[91]},
      {stage1_23[72]}
   );
   gpc1_1 gpc1127 (
      {stage0_23[92]},
      {stage1_23[73]}
   );
   gpc1_1 gpc1128 (
      {stage0_23[93]},
      {stage1_23[74]}
   );
   gpc1_1 gpc1129 (
      {stage0_23[94]},
      {stage1_23[75]}
   );
   gpc1_1 gpc1130 (
      {stage0_23[95]},
      {stage1_23[76]}
   );
   gpc1_1 gpc1131 (
      {stage0_23[96]},
      {stage1_23[77]}
   );
   gpc1_1 gpc1132 (
      {stage0_23[97]},
      {stage1_23[78]}
   );
   gpc1_1 gpc1133 (
      {stage0_23[98]},
      {stage1_23[79]}
   );
   gpc1_1 gpc1134 (
      {stage0_23[99]},
      {stage1_23[80]}
   );
   gpc1_1 gpc1135 (
      {stage0_23[100]},
      {stage1_23[81]}
   );
   gpc1_1 gpc1136 (
      {stage0_23[101]},
      {stage1_23[82]}
   );
   gpc1_1 gpc1137 (
      {stage0_23[102]},
      {stage1_23[83]}
   );
   gpc1_1 gpc1138 (
      {stage0_23[103]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1139 (
      {stage0_23[104]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1140 (
      {stage0_23[105]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1141 (
      {stage0_23[106]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1142 (
      {stage0_23[107]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1143 (
      {stage0_23[108]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1144 (
      {stage0_23[109]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1145 (
      {stage0_23[110]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1146 (
      {stage0_23[111]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1147 (
      {stage0_23[112]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1148 (
      {stage0_23[113]},
      {stage1_23[94]}
   );
   gpc1_1 gpc1149 (
      {stage0_23[114]},
      {stage1_23[95]}
   );
   gpc1_1 gpc1150 (
      {stage0_23[115]},
      {stage1_23[96]}
   );
   gpc1_1 gpc1151 (
      {stage0_23[116]},
      {stage1_23[97]}
   );
   gpc1_1 gpc1152 (
      {stage0_23[117]},
      {stage1_23[98]}
   );
   gpc1_1 gpc1153 (
      {stage0_23[118]},
      {stage1_23[99]}
   );
   gpc1_1 gpc1154 (
      {stage0_23[119]},
      {stage1_23[100]}
   );
   gpc1_1 gpc1155 (
      {stage0_23[120]},
      {stage1_23[101]}
   );
   gpc1_1 gpc1156 (
      {stage0_23[121]},
      {stage1_23[102]}
   );
   gpc1_1 gpc1157 (
      {stage0_23[122]},
      {stage1_23[103]}
   );
   gpc1_1 gpc1158 (
      {stage0_23[123]},
      {stage1_23[104]}
   );
   gpc1_1 gpc1159 (
      {stage0_23[124]},
      {stage1_23[105]}
   );
   gpc1_1 gpc1160 (
      {stage0_23[125]},
      {stage1_23[106]}
   );
   gpc1_1 gpc1161 (
      {stage0_23[126]},
      {stage1_23[107]}
   );
   gpc1_1 gpc1162 (
      {stage0_23[127]},
      {stage1_23[108]}
   );
   gpc1_1 gpc1163 (
      {stage0_23[128]},
      {stage1_23[109]}
   );
   gpc1_1 gpc1164 (
      {stage0_23[129]},
      {stage1_23[110]}
   );
   gpc1_1 gpc1165 (
      {stage0_23[130]},
      {stage1_23[111]}
   );
   gpc1_1 gpc1166 (
      {stage0_23[131]},
      {stage1_23[112]}
   );
   gpc1_1 gpc1167 (
      {stage0_23[132]},
      {stage1_23[113]}
   );
   gpc1_1 gpc1168 (
      {stage0_23[133]},
      {stage1_23[114]}
   );
   gpc1_1 gpc1169 (
      {stage0_23[134]},
      {stage1_23[115]}
   );
   gpc1_1 gpc1170 (
      {stage0_23[135]},
      {stage1_23[116]}
   );
   gpc1_1 gpc1171 (
      {stage0_23[136]},
      {stage1_23[117]}
   );
   gpc1_1 gpc1172 (
      {stage0_23[137]},
      {stage1_23[118]}
   );
   gpc1_1 gpc1173 (
      {stage0_23[138]},
      {stage1_23[119]}
   );
   gpc1_1 gpc1174 (
      {stage0_23[139]},
      {stage1_23[120]}
   );
   gpc1_1 gpc1175 (
      {stage0_23[140]},
      {stage1_23[121]}
   );
   gpc1_1 gpc1176 (
      {stage0_23[141]},
      {stage1_23[122]}
   );
   gpc1_1 gpc1177 (
      {stage0_23[142]},
      {stage1_23[123]}
   );
   gpc1_1 gpc1178 (
      {stage0_23[143]},
      {stage1_23[124]}
   );
   gpc1_1 gpc1179 (
      {stage0_23[144]},
      {stage1_23[125]}
   );
   gpc1_1 gpc1180 (
      {stage0_23[145]},
      {stage1_23[126]}
   );
   gpc1_1 gpc1181 (
      {stage0_23[146]},
      {stage1_23[127]}
   );
   gpc1_1 gpc1182 (
      {stage0_23[147]},
      {stage1_23[128]}
   );
   gpc1_1 gpc1183 (
      {stage0_23[148]},
      {stage1_23[129]}
   );
   gpc1_1 gpc1184 (
      {stage0_23[149]},
      {stage1_23[130]}
   );
   gpc1_1 gpc1185 (
      {stage0_23[150]},
      {stage1_23[131]}
   );
   gpc1_1 gpc1186 (
      {stage0_23[151]},
      {stage1_23[132]}
   );
   gpc1_1 gpc1187 (
      {stage0_23[152]},
      {stage1_23[133]}
   );
   gpc1_1 gpc1188 (
      {stage0_23[153]},
      {stage1_23[134]}
   );
   gpc1_1 gpc1189 (
      {stage0_23[154]},
      {stage1_23[135]}
   );
   gpc1_1 gpc1190 (
      {stage0_23[155]},
      {stage1_23[136]}
   );
   gpc1_1 gpc1191 (
      {stage0_23[156]},
      {stage1_23[137]}
   );
   gpc1_1 gpc1192 (
      {stage0_23[157]},
      {stage1_23[138]}
   );
   gpc1_1 gpc1193 (
      {stage0_23[158]},
      {stage1_23[139]}
   );
   gpc1_1 gpc1194 (
      {stage0_23[159]},
      {stage1_23[140]}
   );
   gpc1_1 gpc1195 (
      {stage0_23[160]},
      {stage1_23[141]}
   );
   gpc1_1 gpc1196 (
      {stage0_23[161]},
      {stage1_23[142]}
   );
   gpc1_1 gpc1197 (
      {stage0_24[126]},
      {stage1_24[47]}
   );
   gpc1_1 gpc1198 (
      {stage0_24[127]},
      {stage1_24[48]}
   );
   gpc1_1 gpc1199 (
      {stage0_24[128]},
      {stage1_24[49]}
   );
   gpc1_1 gpc1200 (
      {stage0_24[129]},
      {stage1_24[50]}
   );
   gpc1_1 gpc1201 (
      {stage0_24[130]},
      {stage1_24[51]}
   );
   gpc1_1 gpc1202 (
      {stage0_24[131]},
      {stage1_24[52]}
   );
   gpc1_1 gpc1203 (
      {stage0_24[132]},
      {stage1_24[53]}
   );
   gpc1_1 gpc1204 (
      {stage0_24[133]},
      {stage1_24[54]}
   );
   gpc1_1 gpc1205 (
      {stage0_24[134]},
      {stage1_24[55]}
   );
   gpc1_1 gpc1206 (
      {stage0_24[135]},
      {stage1_24[56]}
   );
   gpc1_1 gpc1207 (
      {stage0_24[136]},
      {stage1_24[57]}
   );
   gpc1_1 gpc1208 (
      {stage0_24[137]},
      {stage1_24[58]}
   );
   gpc1_1 gpc1209 (
      {stage0_24[138]},
      {stage1_24[59]}
   );
   gpc1_1 gpc1210 (
      {stage0_24[139]},
      {stage1_24[60]}
   );
   gpc1_1 gpc1211 (
      {stage0_24[140]},
      {stage1_24[61]}
   );
   gpc1_1 gpc1212 (
      {stage0_24[141]},
      {stage1_24[62]}
   );
   gpc1_1 gpc1213 (
      {stage0_24[142]},
      {stage1_24[63]}
   );
   gpc1_1 gpc1214 (
      {stage0_24[143]},
      {stage1_24[64]}
   );
   gpc1_1 gpc1215 (
      {stage0_24[144]},
      {stage1_24[65]}
   );
   gpc1_1 gpc1216 (
      {stage0_24[145]},
      {stage1_24[66]}
   );
   gpc1_1 gpc1217 (
      {stage0_24[146]},
      {stage1_24[67]}
   );
   gpc1_1 gpc1218 (
      {stage0_24[147]},
      {stage1_24[68]}
   );
   gpc1_1 gpc1219 (
      {stage0_24[148]},
      {stage1_24[69]}
   );
   gpc1_1 gpc1220 (
      {stage0_24[149]},
      {stage1_24[70]}
   );
   gpc1_1 gpc1221 (
      {stage0_24[150]},
      {stage1_24[71]}
   );
   gpc1_1 gpc1222 (
      {stage0_24[151]},
      {stage1_24[72]}
   );
   gpc1_1 gpc1223 (
      {stage0_24[152]},
      {stage1_24[73]}
   );
   gpc1_1 gpc1224 (
      {stage0_24[153]},
      {stage1_24[74]}
   );
   gpc1_1 gpc1225 (
      {stage0_24[154]},
      {stage1_24[75]}
   );
   gpc1_1 gpc1226 (
      {stage0_24[155]},
      {stage1_24[76]}
   );
   gpc1_1 gpc1227 (
      {stage0_24[156]},
      {stage1_24[77]}
   );
   gpc1_1 gpc1228 (
      {stage0_24[157]},
      {stage1_24[78]}
   );
   gpc1_1 gpc1229 (
      {stage0_24[158]},
      {stage1_24[79]}
   );
   gpc1_1 gpc1230 (
      {stage0_24[159]},
      {stage1_24[80]}
   );
   gpc1_1 gpc1231 (
      {stage0_24[160]},
      {stage1_24[81]}
   );
   gpc1_1 gpc1232 (
      {stage0_24[161]},
      {stage1_24[82]}
   );
   gpc1_1 gpc1233 (
      {stage0_25[127]},
      {stage1_25[50]}
   );
   gpc1_1 gpc1234 (
      {stage0_25[128]},
      {stage1_25[51]}
   );
   gpc1_1 gpc1235 (
      {stage0_25[129]},
      {stage1_25[52]}
   );
   gpc1_1 gpc1236 (
      {stage0_25[130]},
      {stage1_25[53]}
   );
   gpc1_1 gpc1237 (
      {stage0_25[131]},
      {stage1_25[54]}
   );
   gpc1_1 gpc1238 (
      {stage0_25[132]},
      {stage1_25[55]}
   );
   gpc1_1 gpc1239 (
      {stage0_25[133]},
      {stage1_25[56]}
   );
   gpc1_1 gpc1240 (
      {stage0_25[134]},
      {stage1_25[57]}
   );
   gpc1_1 gpc1241 (
      {stage0_25[135]},
      {stage1_25[58]}
   );
   gpc1_1 gpc1242 (
      {stage0_25[136]},
      {stage1_25[59]}
   );
   gpc1_1 gpc1243 (
      {stage0_25[137]},
      {stage1_25[60]}
   );
   gpc1_1 gpc1244 (
      {stage0_25[138]},
      {stage1_25[61]}
   );
   gpc1_1 gpc1245 (
      {stage0_25[139]},
      {stage1_25[62]}
   );
   gpc1_1 gpc1246 (
      {stage0_25[140]},
      {stage1_25[63]}
   );
   gpc1_1 gpc1247 (
      {stage0_25[141]},
      {stage1_25[64]}
   );
   gpc1_1 gpc1248 (
      {stage0_25[142]},
      {stage1_25[65]}
   );
   gpc1_1 gpc1249 (
      {stage0_25[143]},
      {stage1_25[66]}
   );
   gpc1_1 gpc1250 (
      {stage0_25[144]},
      {stage1_25[67]}
   );
   gpc1_1 gpc1251 (
      {stage0_25[145]},
      {stage1_25[68]}
   );
   gpc1_1 gpc1252 (
      {stage0_25[146]},
      {stage1_25[69]}
   );
   gpc1_1 gpc1253 (
      {stage0_25[147]},
      {stage1_25[70]}
   );
   gpc1_1 gpc1254 (
      {stage0_25[148]},
      {stage1_25[71]}
   );
   gpc1_1 gpc1255 (
      {stage0_25[149]},
      {stage1_25[72]}
   );
   gpc1_1 gpc1256 (
      {stage0_25[150]},
      {stage1_25[73]}
   );
   gpc1_1 gpc1257 (
      {stage0_25[151]},
      {stage1_25[74]}
   );
   gpc1_1 gpc1258 (
      {stage0_25[152]},
      {stage1_25[75]}
   );
   gpc1_1 gpc1259 (
      {stage0_25[153]},
      {stage1_25[76]}
   );
   gpc1_1 gpc1260 (
      {stage0_25[154]},
      {stage1_25[77]}
   );
   gpc1_1 gpc1261 (
      {stage0_25[155]},
      {stage1_25[78]}
   );
   gpc1_1 gpc1262 (
      {stage0_25[156]},
      {stage1_25[79]}
   );
   gpc1_1 gpc1263 (
      {stage0_25[157]},
      {stage1_25[80]}
   );
   gpc1_1 gpc1264 (
      {stage0_25[158]},
      {stage1_25[81]}
   );
   gpc1_1 gpc1265 (
      {stage0_25[159]},
      {stage1_25[82]}
   );
   gpc1_1 gpc1266 (
      {stage0_25[160]},
      {stage1_25[83]}
   );
   gpc1_1 gpc1267 (
      {stage0_25[161]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[149]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[150]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[151]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[152]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[153]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[154]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[155]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[156]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[157]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[158]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[159]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[160]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[161]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1281 (
      {stage0_27[142]},
      {stage1_27[54]}
   );
   gpc1_1 gpc1282 (
      {stage0_27[143]},
      {stage1_27[55]}
   );
   gpc1_1 gpc1283 (
      {stage0_27[144]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1284 (
      {stage0_27[145]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1285 (
      {stage0_27[146]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1286 (
      {stage0_27[147]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1287 (
      {stage0_27[148]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1288 (
      {stage0_27[149]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1289 (
      {stage0_27[150]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1290 (
      {stage0_27[151]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1291 (
      {stage0_27[152]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1292 (
      {stage0_27[153]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1293 (
      {stage0_27[154]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1294 (
      {stage0_27[155]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1295 (
      {stage0_27[156]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1296 (
      {stage0_27[157]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1297 (
      {stage0_27[158]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1298 (
      {stage0_27[159]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1299 (
      {stage0_27[160]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1300 (
      {stage0_27[161]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1301 (
      {stage0_28[140]},
      {stage1_28[55]}
   );
   gpc1_1 gpc1302 (
      {stage0_28[141]},
      {stage1_28[56]}
   );
   gpc1_1 gpc1303 (
      {stage0_28[142]},
      {stage1_28[57]}
   );
   gpc1_1 gpc1304 (
      {stage0_28[143]},
      {stage1_28[58]}
   );
   gpc1_1 gpc1305 (
      {stage0_28[144]},
      {stage1_28[59]}
   );
   gpc1_1 gpc1306 (
      {stage0_28[145]},
      {stage1_28[60]}
   );
   gpc1_1 gpc1307 (
      {stage0_28[146]},
      {stage1_28[61]}
   );
   gpc1_1 gpc1308 (
      {stage0_28[147]},
      {stage1_28[62]}
   );
   gpc1_1 gpc1309 (
      {stage0_28[148]},
      {stage1_28[63]}
   );
   gpc1_1 gpc1310 (
      {stage0_28[149]},
      {stage1_28[64]}
   );
   gpc1_1 gpc1311 (
      {stage0_28[150]},
      {stage1_28[65]}
   );
   gpc1_1 gpc1312 (
      {stage0_28[151]},
      {stage1_28[66]}
   );
   gpc1_1 gpc1313 (
      {stage0_28[152]},
      {stage1_28[67]}
   );
   gpc1_1 gpc1314 (
      {stage0_28[153]},
      {stage1_28[68]}
   );
   gpc1_1 gpc1315 (
      {stage0_28[154]},
      {stage1_28[69]}
   );
   gpc1_1 gpc1316 (
      {stage0_28[155]},
      {stage1_28[70]}
   );
   gpc1_1 gpc1317 (
      {stage0_28[156]},
      {stage1_28[71]}
   );
   gpc1_1 gpc1318 (
      {stage0_28[157]},
      {stage1_28[72]}
   );
   gpc1_1 gpc1319 (
      {stage0_28[158]},
      {stage1_28[73]}
   );
   gpc1_1 gpc1320 (
      {stage0_28[159]},
      {stage1_28[74]}
   );
   gpc1_1 gpc1321 (
      {stage0_28[160]},
      {stage1_28[75]}
   );
   gpc1_1 gpc1322 (
      {stage0_28[161]},
      {stage1_28[76]}
   );
   gpc1_1 gpc1323 (
      {stage0_29[144]},
      {stage1_29[63]}
   );
   gpc1_1 gpc1324 (
      {stage0_29[145]},
      {stage1_29[64]}
   );
   gpc1_1 gpc1325 (
      {stage0_29[146]},
      {stage1_29[65]}
   );
   gpc1_1 gpc1326 (
      {stage0_29[147]},
      {stage1_29[66]}
   );
   gpc1_1 gpc1327 (
      {stage0_29[148]},
      {stage1_29[67]}
   );
   gpc1_1 gpc1328 (
      {stage0_29[149]},
      {stage1_29[68]}
   );
   gpc1_1 gpc1329 (
      {stage0_29[150]},
      {stage1_29[69]}
   );
   gpc1_1 gpc1330 (
      {stage0_29[151]},
      {stage1_29[70]}
   );
   gpc1_1 gpc1331 (
      {stage0_29[152]},
      {stage1_29[71]}
   );
   gpc1_1 gpc1332 (
      {stage0_29[153]},
      {stage1_29[72]}
   );
   gpc1_1 gpc1333 (
      {stage0_29[154]},
      {stage1_29[73]}
   );
   gpc1_1 gpc1334 (
      {stage0_29[155]},
      {stage1_29[74]}
   );
   gpc1_1 gpc1335 (
      {stage0_29[156]},
      {stage1_29[75]}
   );
   gpc1_1 gpc1336 (
      {stage0_29[157]},
      {stage1_29[76]}
   );
   gpc1_1 gpc1337 (
      {stage0_29[158]},
      {stage1_29[77]}
   );
   gpc1_1 gpc1338 (
      {stage0_29[159]},
      {stage1_29[78]}
   );
   gpc1_1 gpc1339 (
      {stage0_29[160]},
      {stage1_29[79]}
   );
   gpc1_1 gpc1340 (
      {stage0_29[161]},
      {stage1_29[80]}
   );
   gpc1_1 gpc1341 (
      {stage0_30[111]},
      {stage1_30[56]}
   );
   gpc1_1 gpc1342 (
      {stage0_30[112]},
      {stage1_30[57]}
   );
   gpc1_1 gpc1343 (
      {stage0_30[113]},
      {stage1_30[58]}
   );
   gpc1_1 gpc1344 (
      {stage0_30[114]},
      {stage1_30[59]}
   );
   gpc1_1 gpc1345 (
      {stage0_30[115]},
      {stage1_30[60]}
   );
   gpc1_1 gpc1346 (
      {stage0_30[116]},
      {stage1_30[61]}
   );
   gpc1_1 gpc1347 (
      {stage0_30[117]},
      {stage1_30[62]}
   );
   gpc1_1 gpc1348 (
      {stage0_30[118]},
      {stage1_30[63]}
   );
   gpc1_1 gpc1349 (
      {stage0_30[119]},
      {stage1_30[64]}
   );
   gpc1_1 gpc1350 (
      {stage0_30[120]},
      {stage1_30[65]}
   );
   gpc1_1 gpc1351 (
      {stage0_30[121]},
      {stage1_30[66]}
   );
   gpc1_1 gpc1352 (
      {stage0_30[122]},
      {stage1_30[67]}
   );
   gpc1_1 gpc1353 (
      {stage0_30[123]},
      {stage1_30[68]}
   );
   gpc1_1 gpc1354 (
      {stage0_30[124]},
      {stage1_30[69]}
   );
   gpc1_1 gpc1355 (
      {stage0_30[125]},
      {stage1_30[70]}
   );
   gpc1_1 gpc1356 (
      {stage0_30[126]},
      {stage1_30[71]}
   );
   gpc1_1 gpc1357 (
      {stage0_30[127]},
      {stage1_30[72]}
   );
   gpc1_1 gpc1358 (
      {stage0_30[128]},
      {stage1_30[73]}
   );
   gpc1_1 gpc1359 (
      {stage0_30[129]},
      {stage1_30[74]}
   );
   gpc1_1 gpc1360 (
      {stage0_30[130]},
      {stage1_30[75]}
   );
   gpc1_1 gpc1361 (
      {stage0_30[131]},
      {stage1_30[76]}
   );
   gpc1_1 gpc1362 (
      {stage0_30[132]},
      {stage1_30[77]}
   );
   gpc1_1 gpc1363 (
      {stage0_30[133]},
      {stage1_30[78]}
   );
   gpc1_1 gpc1364 (
      {stage0_30[134]},
      {stage1_30[79]}
   );
   gpc1_1 gpc1365 (
      {stage0_30[135]},
      {stage1_30[80]}
   );
   gpc1_1 gpc1366 (
      {stage0_30[136]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1367 (
      {stage0_30[137]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1368 (
      {stage0_30[138]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1369 (
      {stage0_30[139]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1370 (
      {stage0_30[140]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1371 (
      {stage0_30[141]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1372 (
      {stage0_30[142]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1373 (
      {stage0_30[143]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1374 (
      {stage0_30[144]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1375 (
      {stage0_30[145]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1376 (
      {stage0_30[146]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1377 (
      {stage0_30[147]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1378 (
      {stage0_30[148]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1379 (
      {stage0_30[149]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1380 (
      {stage0_30[150]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1381 (
      {stage0_30[151]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1382 (
      {stage0_30[152]},
      {stage1_30[97]}
   );
   gpc1_1 gpc1383 (
      {stage0_30[153]},
      {stage1_30[98]}
   );
   gpc1_1 gpc1384 (
      {stage0_30[154]},
      {stage1_30[99]}
   );
   gpc1_1 gpc1385 (
      {stage0_30[155]},
      {stage1_30[100]}
   );
   gpc1_1 gpc1386 (
      {stage0_30[156]},
      {stage1_30[101]}
   );
   gpc1_1 gpc1387 (
      {stage0_30[157]},
      {stage1_30[102]}
   );
   gpc1_1 gpc1388 (
      {stage0_30[158]},
      {stage1_30[103]}
   );
   gpc1_1 gpc1389 (
      {stage0_30[159]},
      {stage1_30[104]}
   );
   gpc1_1 gpc1390 (
      {stage0_30[160]},
      {stage1_30[105]}
   );
   gpc1_1 gpc1391 (
      {stage0_30[161]},
      {stage1_30[106]}
   );
   gpc1_1 gpc1392 (
      {stage0_31[109]},
      {stage1_31[44]}
   );
   gpc1_1 gpc1393 (
      {stage0_31[110]},
      {stage1_31[45]}
   );
   gpc1_1 gpc1394 (
      {stage0_31[111]},
      {stage1_31[46]}
   );
   gpc1_1 gpc1395 (
      {stage0_31[112]},
      {stage1_31[47]}
   );
   gpc1_1 gpc1396 (
      {stage0_31[113]},
      {stage1_31[48]}
   );
   gpc1_1 gpc1397 (
      {stage0_31[114]},
      {stage1_31[49]}
   );
   gpc1_1 gpc1398 (
      {stage0_31[115]},
      {stage1_31[50]}
   );
   gpc1_1 gpc1399 (
      {stage0_31[116]},
      {stage1_31[51]}
   );
   gpc1_1 gpc1400 (
      {stage0_31[117]},
      {stage1_31[52]}
   );
   gpc1_1 gpc1401 (
      {stage0_31[118]},
      {stage1_31[53]}
   );
   gpc1_1 gpc1402 (
      {stage0_31[119]},
      {stage1_31[54]}
   );
   gpc1_1 gpc1403 (
      {stage0_31[120]},
      {stage1_31[55]}
   );
   gpc1_1 gpc1404 (
      {stage0_31[121]},
      {stage1_31[56]}
   );
   gpc1_1 gpc1405 (
      {stage0_31[122]},
      {stage1_31[57]}
   );
   gpc1_1 gpc1406 (
      {stage0_31[123]},
      {stage1_31[58]}
   );
   gpc1_1 gpc1407 (
      {stage0_31[124]},
      {stage1_31[59]}
   );
   gpc1_1 gpc1408 (
      {stage0_31[125]},
      {stage1_31[60]}
   );
   gpc1_1 gpc1409 (
      {stage0_31[126]},
      {stage1_31[61]}
   );
   gpc1_1 gpc1410 (
      {stage0_31[127]},
      {stage1_31[62]}
   );
   gpc1_1 gpc1411 (
      {stage0_31[128]},
      {stage1_31[63]}
   );
   gpc1_1 gpc1412 (
      {stage0_31[129]},
      {stage1_31[64]}
   );
   gpc1_1 gpc1413 (
      {stage0_31[130]},
      {stage1_31[65]}
   );
   gpc1_1 gpc1414 (
      {stage0_31[131]},
      {stage1_31[66]}
   );
   gpc1_1 gpc1415 (
      {stage0_31[132]},
      {stage1_31[67]}
   );
   gpc1_1 gpc1416 (
      {stage0_31[133]},
      {stage1_31[68]}
   );
   gpc1_1 gpc1417 (
      {stage0_31[134]},
      {stage1_31[69]}
   );
   gpc1_1 gpc1418 (
      {stage0_31[135]},
      {stage1_31[70]}
   );
   gpc1_1 gpc1419 (
      {stage0_31[136]},
      {stage1_31[71]}
   );
   gpc1_1 gpc1420 (
      {stage0_31[137]},
      {stage1_31[72]}
   );
   gpc1_1 gpc1421 (
      {stage0_31[138]},
      {stage1_31[73]}
   );
   gpc1_1 gpc1422 (
      {stage0_31[139]},
      {stage1_31[74]}
   );
   gpc1_1 gpc1423 (
      {stage0_31[140]},
      {stage1_31[75]}
   );
   gpc1_1 gpc1424 (
      {stage0_31[141]},
      {stage1_31[76]}
   );
   gpc1_1 gpc1425 (
      {stage0_31[142]},
      {stage1_31[77]}
   );
   gpc1_1 gpc1426 (
      {stage0_31[143]},
      {stage1_31[78]}
   );
   gpc1_1 gpc1427 (
      {stage0_31[144]},
      {stage1_31[79]}
   );
   gpc1_1 gpc1428 (
      {stage0_31[145]},
      {stage1_31[80]}
   );
   gpc1_1 gpc1429 (
      {stage0_31[146]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1430 (
      {stage0_31[147]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1431 (
      {stage0_31[148]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1432 (
      {stage0_31[149]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1433 (
      {stage0_31[150]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1434 (
      {stage0_31[151]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1435 (
      {stage0_31[152]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1436 (
      {stage0_31[153]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1437 (
      {stage0_31[154]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1438 (
      {stage0_31[155]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1439 (
      {stage0_31[156]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1440 (
      {stage0_31[157]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1441 (
      {stage0_31[158]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1442 (
      {stage0_31[159]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1443 (
      {stage0_31[160]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1444 (
      {stage0_31[161]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1445 (
      {stage0_32[129]},
      {stage1_32[54]}
   );
   gpc1_1 gpc1446 (
      {stage0_32[130]},
      {stage1_32[55]}
   );
   gpc1_1 gpc1447 (
      {stage0_32[131]},
      {stage1_32[56]}
   );
   gpc1_1 gpc1448 (
      {stage0_32[132]},
      {stage1_32[57]}
   );
   gpc1_1 gpc1449 (
      {stage0_32[133]},
      {stage1_32[58]}
   );
   gpc1_1 gpc1450 (
      {stage0_32[134]},
      {stage1_32[59]}
   );
   gpc1_1 gpc1451 (
      {stage0_32[135]},
      {stage1_32[60]}
   );
   gpc1_1 gpc1452 (
      {stage0_32[136]},
      {stage1_32[61]}
   );
   gpc1_1 gpc1453 (
      {stage0_32[137]},
      {stage1_32[62]}
   );
   gpc1_1 gpc1454 (
      {stage0_32[138]},
      {stage1_32[63]}
   );
   gpc1_1 gpc1455 (
      {stage0_32[139]},
      {stage1_32[64]}
   );
   gpc1_1 gpc1456 (
      {stage0_32[140]},
      {stage1_32[65]}
   );
   gpc1_1 gpc1457 (
      {stage0_32[141]},
      {stage1_32[66]}
   );
   gpc1_1 gpc1458 (
      {stage0_32[142]},
      {stage1_32[67]}
   );
   gpc1_1 gpc1459 (
      {stage0_32[143]},
      {stage1_32[68]}
   );
   gpc1_1 gpc1460 (
      {stage0_32[144]},
      {stage1_32[69]}
   );
   gpc1_1 gpc1461 (
      {stage0_32[145]},
      {stage1_32[70]}
   );
   gpc1_1 gpc1462 (
      {stage0_32[146]},
      {stage1_32[71]}
   );
   gpc1_1 gpc1463 (
      {stage0_32[147]},
      {stage1_32[72]}
   );
   gpc1_1 gpc1464 (
      {stage0_32[148]},
      {stage1_32[73]}
   );
   gpc1_1 gpc1465 (
      {stage0_32[149]},
      {stage1_32[74]}
   );
   gpc1_1 gpc1466 (
      {stage0_32[150]},
      {stage1_32[75]}
   );
   gpc1_1 gpc1467 (
      {stage0_32[151]},
      {stage1_32[76]}
   );
   gpc1_1 gpc1468 (
      {stage0_32[152]},
      {stage1_32[77]}
   );
   gpc1_1 gpc1469 (
      {stage0_32[153]},
      {stage1_32[78]}
   );
   gpc1_1 gpc1470 (
      {stage0_32[154]},
      {stage1_32[79]}
   );
   gpc1_1 gpc1471 (
      {stage0_32[155]},
      {stage1_32[80]}
   );
   gpc1_1 gpc1472 (
      {stage0_32[156]},
      {stage1_32[81]}
   );
   gpc1_1 gpc1473 (
      {stage0_32[157]},
      {stage1_32[82]}
   );
   gpc1_1 gpc1474 (
      {stage0_32[158]},
      {stage1_32[83]}
   );
   gpc1_1 gpc1475 (
      {stage0_32[159]},
      {stage1_32[84]}
   );
   gpc1_1 gpc1476 (
      {stage0_32[160]},
      {stage1_32[85]}
   );
   gpc1_1 gpc1477 (
      {stage0_32[161]},
      {stage1_32[86]}
   );
   gpc1_1 gpc1478 (
      {stage0_33[136]},
      {stage1_33[64]}
   );
   gpc1_1 gpc1479 (
      {stage0_33[137]},
      {stage1_33[65]}
   );
   gpc1_1 gpc1480 (
      {stage0_33[138]},
      {stage1_33[66]}
   );
   gpc1_1 gpc1481 (
      {stage0_33[139]},
      {stage1_33[67]}
   );
   gpc1_1 gpc1482 (
      {stage0_33[140]},
      {stage1_33[68]}
   );
   gpc1_1 gpc1483 (
      {stage0_33[141]},
      {stage1_33[69]}
   );
   gpc1_1 gpc1484 (
      {stage0_33[142]},
      {stage1_33[70]}
   );
   gpc1_1 gpc1485 (
      {stage0_33[143]},
      {stage1_33[71]}
   );
   gpc1_1 gpc1486 (
      {stage0_33[144]},
      {stage1_33[72]}
   );
   gpc1_1 gpc1487 (
      {stage0_33[145]},
      {stage1_33[73]}
   );
   gpc1_1 gpc1488 (
      {stage0_33[146]},
      {stage1_33[74]}
   );
   gpc1_1 gpc1489 (
      {stage0_33[147]},
      {stage1_33[75]}
   );
   gpc1_1 gpc1490 (
      {stage0_33[148]},
      {stage1_33[76]}
   );
   gpc1_1 gpc1491 (
      {stage0_33[149]},
      {stage1_33[77]}
   );
   gpc1_1 gpc1492 (
      {stage0_33[150]},
      {stage1_33[78]}
   );
   gpc1_1 gpc1493 (
      {stage0_33[151]},
      {stage1_33[79]}
   );
   gpc1_1 gpc1494 (
      {stage0_33[152]},
      {stage1_33[80]}
   );
   gpc1_1 gpc1495 (
      {stage0_33[153]},
      {stage1_33[81]}
   );
   gpc1_1 gpc1496 (
      {stage0_33[154]},
      {stage1_33[82]}
   );
   gpc1_1 gpc1497 (
      {stage0_33[155]},
      {stage1_33[83]}
   );
   gpc1_1 gpc1498 (
      {stage0_33[156]},
      {stage1_33[84]}
   );
   gpc1_1 gpc1499 (
      {stage0_33[157]},
      {stage1_33[85]}
   );
   gpc1_1 gpc1500 (
      {stage0_33[158]},
      {stage1_33[86]}
   );
   gpc1_1 gpc1501 (
      {stage0_33[159]},
      {stage1_33[87]}
   );
   gpc1_1 gpc1502 (
      {stage0_33[160]},
      {stage1_33[88]}
   );
   gpc1_1 gpc1503 (
      {stage0_33[161]},
      {stage1_33[89]}
   );
   gpc1_1 gpc1504 (
      {stage0_34[158]},
      {stage1_34[52]}
   );
   gpc1_1 gpc1505 (
      {stage0_34[159]},
      {stage1_34[53]}
   );
   gpc1_1 gpc1506 (
      {stage0_34[160]},
      {stage1_34[54]}
   );
   gpc1_1 gpc1507 (
      {stage0_34[161]},
      {stage1_34[55]}
   );
   gpc1_1 gpc1508 (
      {stage0_35[158]},
      {stage1_35[56]}
   );
   gpc1_1 gpc1509 (
      {stage0_35[159]},
      {stage1_35[57]}
   );
   gpc1_1 gpc1510 (
      {stage0_35[160]},
      {stage1_35[58]}
   );
   gpc1_1 gpc1511 (
      {stage0_35[161]},
      {stage1_35[59]}
   );
   gpc1_1 gpc1512 (
      {stage0_36[146]},
      {stage1_36[67]}
   );
   gpc1_1 gpc1513 (
      {stage0_36[147]},
      {stage1_36[68]}
   );
   gpc1_1 gpc1514 (
      {stage0_36[148]},
      {stage1_36[69]}
   );
   gpc1_1 gpc1515 (
      {stage0_36[149]},
      {stage1_36[70]}
   );
   gpc1_1 gpc1516 (
      {stage0_36[150]},
      {stage1_36[71]}
   );
   gpc1_1 gpc1517 (
      {stage0_36[151]},
      {stage1_36[72]}
   );
   gpc1_1 gpc1518 (
      {stage0_36[152]},
      {stage1_36[73]}
   );
   gpc1_1 gpc1519 (
      {stage0_36[153]},
      {stage1_36[74]}
   );
   gpc1_1 gpc1520 (
      {stage0_36[154]},
      {stage1_36[75]}
   );
   gpc1_1 gpc1521 (
      {stage0_36[155]},
      {stage1_36[76]}
   );
   gpc1_1 gpc1522 (
      {stage0_36[156]},
      {stage1_36[77]}
   );
   gpc1_1 gpc1523 (
      {stage0_36[157]},
      {stage1_36[78]}
   );
   gpc1_1 gpc1524 (
      {stage0_36[158]},
      {stage1_36[79]}
   );
   gpc1_1 gpc1525 (
      {stage0_36[159]},
      {stage1_36[80]}
   );
   gpc1_1 gpc1526 (
      {stage0_36[160]},
      {stage1_36[81]}
   );
   gpc1_1 gpc1527 (
      {stage0_36[161]},
      {stage1_36[82]}
   );
   gpc1_1 gpc1528 (
      {stage0_37[90]},
      {stage1_37[56]}
   );
   gpc1_1 gpc1529 (
      {stage0_37[91]},
      {stage1_37[57]}
   );
   gpc1_1 gpc1530 (
      {stage0_37[92]},
      {stage1_37[58]}
   );
   gpc1_1 gpc1531 (
      {stage0_37[93]},
      {stage1_37[59]}
   );
   gpc1_1 gpc1532 (
      {stage0_37[94]},
      {stage1_37[60]}
   );
   gpc1_1 gpc1533 (
      {stage0_37[95]},
      {stage1_37[61]}
   );
   gpc1_1 gpc1534 (
      {stage0_37[96]},
      {stage1_37[62]}
   );
   gpc1_1 gpc1535 (
      {stage0_37[97]},
      {stage1_37[63]}
   );
   gpc1_1 gpc1536 (
      {stage0_37[98]},
      {stage1_37[64]}
   );
   gpc1_1 gpc1537 (
      {stage0_37[99]},
      {stage1_37[65]}
   );
   gpc1_1 gpc1538 (
      {stage0_37[100]},
      {stage1_37[66]}
   );
   gpc1_1 gpc1539 (
      {stage0_37[101]},
      {stage1_37[67]}
   );
   gpc1_1 gpc1540 (
      {stage0_37[102]},
      {stage1_37[68]}
   );
   gpc1_1 gpc1541 (
      {stage0_37[103]},
      {stage1_37[69]}
   );
   gpc1_1 gpc1542 (
      {stage0_37[104]},
      {stage1_37[70]}
   );
   gpc1_1 gpc1543 (
      {stage0_37[105]},
      {stage1_37[71]}
   );
   gpc1_1 gpc1544 (
      {stage0_37[106]},
      {stage1_37[72]}
   );
   gpc1_1 gpc1545 (
      {stage0_37[107]},
      {stage1_37[73]}
   );
   gpc1_1 gpc1546 (
      {stage0_37[108]},
      {stage1_37[74]}
   );
   gpc1_1 gpc1547 (
      {stage0_37[109]},
      {stage1_37[75]}
   );
   gpc1_1 gpc1548 (
      {stage0_37[110]},
      {stage1_37[76]}
   );
   gpc1_1 gpc1549 (
      {stage0_37[111]},
      {stage1_37[77]}
   );
   gpc1_1 gpc1550 (
      {stage0_37[112]},
      {stage1_37[78]}
   );
   gpc1_1 gpc1551 (
      {stage0_37[113]},
      {stage1_37[79]}
   );
   gpc1_1 gpc1552 (
      {stage0_37[114]},
      {stage1_37[80]}
   );
   gpc1_1 gpc1553 (
      {stage0_37[115]},
      {stage1_37[81]}
   );
   gpc1_1 gpc1554 (
      {stage0_37[116]},
      {stage1_37[82]}
   );
   gpc1_1 gpc1555 (
      {stage0_37[117]},
      {stage1_37[83]}
   );
   gpc1_1 gpc1556 (
      {stage0_37[118]},
      {stage1_37[84]}
   );
   gpc1_1 gpc1557 (
      {stage0_37[119]},
      {stage1_37[85]}
   );
   gpc1_1 gpc1558 (
      {stage0_37[120]},
      {stage1_37[86]}
   );
   gpc1_1 gpc1559 (
      {stage0_37[121]},
      {stage1_37[87]}
   );
   gpc1_1 gpc1560 (
      {stage0_37[122]},
      {stage1_37[88]}
   );
   gpc1_1 gpc1561 (
      {stage0_37[123]},
      {stage1_37[89]}
   );
   gpc1_1 gpc1562 (
      {stage0_37[124]},
      {stage1_37[90]}
   );
   gpc1_1 gpc1563 (
      {stage0_37[125]},
      {stage1_37[91]}
   );
   gpc1_1 gpc1564 (
      {stage0_37[126]},
      {stage1_37[92]}
   );
   gpc1_1 gpc1565 (
      {stage0_37[127]},
      {stage1_37[93]}
   );
   gpc1_1 gpc1566 (
      {stage0_37[128]},
      {stage1_37[94]}
   );
   gpc1_1 gpc1567 (
      {stage0_37[129]},
      {stage1_37[95]}
   );
   gpc1_1 gpc1568 (
      {stage0_37[130]},
      {stage1_37[96]}
   );
   gpc1_1 gpc1569 (
      {stage0_37[131]},
      {stage1_37[97]}
   );
   gpc1_1 gpc1570 (
      {stage0_37[132]},
      {stage1_37[98]}
   );
   gpc1_1 gpc1571 (
      {stage0_37[133]},
      {stage1_37[99]}
   );
   gpc1_1 gpc1572 (
      {stage0_37[134]},
      {stage1_37[100]}
   );
   gpc1_1 gpc1573 (
      {stage0_37[135]},
      {stage1_37[101]}
   );
   gpc1_1 gpc1574 (
      {stage0_37[136]},
      {stage1_37[102]}
   );
   gpc1_1 gpc1575 (
      {stage0_37[137]},
      {stage1_37[103]}
   );
   gpc1_1 gpc1576 (
      {stage0_37[138]},
      {stage1_37[104]}
   );
   gpc1_1 gpc1577 (
      {stage0_37[139]},
      {stage1_37[105]}
   );
   gpc1_1 gpc1578 (
      {stage0_37[140]},
      {stage1_37[106]}
   );
   gpc1_1 gpc1579 (
      {stage0_37[141]},
      {stage1_37[107]}
   );
   gpc1_1 gpc1580 (
      {stage0_37[142]},
      {stage1_37[108]}
   );
   gpc1_1 gpc1581 (
      {stage0_37[143]},
      {stage1_37[109]}
   );
   gpc1_1 gpc1582 (
      {stage0_37[144]},
      {stage1_37[110]}
   );
   gpc1_1 gpc1583 (
      {stage0_37[145]},
      {stage1_37[111]}
   );
   gpc1_1 gpc1584 (
      {stage0_37[146]},
      {stage1_37[112]}
   );
   gpc1_1 gpc1585 (
      {stage0_37[147]},
      {stage1_37[113]}
   );
   gpc1_1 gpc1586 (
      {stage0_37[148]},
      {stage1_37[114]}
   );
   gpc1_1 gpc1587 (
      {stage0_37[149]},
      {stage1_37[115]}
   );
   gpc1_1 gpc1588 (
      {stage0_37[150]},
      {stage1_37[116]}
   );
   gpc1_1 gpc1589 (
      {stage0_37[151]},
      {stage1_37[117]}
   );
   gpc1_1 gpc1590 (
      {stage0_37[152]},
      {stage1_37[118]}
   );
   gpc1_1 gpc1591 (
      {stage0_37[153]},
      {stage1_37[119]}
   );
   gpc1_1 gpc1592 (
      {stage0_37[154]},
      {stage1_37[120]}
   );
   gpc1_1 gpc1593 (
      {stage0_37[155]},
      {stage1_37[121]}
   );
   gpc1_1 gpc1594 (
      {stage0_37[156]},
      {stage1_37[122]}
   );
   gpc1_1 gpc1595 (
      {stage0_37[157]},
      {stage1_37[123]}
   );
   gpc1_1 gpc1596 (
      {stage0_37[158]},
      {stage1_37[124]}
   );
   gpc1_1 gpc1597 (
      {stage0_37[159]},
      {stage1_37[125]}
   );
   gpc1_1 gpc1598 (
      {stage0_37[160]},
      {stage1_37[126]}
   );
   gpc1_1 gpc1599 (
      {stage0_37[161]},
      {stage1_37[127]}
   );
   gpc1_1 gpc1600 (
      {stage0_38[148]},
      {stage1_38[52]}
   );
   gpc1_1 gpc1601 (
      {stage0_38[149]},
      {stage1_38[53]}
   );
   gpc1_1 gpc1602 (
      {stage0_38[150]},
      {stage1_38[54]}
   );
   gpc1_1 gpc1603 (
      {stage0_38[151]},
      {stage1_38[55]}
   );
   gpc1_1 gpc1604 (
      {stage0_38[152]},
      {stage1_38[56]}
   );
   gpc1_1 gpc1605 (
      {stage0_38[153]},
      {stage1_38[57]}
   );
   gpc1_1 gpc1606 (
      {stage0_38[154]},
      {stage1_38[58]}
   );
   gpc1_1 gpc1607 (
      {stage0_38[155]},
      {stage1_38[59]}
   );
   gpc1_1 gpc1608 (
      {stage0_38[156]},
      {stage1_38[60]}
   );
   gpc1_1 gpc1609 (
      {stage0_38[157]},
      {stage1_38[61]}
   );
   gpc1_1 gpc1610 (
      {stage0_38[158]},
      {stage1_38[62]}
   );
   gpc1_1 gpc1611 (
      {stage0_38[159]},
      {stage1_38[63]}
   );
   gpc1_1 gpc1612 (
      {stage0_38[160]},
      {stage1_38[64]}
   );
   gpc1_1 gpc1613 (
      {stage0_38[161]},
      {stage1_38[65]}
   );
   gpc1_1 gpc1614 (
      {stage0_39[156]},
      {stage1_39[62]}
   );
   gpc1_1 gpc1615 (
      {stage0_39[157]},
      {stage1_39[63]}
   );
   gpc1_1 gpc1616 (
      {stage0_39[158]},
      {stage1_39[64]}
   );
   gpc1_1 gpc1617 (
      {stage0_39[159]},
      {stage1_39[65]}
   );
   gpc1_1 gpc1618 (
      {stage0_39[160]},
      {stage1_39[66]}
   );
   gpc1_1 gpc1619 (
      {stage0_39[161]},
      {stage1_39[67]}
   );
   gpc1_1 gpc1620 (
      {stage0_40[140]},
      {stage1_40[60]}
   );
   gpc1_1 gpc1621 (
      {stage0_40[141]},
      {stage1_40[61]}
   );
   gpc1_1 gpc1622 (
      {stage0_40[142]},
      {stage1_40[62]}
   );
   gpc1_1 gpc1623 (
      {stage0_40[143]},
      {stage1_40[63]}
   );
   gpc1_1 gpc1624 (
      {stage0_40[144]},
      {stage1_40[64]}
   );
   gpc1_1 gpc1625 (
      {stage0_40[145]},
      {stage1_40[65]}
   );
   gpc1_1 gpc1626 (
      {stage0_40[146]},
      {stage1_40[66]}
   );
   gpc1_1 gpc1627 (
      {stage0_40[147]},
      {stage1_40[67]}
   );
   gpc1_1 gpc1628 (
      {stage0_40[148]},
      {stage1_40[68]}
   );
   gpc1_1 gpc1629 (
      {stage0_40[149]},
      {stage1_40[69]}
   );
   gpc1_1 gpc1630 (
      {stage0_40[150]},
      {stage1_40[70]}
   );
   gpc1_1 gpc1631 (
      {stage0_40[151]},
      {stage1_40[71]}
   );
   gpc1_1 gpc1632 (
      {stage0_40[152]},
      {stage1_40[72]}
   );
   gpc1_1 gpc1633 (
      {stage0_40[153]},
      {stage1_40[73]}
   );
   gpc1_1 gpc1634 (
      {stage0_40[154]},
      {stage1_40[74]}
   );
   gpc1_1 gpc1635 (
      {stage0_40[155]},
      {stage1_40[75]}
   );
   gpc1_1 gpc1636 (
      {stage0_40[156]},
      {stage1_40[76]}
   );
   gpc1_1 gpc1637 (
      {stage0_40[157]},
      {stage1_40[77]}
   );
   gpc1_1 gpc1638 (
      {stage0_40[158]},
      {stage1_40[78]}
   );
   gpc1_1 gpc1639 (
      {stage0_40[159]},
      {stage1_40[79]}
   );
   gpc1_1 gpc1640 (
      {stage0_40[160]},
      {stage1_40[80]}
   );
   gpc1_1 gpc1641 (
      {stage0_40[161]},
      {stage1_40[81]}
   );
   gpc1_1 gpc1642 (
      {stage0_41[138]},
      {stage1_41[50]}
   );
   gpc1_1 gpc1643 (
      {stage0_41[139]},
      {stage1_41[51]}
   );
   gpc1_1 gpc1644 (
      {stage0_41[140]},
      {stage1_41[52]}
   );
   gpc1_1 gpc1645 (
      {stage0_41[141]},
      {stage1_41[53]}
   );
   gpc1_1 gpc1646 (
      {stage0_41[142]},
      {stage1_41[54]}
   );
   gpc1_1 gpc1647 (
      {stage0_41[143]},
      {stage1_41[55]}
   );
   gpc1_1 gpc1648 (
      {stage0_41[144]},
      {stage1_41[56]}
   );
   gpc1_1 gpc1649 (
      {stage0_41[145]},
      {stage1_41[57]}
   );
   gpc1_1 gpc1650 (
      {stage0_41[146]},
      {stage1_41[58]}
   );
   gpc1_1 gpc1651 (
      {stage0_41[147]},
      {stage1_41[59]}
   );
   gpc1_1 gpc1652 (
      {stage0_41[148]},
      {stage1_41[60]}
   );
   gpc1_1 gpc1653 (
      {stage0_41[149]},
      {stage1_41[61]}
   );
   gpc1_1 gpc1654 (
      {stage0_41[150]},
      {stage1_41[62]}
   );
   gpc1_1 gpc1655 (
      {stage0_41[151]},
      {stage1_41[63]}
   );
   gpc1_1 gpc1656 (
      {stage0_41[152]},
      {stage1_41[64]}
   );
   gpc1_1 gpc1657 (
      {stage0_41[153]},
      {stage1_41[65]}
   );
   gpc1_1 gpc1658 (
      {stage0_41[154]},
      {stage1_41[66]}
   );
   gpc1_1 gpc1659 (
      {stage0_41[155]},
      {stage1_41[67]}
   );
   gpc1_1 gpc1660 (
      {stage0_41[156]},
      {stage1_41[68]}
   );
   gpc1_1 gpc1661 (
      {stage0_41[157]},
      {stage1_41[69]}
   );
   gpc1_1 gpc1662 (
      {stage0_41[158]},
      {stage1_41[70]}
   );
   gpc1_1 gpc1663 (
      {stage0_41[159]},
      {stage1_41[71]}
   );
   gpc1_1 gpc1664 (
      {stage0_41[160]},
      {stage1_41[72]}
   );
   gpc1_1 gpc1665 (
      {stage0_41[161]},
      {stage1_41[73]}
   );
   gpc1_1 gpc1666 (
      {stage0_42[126]},
      {stage1_42[60]}
   );
   gpc1_1 gpc1667 (
      {stage0_42[127]},
      {stage1_42[61]}
   );
   gpc1_1 gpc1668 (
      {stage0_42[128]},
      {stage1_42[62]}
   );
   gpc1_1 gpc1669 (
      {stage0_42[129]},
      {stage1_42[63]}
   );
   gpc1_1 gpc1670 (
      {stage0_42[130]},
      {stage1_42[64]}
   );
   gpc1_1 gpc1671 (
      {stage0_42[131]},
      {stage1_42[65]}
   );
   gpc1_1 gpc1672 (
      {stage0_42[132]},
      {stage1_42[66]}
   );
   gpc1_1 gpc1673 (
      {stage0_42[133]},
      {stage1_42[67]}
   );
   gpc1_1 gpc1674 (
      {stage0_42[134]},
      {stage1_42[68]}
   );
   gpc1_1 gpc1675 (
      {stage0_42[135]},
      {stage1_42[69]}
   );
   gpc1_1 gpc1676 (
      {stage0_42[136]},
      {stage1_42[70]}
   );
   gpc1_1 gpc1677 (
      {stage0_42[137]},
      {stage1_42[71]}
   );
   gpc1_1 gpc1678 (
      {stage0_42[138]},
      {stage1_42[72]}
   );
   gpc1_1 gpc1679 (
      {stage0_42[139]},
      {stage1_42[73]}
   );
   gpc1_1 gpc1680 (
      {stage0_42[140]},
      {stage1_42[74]}
   );
   gpc1_1 gpc1681 (
      {stage0_42[141]},
      {stage1_42[75]}
   );
   gpc1_1 gpc1682 (
      {stage0_42[142]},
      {stage1_42[76]}
   );
   gpc1_1 gpc1683 (
      {stage0_42[143]},
      {stage1_42[77]}
   );
   gpc1_1 gpc1684 (
      {stage0_42[144]},
      {stage1_42[78]}
   );
   gpc1_1 gpc1685 (
      {stage0_42[145]},
      {stage1_42[79]}
   );
   gpc1_1 gpc1686 (
      {stage0_42[146]},
      {stage1_42[80]}
   );
   gpc1_1 gpc1687 (
      {stage0_42[147]},
      {stage1_42[81]}
   );
   gpc1_1 gpc1688 (
      {stage0_42[148]},
      {stage1_42[82]}
   );
   gpc1_1 gpc1689 (
      {stage0_42[149]},
      {stage1_42[83]}
   );
   gpc1_1 gpc1690 (
      {stage0_42[150]},
      {stage1_42[84]}
   );
   gpc1_1 gpc1691 (
      {stage0_42[151]},
      {stage1_42[85]}
   );
   gpc1_1 gpc1692 (
      {stage0_42[152]},
      {stage1_42[86]}
   );
   gpc1_1 gpc1693 (
      {stage0_42[153]},
      {stage1_42[87]}
   );
   gpc1_1 gpc1694 (
      {stage0_42[154]},
      {stage1_42[88]}
   );
   gpc1_1 gpc1695 (
      {stage0_42[155]},
      {stage1_42[89]}
   );
   gpc1_1 gpc1696 (
      {stage0_42[156]},
      {stage1_42[90]}
   );
   gpc1_1 gpc1697 (
      {stage0_42[157]},
      {stage1_42[91]}
   );
   gpc1_1 gpc1698 (
      {stage0_42[158]},
      {stage1_42[92]}
   );
   gpc1_1 gpc1699 (
      {stage0_42[159]},
      {stage1_42[93]}
   );
   gpc1_1 gpc1700 (
      {stage0_42[160]},
      {stage1_42[94]}
   );
   gpc1_1 gpc1701 (
      {stage0_42[161]},
      {stage1_42[95]}
   );
   gpc1_1 gpc1702 (
      {stage0_43[78]},
      {stage1_43[54]}
   );
   gpc1_1 gpc1703 (
      {stage0_43[79]},
      {stage1_43[55]}
   );
   gpc1_1 gpc1704 (
      {stage0_43[80]},
      {stage1_43[56]}
   );
   gpc1_1 gpc1705 (
      {stage0_43[81]},
      {stage1_43[57]}
   );
   gpc1_1 gpc1706 (
      {stage0_43[82]},
      {stage1_43[58]}
   );
   gpc1_1 gpc1707 (
      {stage0_43[83]},
      {stage1_43[59]}
   );
   gpc1_1 gpc1708 (
      {stage0_43[84]},
      {stage1_43[60]}
   );
   gpc1_1 gpc1709 (
      {stage0_43[85]},
      {stage1_43[61]}
   );
   gpc1_1 gpc1710 (
      {stage0_43[86]},
      {stage1_43[62]}
   );
   gpc1_1 gpc1711 (
      {stage0_43[87]},
      {stage1_43[63]}
   );
   gpc1_1 gpc1712 (
      {stage0_43[88]},
      {stage1_43[64]}
   );
   gpc1_1 gpc1713 (
      {stage0_43[89]},
      {stage1_43[65]}
   );
   gpc1_1 gpc1714 (
      {stage0_43[90]},
      {stage1_43[66]}
   );
   gpc1_1 gpc1715 (
      {stage0_43[91]},
      {stage1_43[67]}
   );
   gpc1_1 gpc1716 (
      {stage0_43[92]},
      {stage1_43[68]}
   );
   gpc1_1 gpc1717 (
      {stage0_43[93]},
      {stage1_43[69]}
   );
   gpc1_1 gpc1718 (
      {stage0_43[94]},
      {stage1_43[70]}
   );
   gpc1_1 gpc1719 (
      {stage0_43[95]},
      {stage1_43[71]}
   );
   gpc1_1 gpc1720 (
      {stage0_43[96]},
      {stage1_43[72]}
   );
   gpc1_1 gpc1721 (
      {stage0_43[97]},
      {stage1_43[73]}
   );
   gpc1_1 gpc1722 (
      {stage0_43[98]},
      {stage1_43[74]}
   );
   gpc1_1 gpc1723 (
      {stage0_43[99]},
      {stage1_43[75]}
   );
   gpc1_1 gpc1724 (
      {stage0_43[100]},
      {stage1_43[76]}
   );
   gpc1_1 gpc1725 (
      {stage0_43[101]},
      {stage1_43[77]}
   );
   gpc1_1 gpc1726 (
      {stage0_43[102]},
      {stage1_43[78]}
   );
   gpc1_1 gpc1727 (
      {stage0_43[103]},
      {stage1_43[79]}
   );
   gpc1_1 gpc1728 (
      {stage0_43[104]},
      {stage1_43[80]}
   );
   gpc1_1 gpc1729 (
      {stage0_43[105]},
      {stage1_43[81]}
   );
   gpc1_1 gpc1730 (
      {stage0_43[106]},
      {stage1_43[82]}
   );
   gpc1_1 gpc1731 (
      {stage0_43[107]},
      {stage1_43[83]}
   );
   gpc1_1 gpc1732 (
      {stage0_43[108]},
      {stage1_43[84]}
   );
   gpc1_1 gpc1733 (
      {stage0_43[109]},
      {stage1_43[85]}
   );
   gpc1_1 gpc1734 (
      {stage0_43[110]},
      {stage1_43[86]}
   );
   gpc1_1 gpc1735 (
      {stage0_43[111]},
      {stage1_43[87]}
   );
   gpc1_1 gpc1736 (
      {stage0_43[112]},
      {stage1_43[88]}
   );
   gpc1_1 gpc1737 (
      {stage0_43[113]},
      {stage1_43[89]}
   );
   gpc1_1 gpc1738 (
      {stage0_43[114]},
      {stage1_43[90]}
   );
   gpc1_1 gpc1739 (
      {stage0_43[115]},
      {stage1_43[91]}
   );
   gpc1_1 gpc1740 (
      {stage0_43[116]},
      {stage1_43[92]}
   );
   gpc1_1 gpc1741 (
      {stage0_43[117]},
      {stage1_43[93]}
   );
   gpc1_1 gpc1742 (
      {stage0_43[118]},
      {stage1_43[94]}
   );
   gpc1_1 gpc1743 (
      {stage0_43[119]},
      {stage1_43[95]}
   );
   gpc1_1 gpc1744 (
      {stage0_43[120]},
      {stage1_43[96]}
   );
   gpc1_1 gpc1745 (
      {stage0_43[121]},
      {stage1_43[97]}
   );
   gpc1_1 gpc1746 (
      {stage0_43[122]},
      {stage1_43[98]}
   );
   gpc1_1 gpc1747 (
      {stage0_43[123]},
      {stage1_43[99]}
   );
   gpc1_1 gpc1748 (
      {stage0_43[124]},
      {stage1_43[100]}
   );
   gpc1_1 gpc1749 (
      {stage0_43[125]},
      {stage1_43[101]}
   );
   gpc1_1 gpc1750 (
      {stage0_43[126]},
      {stage1_43[102]}
   );
   gpc1_1 gpc1751 (
      {stage0_43[127]},
      {stage1_43[103]}
   );
   gpc1_1 gpc1752 (
      {stage0_43[128]},
      {stage1_43[104]}
   );
   gpc1_1 gpc1753 (
      {stage0_43[129]},
      {stage1_43[105]}
   );
   gpc1_1 gpc1754 (
      {stage0_43[130]},
      {stage1_43[106]}
   );
   gpc1_1 gpc1755 (
      {stage0_43[131]},
      {stage1_43[107]}
   );
   gpc1_1 gpc1756 (
      {stage0_43[132]},
      {stage1_43[108]}
   );
   gpc1_1 gpc1757 (
      {stage0_43[133]},
      {stage1_43[109]}
   );
   gpc1_1 gpc1758 (
      {stage0_43[134]},
      {stage1_43[110]}
   );
   gpc1_1 gpc1759 (
      {stage0_43[135]},
      {stage1_43[111]}
   );
   gpc1_1 gpc1760 (
      {stage0_43[136]},
      {stage1_43[112]}
   );
   gpc1_1 gpc1761 (
      {stage0_43[137]},
      {stage1_43[113]}
   );
   gpc1_1 gpc1762 (
      {stage0_43[138]},
      {stage1_43[114]}
   );
   gpc1_1 gpc1763 (
      {stage0_43[139]},
      {stage1_43[115]}
   );
   gpc1_1 gpc1764 (
      {stage0_43[140]},
      {stage1_43[116]}
   );
   gpc1_1 gpc1765 (
      {stage0_43[141]},
      {stage1_43[117]}
   );
   gpc1_1 gpc1766 (
      {stage0_43[142]},
      {stage1_43[118]}
   );
   gpc1_1 gpc1767 (
      {stage0_43[143]},
      {stage1_43[119]}
   );
   gpc1_1 gpc1768 (
      {stage0_43[144]},
      {stage1_43[120]}
   );
   gpc1_1 gpc1769 (
      {stage0_43[145]},
      {stage1_43[121]}
   );
   gpc1_1 gpc1770 (
      {stage0_43[146]},
      {stage1_43[122]}
   );
   gpc1_1 gpc1771 (
      {stage0_43[147]},
      {stage1_43[123]}
   );
   gpc1_1 gpc1772 (
      {stage0_43[148]},
      {stage1_43[124]}
   );
   gpc1_1 gpc1773 (
      {stage0_43[149]},
      {stage1_43[125]}
   );
   gpc1_1 gpc1774 (
      {stage0_43[150]},
      {stage1_43[126]}
   );
   gpc1_1 gpc1775 (
      {stage0_43[151]},
      {stage1_43[127]}
   );
   gpc1_1 gpc1776 (
      {stage0_43[152]},
      {stage1_43[128]}
   );
   gpc1_1 gpc1777 (
      {stage0_43[153]},
      {stage1_43[129]}
   );
   gpc1_1 gpc1778 (
      {stage0_43[154]},
      {stage1_43[130]}
   );
   gpc1_1 gpc1779 (
      {stage0_43[155]},
      {stage1_43[131]}
   );
   gpc1_1 gpc1780 (
      {stage0_43[156]},
      {stage1_43[132]}
   );
   gpc1_1 gpc1781 (
      {stage0_43[157]},
      {stage1_43[133]}
   );
   gpc1_1 gpc1782 (
      {stage0_43[158]},
      {stage1_43[134]}
   );
   gpc1_1 gpc1783 (
      {stage0_43[159]},
      {stage1_43[135]}
   );
   gpc1_1 gpc1784 (
      {stage0_43[160]},
      {stage1_43[136]}
   );
   gpc1_1 gpc1785 (
      {stage0_43[161]},
      {stage1_43[137]}
   );
   gpc1_1 gpc1786 (
      {stage0_44[160]},
      {stage1_44[44]}
   );
   gpc1_1 gpc1787 (
      {stage0_44[161]},
      {stage1_44[45]}
   );
   gpc1_1 gpc1788 (
      {stage0_45[121]},
      {stage1_45[52]}
   );
   gpc1_1 gpc1789 (
      {stage0_45[122]},
      {stage1_45[53]}
   );
   gpc1_1 gpc1790 (
      {stage0_45[123]},
      {stage1_45[54]}
   );
   gpc1_1 gpc1791 (
      {stage0_45[124]},
      {stage1_45[55]}
   );
   gpc1_1 gpc1792 (
      {stage0_45[125]},
      {stage1_45[56]}
   );
   gpc1_1 gpc1793 (
      {stage0_45[126]},
      {stage1_45[57]}
   );
   gpc1_1 gpc1794 (
      {stage0_45[127]},
      {stage1_45[58]}
   );
   gpc1_1 gpc1795 (
      {stage0_45[128]},
      {stage1_45[59]}
   );
   gpc1_1 gpc1796 (
      {stage0_45[129]},
      {stage1_45[60]}
   );
   gpc1_1 gpc1797 (
      {stage0_45[130]},
      {stage1_45[61]}
   );
   gpc1_1 gpc1798 (
      {stage0_45[131]},
      {stage1_45[62]}
   );
   gpc1_1 gpc1799 (
      {stage0_45[132]},
      {stage1_45[63]}
   );
   gpc1_1 gpc1800 (
      {stage0_45[133]},
      {stage1_45[64]}
   );
   gpc1_1 gpc1801 (
      {stage0_45[134]},
      {stage1_45[65]}
   );
   gpc1_1 gpc1802 (
      {stage0_45[135]},
      {stage1_45[66]}
   );
   gpc1_1 gpc1803 (
      {stage0_45[136]},
      {stage1_45[67]}
   );
   gpc1_1 gpc1804 (
      {stage0_45[137]},
      {stage1_45[68]}
   );
   gpc1_1 gpc1805 (
      {stage0_45[138]},
      {stage1_45[69]}
   );
   gpc1_1 gpc1806 (
      {stage0_45[139]},
      {stage1_45[70]}
   );
   gpc1_1 gpc1807 (
      {stage0_45[140]},
      {stage1_45[71]}
   );
   gpc1_1 gpc1808 (
      {stage0_45[141]},
      {stage1_45[72]}
   );
   gpc1_1 gpc1809 (
      {stage0_45[142]},
      {stage1_45[73]}
   );
   gpc1_1 gpc1810 (
      {stage0_45[143]},
      {stage1_45[74]}
   );
   gpc1_1 gpc1811 (
      {stage0_45[144]},
      {stage1_45[75]}
   );
   gpc1_1 gpc1812 (
      {stage0_45[145]},
      {stage1_45[76]}
   );
   gpc1_1 gpc1813 (
      {stage0_45[146]},
      {stage1_45[77]}
   );
   gpc1_1 gpc1814 (
      {stage0_45[147]},
      {stage1_45[78]}
   );
   gpc1_1 gpc1815 (
      {stage0_45[148]},
      {stage1_45[79]}
   );
   gpc1_1 gpc1816 (
      {stage0_45[149]},
      {stage1_45[80]}
   );
   gpc1_1 gpc1817 (
      {stage0_45[150]},
      {stage1_45[81]}
   );
   gpc1_1 gpc1818 (
      {stage0_45[151]},
      {stage1_45[82]}
   );
   gpc1_1 gpc1819 (
      {stage0_45[152]},
      {stage1_45[83]}
   );
   gpc1_1 gpc1820 (
      {stage0_45[153]},
      {stage1_45[84]}
   );
   gpc1_1 gpc1821 (
      {stage0_45[154]},
      {stage1_45[85]}
   );
   gpc1_1 gpc1822 (
      {stage0_45[155]},
      {stage1_45[86]}
   );
   gpc1_1 gpc1823 (
      {stage0_45[156]},
      {stage1_45[87]}
   );
   gpc1_1 gpc1824 (
      {stage0_45[157]},
      {stage1_45[88]}
   );
   gpc1_1 gpc1825 (
      {stage0_45[158]},
      {stage1_45[89]}
   );
   gpc1_1 gpc1826 (
      {stage0_45[159]},
      {stage1_45[90]}
   );
   gpc1_1 gpc1827 (
      {stage0_45[160]},
      {stage1_45[91]}
   );
   gpc1_1 gpc1828 (
      {stage0_45[161]},
      {stage1_45[92]}
   );
   gpc1_1 gpc1829 (
      {stage0_46[161]},
      {stage1_46[63]}
   );
   gpc1_1 gpc1830 (
      {stage0_48[161]},
      {stage1_48[71]}
   );
   gpc1_1 gpc1831 (
      {stage0_49[147]},
      {stage1_49[72]}
   );
   gpc1_1 gpc1832 (
      {stage0_49[148]},
      {stage1_49[73]}
   );
   gpc1_1 gpc1833 (
      {stage0_49[149]},
      {stage1_49[74]}
   );
   gpc1_1 gpc1834 (
      {stage0_49[150]},
      {stage1_49[75]}
   );
   gpc1_1 gpc1835 (
      {stage0_49[151]},
      {stage1_49[76]}
   );
   gpc1_1 gpc1836 (
      {stage0_49[152]},
      {stage1_49[77]}
   );
   gpc1_1 gpc1837 (
      {stage0_49[153]},
      {stage1_49[78]}
   );
   gpc1_1 gpc1838 (
      {stage0_49[154]},
      {stage1_49[79]}
   );
   gpc1_1 gpc1839 (
      {stage0_49[155]},
      {stage1_49[80]}
   );
   gpc1_1 gpc1840 (
      {stage0_49[156]},
      {stage1_49[81]}
   );
   gpc1_1 gpc1841 (
      {stage0_49[157]},
      {stage1_49[82]}
   );
   gpc1_1 gpc1842 (
      {stage0_49[158]},
      {stage1_49[83]}
   );
   gpc1_1 gpc1843 (
      {stage0_49[159]},
      {stage1_49[84]}
   );
   gpc1_1 gpc1844 (
      {stage0_49[160]},
      {stage1_49[85]}
   );
   gpc1_1 gpc1845 (
      {stage0_49[161]},
      {stage1_49[86]}
   );
   gpc1_1 gpc1846 (
      {stage0_50[159]},
      {stage1_50[55]}
   );
   gpc1_1 gpc1847 (
      {stage0_50[160]},
      {stage1_50[56]}
   );
   gpc1_1 gpc1848 (
      {stage0_50[161]},
      {stage1_50[57]}
   );
   gpc1_1 gpc1849 (
      {stage0_51[126]},
      {stage1_51[58]}
   );
   gpc1_1 gpc1850 (
      {stage0_51[127]},
      {stage1_51[59]}
   );
   gpc1_1 gpc1851 (
      {stage0_51[128]},
      {stage1_51[60]}
   );
   gpc1_1 gpc1852 (
      {stage0_51[129]},
      {stage1_51[61]}
   );
   gpc1_1 gpc1853 (
      {stage0_51[130]},
      {stage1_51[62]}
   );
   gpc1_1 gpc1854 (
      {stage0_51[131]},
      {stage1_51[63]}
   );
   gpc1_1 gpc1855 (
      {stage0_51[132]},
      {stage1_51[64]}
   );
   gpc1_1 gpc1856 (
      {stage0_51[133]},
      {stage1_51[65]}
   );
   gpc1_1 gpc1857 (
      {stage0_51[134]},
      {stage1_51[66]}
   );
   gpc1_1 gpc1858 (
      {stage0_51[135]},
      {stage1_51[67]}
   );
   gpc1_1 gpc1859 (
      {stage0_51[136]},
      {stage1_51[68]}
   );
   gpc1_1 gpc1860 (
      {stage0_51[137]},
      {stage1_51[69]}
   );
   gpc1_1 gpc1861 (
      {stage0_51[138]},
      {stage1_51[70]}
   );
   gpc1_1 gpc1862 (
      {stage0_51[139]},
      {stage1_51[71]}
   );
   gpc1_1 gpc1863 (
      {stage0_51[140]},
      {stage1_51[72]}
   );
   gpc1_1 gpc1864 (
      {stage0_51[141]},
      {stage1_51[73]}
   );
   gpc1_1 gpc1865 (
      {stage0_51[142]},
      {stage1_51[74]}
   );
   gpc1_1 gpc1866 (
      {stage0_51[143]},
      {stage1_51[75]}
   );
   gpc1_1 gpc1867 (
      {stage0_51[144]},
      {stage1_51[76]}
   );
   gpc1_1 gpc1868 (
      {stage0_51[145]},
      {stage1_51[77]}
   );
   gpc1_1 gpc1869 (
      {stage0_51[146]},
      {stage1_51[78]}
   );
   gpc1_1 gpc1870 (
      {stage0_51[147]},
      {stage1_51[79]}
   );
   gpc1_1 gpc1871 (
      {stage0_51[148]},
      {stage1_51[80]}
   );
   gpc1_1 gpc1872 (
      {stage0_51[149]},
      {stage1_51[81]}
   );
   gpc1_1 gpc1873 (
      {stage0_51[150]},
      {stage1_51[82]}
   );
   gpc1_1 gpc1874 (
      {stage0_51[151]},
      {stage1_51[83]}
   );
   gpc1_1 gpc1875 (
      {stage0_51[152]},
      {stage1_51[84]}
   );
   gpc1_1 gpc1876 (
      {stage0_51[153]},
      {stage1_51[85]}
   );
   gpc1_1 gpc1877 (
      {stage0_51[154]},
      {stage1_51[86]}
   );
   gpc1_1 gpc1878 (
      {stage0_51[155]},
      {stage1_51[87]}
   );
   gpc1_1 gpc1879 (
      {stage0_51[156]},
      {stage1_51[88]}
   );
   gpc1_1 gpc1880 (
      {stage0_51[157]},
      {stage1_51[89]}
   );
   gpc1_1 gpc1881 (
      {stage0_51[158]},
      {stage1_51[90]}
   );
   gpc1_1 gpc1882 (
      {stage0_51[159]},
      {stage1_51[91]}
   );
   gpc1_1 gpc1883 (
      {stage0_51[160]},
      {stage1_51[92]}
   );
   gpc1_1 gpc1884 (
      {stage0_51[161]},
      {stage1_51[93]}
   );
   gpc1_1 gpc1885 (
      {stage0_52[153]},
      {stage1_52[68]}
   );
   gpc1_1 gpc1886 (
      {stage0_52[154]},
      {stage1_52[69]}
   );
   gpc1_1 gpc1887 (
      {stage0_52[155]},
      {stage1_52[70]}
   );
   gpc1_1 gpc1888 (
      {stage0_52[156]},
      {stage1_52[71]}
   );
   gpc1_1 gpc1889 (
      {stage0_52[157]},
      {stage1_52[72]}
   );
   gpc1_1 gpc1890 (
      {stage0_52[158]},
      {stage1_52[73]}
   );
   gpc1_1 gpc1891 (
      {stage0_52[159]},
      {stage1_52[74]}
   );
   gpc1_1 gpc1892 (
      {stage0_52[160]},
      {stage1_52[75]}
   );
   gpc1_1 gpc1893 (
      {stage0_52[161]},
      {stage1_52[76]}
   );
   gpc1_1 gpc1894 (
      {stage0_53[159]},
      {stage1_53[63]}
   );
   gpc1_1 gpc1895 (
      {stage0_53[160]},
      {stage1_53[64]}
   );
   gpc1_1 gpc1896 (
      {stage0_53[161]},
      {stage1_53[65]}
   );
   gpc1_1 gpc1897 (
      {stage0_55[122]},
      {stage1_55[58]}
   );
   gpc1_1 gpc1898 (
      {stage0_55[123]},
      {stage1_55[59]}
   );
   gpc1_1 gpc1899 (
      {stage0_55[124]},
      {stage1_55[60]}
   );
   gpc1_1 gpc1900 (
      {stage0_55[125]},
      {stage1_55[61]}
   );
   gpc1_1 gpc1901 (
      {stage0_55[126]},
      {stage1_55[62]}
   );
   gpc1_1 gpc1902 (
      {stage0_55[127]},
      {stage1_55[63]}
   );
   gpc1_1 gpc1903 (
      {stage0_55[128]},
      {stage1_55[64]}
   );
   gpc1_1 gpc1904 (
      {stage0_55[129]},
      {stage1_55[65]}
   );
   gpc1_1 gpc1905 (
      {stage0_55[130]},
      {stage1_55[66]}
   );
   gpc1_1 gpc1906 (
      {stage0_55[131]},
      {stage1_55[67]}
   );
   gpc1_1 gpc1907 (
      {stage0_55[132]},
      {stage1_55[68]}
   );
   gpc1_1 gpc1908 (
      {stage0_55[133]},
      {stage1_55[69]}
   );
   gpc1_1 gpc1909 (
      {stage0_55[134]},
      {stage1_55[70]}
   );
   gpc1_1 gpc1910 (
      {stage0_55[135]},
      {stage1_55[71]}
   );
   gpc1_1 gpc1911 (
      {stage0_55[136]},
      {stage1_55[72]}
   );
   gpc1_1 gpc1912 (
      {stage0_55[137]},
      {stage1_55[73]}
   );
   gpc1_1 gpc1913 (
      {stage0_55[138]},
      {stage1_55[74]}
   );
   gpc1_1 gpc1914 (
      {stage0_55[139]},
      {stage1_55[75]}
   );
   gpc1_1 gpc1915 (
      {stage0_55[140]},
      {stage1_55[76]}
   );
   gpc1_1 gpc1916 (
      {stage0_55[141]},
      {stage1_55[77]}
   );
   gpc1_1 gpc1917 (
      {stage0_55[142]},
      {stage1_55[78]}
   );
   gpc1_1 gpc1918 (
      {stage0_55[143]},
      {stage1_55[79]}
   );
   gpc1_1 gpc1919 (
      {stage0_55[144]},
      {stage1_55[80]}
   );
   gpc1_1 gpc1920 (
      {stage0_55[145]},
      {stage1_55[81]}
   );
   gpc1_1 gpc1921 (
      {stage0_55[146]},
      {stage1_55[82]}
   );
   gpc1_1 gpc1922 (
      {stage0_55[147]},
      {stage1_55[83]}
   );
   gpc1_1 gpc1923 (
      {stage0_55[148]},
      {stage1_55[84]}
   );
   gpc1_1 gpc1924 (
      {stage0_55[149]},
      {stage1_55[85]}
   );
   gpc1_1 gpc1925 (
      {stage0_55[150]},
      {stage1_55[86]}
   );
   gpc1_1 gpc1926 (
      {stage0_55[151]},
      {stage1_55[87]}
   );
   gpc1_1 gpc1927 (
      {stage0_55[152]},
      {stage1_55[88]}
   );
   gpc1_1 gpc1928 (
      {stage0_55[153]},
      {stage1_55[89]}
   );
   gpc1_1 gpc1929 (
      {stage0_55[154]},
      {stage1_55[90]}
   );
   gpc1_1 gpc1930 (
      {stage0_55[155]},
      {stage1_55[91]}
   );
   gpc1_1 gpc1931 (
      {stage0_55[156]},
      {stage1_55[92]}
   );
   gpc1_1 gpc1932 (
      {stage0_55[157]},
      {stage1_55[93]}
   );
   gpc1_1 gpc1933 (
      {stage0_55[158]},
      {stage1_55[94]}
   );
   gpc1_1 gpc1934 (
      {stage0_55[159]},
      {stage1_55[95]}
   );
   gpc1_1 gpc1935 (
      {stage0_55[160]},
      {stage1_55[96]}
   );
   gpc1_1 gpc1936 (
      {stage0_55[161]},
      {stage1_55[97]}
   );
   gpc1_1 gpc1937 (
      {stage0_56[148]},
      {stage1_56[66]}
   );
   gpc1_1 gpc1938 (
      {stage0_56[149]},
      {stage1_56[67]}
   );
   gpc1_1 gpc1939 (
      {stage0_56[150]},
      {stage1_56[68]}
   );
   gpc1_1 gpc1940 (
      {stage0_56[151]},
      {stage1_56[69]}
   );
   gpc1_1 gpc1941 (
      {stage0_56[152]},
      {stage1_56[70]}
   );
   gpc1_1 gpc1942 (
      {stage0_56[153]},
      {stage1_56[71]}
   );
   gpc1_1 gpc1943 (
      {stage0_56[154]},
      {stage1_56[72]}
   );
   gpc1_1 gpc1944 (
      {stage0_56[155]},
      {stage1_56[73]}
   );
   gpc1_1 gpc1945 (
      {stage0_56[156]},
      {stage1_56[74]}
   );
   gpc1_1 gpc1946 (
      {stage0_56[157]},
      {stage1_56[75]}
   );
   gpc1_1 gpc1947 (
      {stage0_56[158]},
      {stage1_56[76]}
   );
   gpc1_1 gpc1948 (
      {stage0_56[159]},
      {stage1_56[77]}
   );
   gpc1_1 gpc1949 (
      {stage0_56[160]},
      {stage1_56[78]}
   );
   gpc1_1 gpc1950 (
      {stage0_56[161]},
      {stage1_56[79]}
   );
   gpc1_1 gpc1951 (
      {stage0_57[156]},
      {stage1_57[66]}
   );
   gpc1_1 gpc1952 (
      {stage0_57[157]},
      {stage1_57[67]}
   );
   gpc1_1 gpc1953 (
      {stage0_57[158]},
      {stage1_57[68]}
   );
   gpc1_1 gpc1954 (
      {stage0_57[159]},
      {stage1_57[69]}
   );
   gpc1_1 gpc1955 (
      {stage0_57[160]},
      {stage1_57[70]}
   );
   gpc1_1 gpc1956 (
      {stage0_57[161]},
      {stage1_57[71]}
   );
   gpc1_1 gpc1957 (
      {stage0_58[144]},
      {stage1_58[56]}
   );
   gpc1_1 gpc1958 (
      {stage0_58[145]},
      {stage1_58[57]}
   );
   gpc1_1 gpc1959 (
      {stage0_58[146]},
      {stage1_58[58]}
   );
   gpc1_1 gpc1960 (
      {stage0_58[147]},
      {stage1_58[59]}
   );
   gpc1_1 gpc1961 (
      {stage0_58[148]},
      {stage1_58[60]}
   );
   gpc1_1 gpc1962 (
      {stage0_58[149]},
      {stage1_58[61]}
   );
   gpc1_1 gpc1963 (
      {stage0_58[150]},
      {stage1_58[62]}
   );
   gpc1_1 gpc1964 (
      {stage0_58[151]},
      {stage1_58[63]}
   );
   gpc1_1 gpc1965 (
      {stage0_58[152]},
      {stage1_58[64]}
   );
   gpc1_1 gpc1966 (
      {stage0_58[153]},
      {stage1_58[65]}
   );
   gpc1_1 gpc1967 (
      {stage0_58[154]},
      {stage1_58[66]}
   );
   gpc1_1 gpc1968 (
      {stage0_58[155]},
      {stage1_58[67]}
   );
   gpc1_1 gpc1969 (
      {stage0_58[156]},
      {stage1_58[68]}
   );
   gpc1_1 gpc1970 (
      {stage0_58[157]},
      {stage1_58[69]}
   );
   gpc1_1 gpc1971 (
      {stage0_58[158]},
      {stage1_58[70]}
   );
   gpc1_1 gpc1972 (
      {stage0_58[159]},
      {stage1_58[71]}
   );
   gpc1_1 gpc1973 (
      {stage0_58[160]},
      {stage1_58[72]}
   );
   gpc1_1 gpc1974 (
      {stage0_58[161]},
      {stage1_58[73]}
   );
   gpc1_1 gpc1975 (
      {stage0_59[132]},
      {stage1_59[50]}
   );
   gpc1_1 gpc1976 (
      {stage0_59[133]},
      {stage1_59[51]}
   );
   gpc1_1 gpc1977 (
      {stage0_59[134]},
      {stage1_59[52]}
   );
   gpc1_1 gpc1978 (
      {stage0_59[135]},
      {stage1_59[53]}
   );
   gpc1_1 gpc1979 (
      {stage0_59[136]},
      {stage1_59[54]}
   );
   gpc1_1 gpc1980 (
      {stage0_59[137]},
      {stage1_59[55]}
   );
   gpc1_1 gpc1981 (
      {stage0_59[138]},
      {stage1_59[56]}
   );
   gpc1_1 gpc1982 (
      {stage0_59[139]},
      {stage1_59[57]}
   );
   gpc1_1 gpc1983 (
      {stage0_59[140]},
      {stage1_59[58]}
   );
   gpc1_1 gpc1984 (
      {stage0_59[141]},
      {stage1_59[59]}
   );
   gpc1_1 gpc1985 (
      {stage0_59[142]},
      {stage1_59[60]}
   );
   gpc1_1 gpc1986 (
      {stage0_59[143]},
      {stage1_59[61]}
   );
   gpc1_1 gpc1987 (
      {stage0_59[144]},
      {stage1_59[62]}
   );
   gpc1_1 gpc1988 (
      {stage0_59[145]},
      {stage1_59[63]}
   );
   gpc1_1 gpc1989 (
      {stage0_59[146]},
      {stage1_59[64]}
   );
   gpc1_1 gpc1990 (
      {stage0_59[147]},
      {stage1_59[65]}
   );
   gpc1_1 gpc1991 (
      {stage0_59[148]},
      {stage1_59[66]}
   );
   gpc1_1 gpc1992 (
      {stage0_59[149]},
      {stage1_59[67]}
   );
   gpc1_1 gpc1993 (
      {stage0_59[150]},
      {stage1_59[68]}
   );
   gpc1_1 gpc1994 (
      {stage0_59[151]},
      {stage1_59[69]}
   );
   gpc1_1 gpc1995 (
      {stage0_59[152]},
      {stage1_59[70]}
   );
   gpc1_1 gpc1996 (
      {stage0_59[153]},
      {stage1_59[71]}
   );
   gpc1_1 gpc1997 (
      {stage0_59[154]},
      {stage1_59[72]}
   );
   gpc1_1 gpc1998 (
      {stage0_59[155]},
      {stage1_59[73]}
   );
   gpc1_1 gpc1999 (
      {stage0_59[156]},
      {stage1_59[74]}
   );
   gpc1_1 gpc2000 (
      {stage0_59[157]},
      {stage1_59[75]}
   );
   gpc1_1 gpc2001 (
      {stage0_59[158]},
      {stage1_59[76]}
   );
   gpc1_1 gpc2002 (
      {stage0_59[159]},
      {stage1_59[77]}
   );
   gpc1_1 gpc2003 (
      {stage0_59[160]},
      {stage1_59[78]}
   );
   gpc1_1 gpc2004 (
      {stage0_59[161]},
      {stage1_59[79]}
   );
   gpc1_1 gpc2005 (
      {stage0_61[144]},
      {stage1_61[73]}
   );
   gpc1_1 gpc2006 (
      {stage0_61[145]},
      {stage1_61[74]}
   );
   gpc1_1 gpc2007 (
      {stage0_61[146]},
      {stage1_61[75]}
   );
   gpc1_1 gpc2008 (
      {stage0_61[147]},
      {stage1_61[76]}
   );
   gpc1_1 gpc2009 (
      {stage0_61[148]},
      {stage1_61[77]}
   );
   gpc1_1 gpc2010 (
      {stage0_61[149]},
      {stage1_61[78]}
   );
   gpc1_1 gpc2011 (
      {stage0_61[150]},
      {stage1_61[79]}
   );
   gpc1_1 gpc2012 (
      {stage0_61[151]},
      {stage1_61[80]}
   );
   gpc1_1 gpc2013 (
      {stage0_61[152]},
      {stage1_61[81]}
   );
   gpc1_1 gpc2014 (
      {stage0_61[153]},
      {stage1_61[82]}
   );
   gpc1_1 gpc2015 (
      {stage0_61[154]},
      {stage1_61[83]}
   );
   gpc1_1 gpc2016 (
      {stage0_61[155]},
      {stage1_61[84]}
   );
   gpc1_1 gpc2017 (
      {stage0_61[156]},
      {stage1_61[85]}
   );
   gpc1_1 gpc2018 (
      {stage0_61[157]},
      {stage1_61[86]}
   );
   gpc1_1 gpc2019 (
      {stage0_61[158]},
      {stage1_61[87]}
   );
   gpc1_1 gpc2020 (
      {stage0_61[159]},
      {stage1_61[88]}
   );
   gpc1_1 gpc2021 (
      {stage0_61[160]},
      {stage1_61[89]}
   );
   gpc1_1 gpc2022 (
      {stage0_61[161]},
      {stage1_61[90]}
   );
   gpc1_1 gpc2023 (
      {stage0_62[126]},
      {stage1_62[51]}
   );
   gpc1_1 gpc2024 (
      {stage0_62[127]},
      {stage1_62[52]}
   );
   gpc1_1 gpc2025 (
      {stage0_62[128]},
      {stage1_62[53]}
   );
   gpc1_1 gpc2026 (
      {stage0_62[129]},
      {stage1_62[54]}
   );
   gpc1_1 gpc2027 (
      {stage0_62[130]},
      {stage1_62[55]}
   );
   gpc1_1 gpc2028 (
      {stage0_62[131]},
      {stage1_62[56]}
   );
   gpc1_1 gpc2029 (
      {stage0_62[132]},
      {stage1_62[57]}
   );
   gpc1_1 gpc2030 (
      {stage0_62[133]},
      {stage1_62[58]}
   );
   gpc1_1 gpc2031 (
      {stage0_62[134]},
      {stage1_62[59]}
   );
   gpc1_1 gpc2032 (
      {stage0_62[135]},
      {stage1_62[60]}
   );
   gpc1_1 gpc2033 (
      {stage0_62[136]},
      {stage1_62[61]}
   );
   gpc1_1 gpc2034 (
      {stage0_62[137]},
      {stage1_62[62]}
   );
   gpc1_1 gpc2035 (
      {stage0_62[138]},
      {stage1_62[63]}
   );
   gpc1_1 gpc2036 (
      {stage0_62[139]},
      {stage1_62[64]}
   );
   gpc1_1 gpc2037 (
      {stage0_62[140]},
      {stage1_62[65]}
   );
   gpc1_1 gpc2038 (
      {stage0_62[141]},
      {stage1_62[66]}
   );
   gpc1_1 gpc2039 (
      {stage0_62[142]},
      {stage1_62[67]}
   );
   gpc1_1 gpc2040 (
      {stage0_62[143]},
      {stage1_62[68]}
   );
   gpc1_1 gpc2041 (
      {stage0_62[144]},
      {stage1_62[69]}
   );
   gpc1_1 gpc2042 (
      {stage0_62[145]},
      {stage1_62[70]}
   );
   gpc1_1 gpc2043 (
      {stage0_62[146]},
      {stage1_62[71]}
   );
   gpc1_1 gpc2044 (
      {stage0_62[147]},
      {stage1_62[72]}
   );
   gpc1_1 gpc2045 (
      {stage0_62[148]},
      {stage1_62[73]}
   );
   gpc1_1 gpc2046 (
      {stage0_62[149]},
      {stage1_62[74]}
   );
   gpc1_1 gpc2047 (
      {stage0_62[150]},
      {stage1_62[75]}
   );
   gpc1_1 gpc2048 (
      {stage0_62[151]},
      {stage1_62[76]}
   );
   gpc1_1 gpc2049 (
      {stage0_62[152]},
      {stage1_62[77]}
   );
   gpc1_1 gpc2050 (
      {stage0_62[153]},
      {stage1_62[78]}
   );
   gpc1_1 gpc2051 (
      {stage0_62[154]},
      {stage1_62[79]}
   );
   gpc1_1 gpc2052 (
      {stage0_62[155]},
      {stage1_62[80]}
   );
   gpc1_1 gpc2053 (
      {stage0_62[156]},
      {stage1_62[81]}
   );
   gpc1_1 gpc2054 (
      {stage0_62[157]},
      {stage1_62[82]}
   );
   gpc1_1 gpc2055 (
      {stage0_62[158]},
      {stage1_62[83]}
   );
   gpc1_1 gpc2056 (
      {stage0_62[159]},
      {stage1_62[84]}
   );
   gpc1_1 gpc2057 (
      {stage0_62[160]},
      {stage1_62[85]}
   );
   gpc1_1 gpc2058 (
      {stage0_62[161]},
      {stage1_62[86]}
   );
   gpc1_1 gpc2059 (
      {stage0_63[144]},
      {stage1_63[45]}
   );
   gpc1_1 gpc2060 (
      {stage0_63[145]},
      {stage1_63[46]}
   );
   gpc1_1 gpc2061 (
      {stage0_63[146]},
      {stage1_63[47]}
   );
   gpc1_1 gpc2062 (
      {stage0_63[147]},
      {stage1_63[48]}
   );
   gpc1_1 gpc2063 (
      {stage0_63[148]},
      {stage1_63[49]}
   );
   gpc1_1 gpc2064 (
      {stage0_63[149]},
      {stage1_63[50]}
   );
   gpc1_1 gpc2065 (
      {stage0_63[150]},
      {stage1_63[51]}
   );
   gpc1_1 gpc2066 (
      {stage0_63[151]},
      {stage1_63[52]}
   );
   gpc1_1 gpc2067 (
      {stage0_63[152]},
      {stage1_63[53]}
   );
   gpc1_1 gpc2068 (
      {stage0_63[153]},
      {stage1_63[54]}
   );
   gpc1_1 gpc2069 (
      {stage0_63[154]},
      {stage1_63[55]}
   );
   gpc1_1 gpc2070 (
      {stage0_63[155]},
      {stage1_63[56]}
   );
   gpc1_1 gpc2071 (
      {stage0_63[156]},
      {stage1_63[57]}
   );
   gpc1_1 gpc2072 (
      {stage0_63[157]},
      {stage1_63[58]}
   );
   gpc1_1 gpc2073 (
      {stage0_63[158]},
      {stage1_63[59]}
   );
   gpc1_1 gpc2074 (
      {stage0_63[159]},
      {stage1_63[60]}
   );
   gpc1_1 gpc2075 (
      {stage0_63[160]},
      {stage1_63[61]}
   );
   gpc1_1 gpc2076 (
      {stage0_63[161]},
      {stage1_63[62]}
   );
   gpc1163_5 gpc2077 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc2078 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc2079 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2080 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2081 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2082 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_1[18]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2083 (
      {stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30]},
      {stage1_1[19]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2084 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc2085 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc2086 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc1163_5 gpc2087 (
      {stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_5[0]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[0],stage2_5[3],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc2088 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[6]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[1],stage2_6[1],stage2_5[4],stage2_4[11],stage2_3[11]}
   );
   gpc615_5 gpc2089 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[7]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[2],stage2_6[2],stage2_5[5],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc2090 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[8]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[3],stage2_6[3],stage2_5[6],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc2091 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[9]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[4],stage2_6[4],stage2_5[7],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc2092 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[10]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[5],stage2_6[5],stage2_5[8],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc2093 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[11]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[6],stage2_6[6],stage2_5[9],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc2094 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[12]},
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage2_7[7],stage2_6[7],stage2_5[10],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc2095 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[13]},
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage2_7[8],stage2_6[8],stage2_5[11],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc2096 (
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68]},
      {stage1_4[14]},
      {stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54]},
      {stage2_7[9],stage2_6[9],stage2_5[12],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc2097 (
      {stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage1_4[15]},
      {stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60]},
      {stage2_7[10],stage2_6[10],stage2_5[13],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc2098 (
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78]},
      {stage1_4[16]},
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage2_7[11],stage2_6[11],stage2_5[14],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc2099 (
      {stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage1_4[17]},
      {stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72]},
      {stage2_7[12],stage2_6[12],stage2_5[15],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc2100 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[0],stage2_7[13],stage2_6[13],stage2_5[16],stage2_4[23]}
   );
   gpc606_5 gpc2101 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[1],stage2_7[14],stage2_6[14],stage2_5[17],stage2_4[24]}
   );
   gpc606_5 gpc2102 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[2],stage2_7[15],stage2_6[15],stage2_5[18],stage2_4[25]}
   );
   gpc606_5 gpc2103 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[3],stage2_7[16],stage2_6[16],stage2_5[19],stage2_4[26]}
   );
   gpc606_5 gpc2104 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[4],stage2_7[17],stage2_6[17],stage2_5[20],stage2_4[27]}
   );
   gpc606_5 gpc2105 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[5],stage2_7[18],stage2_6[18],stage2_5[21],stage2_4[28]}
   );
   gpc606_5 gpc2106 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[6],stage2_7[19],stage2_6[19],stage2_5[22],stage2_4[29]}
   );
   gpc606_5 gpc2107 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[7],stage2_7[20],stage2_6[20],stage2_5[23],stage2_4[30]}
   );
   gpc606_5 gpc2108 (
      {stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[8],stage2_7[21],stage2_6[21],stage2_5[24]}
   );
   gpc606_5 gpc2109 (
      {stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[9],stage2_7[22],stage2_6[22],stage2_5[25]}
   );
   gpc606_5 gpc2110 (
      {stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[10],stage2_7[23],stage2_6[23],stage2_5[26]}
   );
   gpc606_5 gpc2111 (
      {stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[11],stage2_7[24],stage2_6[24],stage2_5[27]}
   );
   gpc606_5 gpc2112 (
      {stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[12],stage2_7[25],stage2_6[25],stage2_5[28]}
   );
   gpc606_5 gpc2113 (
      {stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[13],stage2_7[26],stage2_6[26],stage2_5[29]}
   );
   gpc615_5 gpc2114 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_7[36]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[6],stage2_8[14],stage2_7[27],stage2_6[27]}
   );
   gpc615_5 gpc2115 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], 1'b0},
      {stage1_7[37]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[7],stage2_8[15],stage2_7[28],stage2_6[28]}
   );
   gpc606_5 gpc2116 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[8],stage2_8[16],stage2_7[29]}
   );
   gpc615_5 gpc2117 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[12]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[9],stage2_8[17],stage2_7[30]}
   );
   gpc615_5 gpc2118 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[13]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[4],stage2_9[10],stage2_8[18],stage2_7[31]}
   );
   gpc615_5 gpc2119 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[14]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[5],stage2_9[11],stage2_8[19],stage2_7[32]}
   );
   gpc615_5 gpc2120 (
      {stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63]},
      {stage1_8[15]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[6],stage2_9[12],stage2_8[20],stage2_7[33]}
   );
   gpc606_5 gpc2121 (
      {stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[5],stage2_10[7],stage2_9[13],stage2_8[21]}
   );
   gpc606_5 gpc2122 (
      {stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[6],stage2_10[8],stage2_9[14],stage2_8[22]}
   );
   gpc606_5 gpc2123 (
      {stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[7],stage2_10[9],stage2_9[15],stage2_8[23]}
   );
   gpc606_5 gpc2124 (
      {stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[8],stage2_10[10],stage2_9[16],stage2_8[24]}
   );
   gpc606_5 gpc2125 (
      {stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[9],stage2_10[11],stage2_9[17],stage2_8[25]}
   );
   gpc606_5 gpc2126 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[10],stage2_10[12],stage2_9[18]}
   );
   gpc606_5 gpc2127 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[11],stage2_10[13],stage2_9[19]}
   );
   gpc606_5 gpc2128 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[12],stage2_10[14],stage2_9[20]}
   );
   gpc606_5 gpc2129 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[13],stage2_10[15],stage2_9[21]}
   );
   gpc606_5 gpc2130 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[14],stage2_10[16]}
   );
   gpc606_5 gpc2131 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[15],stage2_10[17]}
   );
   gpc606_5 gpc2132 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[16],stage2_10[18]}
   );
   gpc606_5 gpc2133 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[17],stage2_10[19]}
   );
   gpc615_5 gpc2134 (
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58]},
      {stage1_11[24]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[18],stage2_10[20]}
   );
   gpc615_5 gpc2135 (
      {stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63]},
      {stage1_11[25]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[19],stage2_10[21]}
   );
   gpc615_5 gpc2136 (
      {stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_11[26]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[20],stage2_10[22]}
   );
   gpc615_5 gpc2137 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage1_11[27]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[21],stage2_10[23]}
   );
   gpc615_5 gpc2138 (
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[28]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[22],stage2_10[24]}
   );
   gpc615_5 gpc2139 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[54]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[23]}
   );
   gpc615_5 gpc2140 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[55]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[24]}
   );
   gpc615_5 gpc2141 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[56]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[25]}
   );
   gpc615_5 gpc2142 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[57]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[26]}
   );
   gpc615_5 gpc2143 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[58]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[13],stage2_13[17],stage2_12[22],stage2_11[27]}
   );
   gpc615_5 gpc2144 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[59]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[14],stage2_13[18],stage2_12[23],stage2_11[28]}
   );
   gpc615_5 gpc2145 (
      {stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63]},
      {stage1_12[60]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[15],stage2_13[19],stage2_12[24],stage2_11[29]}
   );
   gpc615_5 gpc2146 (
      {stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67], stage1_11[68]},
      {stage1_12[61]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[16],stage2_13[20],stage2_12[25],stage2_11[30]}
   );
   gpc615_5 gpc2147 (
      {stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72], stage1_11[73]},
      {stage1_12[62]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[17],stage2_13[21],stage2_12[26],stage2_11[31]}
   );
   gpc606_5 gpc2148 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[9],stage2_14[18],stage2_13[22]}
   );
   gpc606_5 gpc2149 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[10],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc2150 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4]},
      {stage1_15[12]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[11],stage2_14[20]}
   );
   gpc615_5 gpc2151 (
      {stage1_14[5], stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[13]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[12],stage2_14[21]}
   );
   gpc606_5 gpc2152 (
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[13]}
   );
   gpc606_5 gpc2153 (
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[14]}
   );
   gpc606_5 gpc2154 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[6],stage2_15[15]}
   );
   gpc606_5 gpc2155 (
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[7],stage2_15[16]}
   );
   gpc606_5 gpc2156 (
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[8],stage2_15[17]}
   );
   gpc606_5 gpc2157 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[9],stage2_15[18]}
   );
   gpc606_5 gpc2158 (
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[10],stage2_15[19]}
   );
   gpc606_5 gpc2159 (
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[11],stage2_16[11],stage2_15[20]}
   );
   gpc606_5 gpc2160 (
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[12],stage2_16[12],stage2_15[21]}
   );
   gpc606_5 gpc2161 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[13],stage2_16[13],stage2_15[22]}
   );
   gpc606_5 gpc2162 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[14],stage2_16[14],stage2_15[23]}
   );
   gpc606_5 gpc2163 (
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[15],stage2_16[15],stage2_15[24]}
   );
   gpc606_5 gpc2164 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[14],stage2_17[16],stage2_16[16]}
   );
   gpc606_5 gpc2165 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[15],stage2_17[17],stage2_16[17]}
   );
   gpc606_5 gpc2166 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[16],stage2_17[18],stage2_16[18]}
   );
   gpc606_5 gpc2167 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[17],stage2_17[19],stage2_16[19]}
   );
   gpc606_5 gpc2168 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[18],stage2_17[20],stage2_16[20]}
   );
   gpc606_5 gpc2169 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[5],stage2_19[17],stage2_18[19],stage2_17[21]}
   );
   gpc606_5 gpc2170 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[6],stage2_19[18],stage2_18[20],stage2_17[22]}
   );
   gpc606_5 gpc2171 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[7],stage2_19[19],stage2_18[21],stage2_17[23]}
   );
   gpc615_5 gpc2172 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94]},
      {stage1_18[30]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[8],stage2_19[20],stage2_18[22],stage2_17[24]}
   );
   gpc615_5 gpc2173 (
      {stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_18[31]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[9],stage2_19[21],stage2_18[23],stage2_17[25]}
   );
   gpc615_5 gpc2174 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage1_19[30]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[5],stage2_20[10],stage2_19[22],stage2_18[24]}
   );
   gpc615_5 gpc2175 (
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_19[31]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[6],stage2_20[11],stage2_19[23],stage2_18[25]}
   );
   gpc615_5 gpc2176 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46]},
      {stage1_19[32]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[7],stage2_20[12],stage2_19[24],stage2_18[26]}
   );
   gpc615_5 gpc2177 (
      {stage1_19[33], stage1_19[34], stage1_19[35], stage1_19[36], stage1_19[37]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[8],stage2_20[13],stage2_19[25]}
   );
   gpc615_5 gpc2178 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[19]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[9],stage2_20[14],stage2_19[26]}
   );
   gpc615_5 gpc2179 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[20]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[5],stage2_21[10],stage2_20[15],stage2_19[27]}
   );
   gpc606_5 gpc2180 (
      {stage1_20[21], stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[3],stage2_22[6],stage2_21[11],stage2_20[16]}
   );
   gpc606_5 gpc2181 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[4],stage2_22[7],stage2_21[12]}
   );
   gpc606_5 gpc2182 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[5],stage2_22[8],stage2_21[13]}
   );
   gpc606_5 gpc2183 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[6],stage2_22[9],stage2_21[14]}
   );
   gpc606_5 gpc2184 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[4],stage2_23[7],stage2_22[10],stage2_21[15]}
   );
   gpc606_5 gpc2185 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[5],stage2_23[8],stage2_22[11],stage2_21[16]}
   );
   gpc1163_5 gpc2186 (
      {stage1_22[6], stage1_22[7], stage1_22[8]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage1_24[0]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[5],stage2_24[6],stage2_23[9],stage2_22[12]}
   );
   gpc1163_5 gpc2187 (
      {stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage1_24[1]},
      {stage1_25[1]},
      {stage2_26[1],stage2_25[6],stage2_24[7],stage2_23[10],stage2_22[13]}
   );
   gpc1163_5 gpc2188 (
      {stage1_22[12], stage1_22[13], stage1_22[14]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[2]},
      {stage1_25[2]},
      {stage2_26[2],stage2_25[7],stage2_24[8],stage2_23[11],stage2_22[14]}
   );
   gpc1163_5 gpc2189 (
      {stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_24[3]},
      {stage1_25[3]},
      {stage2_26[3],stage2_25[8],stage2_24[9],stage2_23[12],stage2_22[15]}
   );
   gpc1163_5 gpc2190 (
      {stage1_22[18], stage1_22[19], stage1_22[20]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_24[4]},
      {stage1_25[4]},
      {stage2_26[4],stage2_25[9],stage2_24[10],stage2_23[13],stage2_22[16]}
   );
   gpc1163_5 gpc2191 (
      {stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_24[5]},
      {stage1_25[5]},
      {stage2_26[5],stage2_25[10],stage2_24[11],stage2_23[14],stage2_22[17]}
   );
   gpc1163_5 gpc2192 (
      {stage1_22[24], stage1_22[25], stage1_22[26]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_24[6]},
      {stage1_25[6]},
      {stage2_26[6],stage2_25[11],stage2_24[12],stage2_23[15],stage2_22[18]}
   );
   gpc615_5 gpc2193 (
      {stage1_22[27], stage1_22[28], stage1_22[29], stage1_22[30], stage1_22[31]},
      {stage1_23[72]},
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12]},
      {stage2_26[7],stage2_25[12],stage2_24[13],stage2_23[16],stage2_22[19]}
   );
   gpc615_5 gpc2194 (
      {stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35], stage1_22[36]},
      {stage1_23[73]},
      {stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage2_26[8],stage2_25[13],stage2_24[14],stage2_23[17],stage2_22[20]}
   );
   gpc615_5 gpc2195 (
      {stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_23[74]},
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24]},
      {stage2_26[9],stage2_25[14],stage2_24[15],stage2_23[18],stage2_22[21]}
   );
   gpc615_5 gpc2196 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46]},
      {stage1_23[75]},
      {stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30]},
      {stage2_26[10],stage2_25[15],stage2_24[16],stage2_23[19],stage2_22[22]}
   );
   gpc615_5 gpc2197 (
      {stage1_22[47], stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51]},
      {stage1_23[76]},
      {stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36]},
      {stage2_26[11],stage2_25[16],stage2_24[17],stage2_23[20],stage2_22[23]}
   );
   gpc615_5 gpc2198 (
      {stage1_22[52], stage1_22[53], stage1_22[54], stage1_22[55], stage1_22[56]},
      {stage1_23[77]},
      {stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42]},
      {stage2_26[12],stage2_25[17],stage2_24[18],stage2_23[21],stage2_22[24]}
   );
   gpc615_5 gpc2199 (
      {stage1_22[57], stage1_22[58], stage1_22[59], stage1_22[60], stage1_22[61]},
      {stage1_23[78]},
      {stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48]},
      {stage2_26[13],stage2_25[18],stage2_24[19],stage2_23[22],stage2_22[25]}
   );
   gpc606_5 gpc2200 (
      {stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[0],stage2_26[14],stage2_25[19],stage2_24[20],stage2_23[23]}
   );
   gpc606_5 gpc2201 (
      {stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[1],stage2_26[15],stage2_25[20],stage2_24[21],stage2_23[24]}
   );
   gpc606_5 gpc2202 (
      {stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[2],stage2_26[16],stage2_25[21],stage2_24[22],stage2_23[25]}
   );
   gpc606_5 gpc2203 (
      {stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[3],stage2_26[17],stage2_25[22],stage2_24[23],stage2_23[26]}
   );
   gpc606_5 gpc2204 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108]},
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage2_27[4],stage2_26[18],stage2_25[23],stage2_24[24],stage2_23[27]}
   );
   gpc606_5 gpc2205 (
      {stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114]},
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage2_27[5],stage2_26[19],stage2_25[24],stage2_24[25],stage2_23[28]}
   );
   gpc606_5 gpc2206 (
      {stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120]},
      {stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47], stage1_25[48]},
      {stage2_27[6],stage2_26[20],stage2_25[25],stage2_24[26],stage2_23[29]}
   );
   gpc606_5 gpc2207 (
      {stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126]},
      {stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53], stage1_25[54]},
      {stage2_27[7],stage2_26[21],stage2_25[26],stage2_24[27],stage2_23[30]}
   );
   gpc615_5 gpc2208 (
      {stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_25[55]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[22],stage2_25[27],stage2_24[28]}
   );
   gpc615_5 gpc2209 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58]},
      {stage1_25[56]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[23],stage2_25[28],stage2_24[29]}
   );
   gpc615_5 gpc2210 (
      {stage1_24[59], stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63]},
      {stage1_25[57]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[24],stage2_25[29],stage2_24[30]}
   );
   gpc615_5 gpc2211 (
      {stage1_24[64], stage1_24[65], stage1_24[66], stage1_24[67], stage1_24[68]},
      {stage1_25[58]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[25],stage2_25[30],stage2_24[31]}
   );
   gpc606_5 gpc2212 (
      {stage1_25[59], stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[4],stage2_27[12],stage2_26[26],stage2_25[31]}
   );
   gpc606_5 gpc2213 (
      {stage1_25[65], stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[5],stage2_27[13],stage2_26[27],stage2_25[32]}
   );
   gpc606_5 gpc2214 (
      {stage1_25[71], stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[6],stage2_27[14],stage2_26[28],stage2_25[33]}
   );
   gpc606_5 gpc2215 (
      {stage1_25[77], stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[7],stage2_27[15],stage2_26[29],stage2_25[34]}
   );
   gpc2116_5 gpc2216 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_27[24]},
      {stage1_28[0]},
      {stage1_29[0], stage1_29[1]},
      {stage2_30[0],stage2_29[4],stage2_28[8],stage2_27[16],stage2_26[30]}
   );
   gpc2116_5 gpc2217 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[25]},
      {stage1_28[1]},
      {stage1_29[2], stage1_29[3]},
      {stage2_30[1],stage2_29[5],stage2_28[9],stage2_27[17],stage2_26[31]}
   );
   gpc2116_5 gpc2218 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_27[26]},
      {stage1_28[2]},
      {stage1_29[4], stage1_29[5]},
      {stage2_30[2],stage2_29[6],stage2_28[10],stage2_27[18],stage2_26[32]}
   );
   gpc2116_5 gpc2219 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_27[27]},
      {stage1_28[3]},
      {stage1_29[6], stage1_29[7]},
      {stage2_30[3],stage2_29[7],stage2_28[11],stage2_27[19],stage2_26[33]}
   );
   gpc2116_5 gpc2220 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_27[28]},
      {stage1_28[4]},
      {stage1_29[8], stage1_29[9]},
      {stage2_30[4],stage2_29[8],stage2_28[12],stage2_27[20],stage2_26[34]}
   );
   gpc615_5 gpc2221 (
      {stage1_27[29], stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33]},
      {stage1_28[5]},
      {stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15]},
      {stage2_31[0],stage2_30[5],stage2_29[9],stage2_28[13],stage2_27[21]}
   );
   gpc615_5 gpc2222 (
      {stage1_27[34], stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38]},
      {stage1_28[6]},
      {stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21]},
      {stage2_31[1],stage2_30[6],stage2_29[10],stage2_28[14],stage2_27[22]}
   );
   gpc615_5 gpc2223 (
      {stage1_27[39], stage1_27[40], stage1_27[41], stage1_27[42], stage1_27[43]},
      {stage1_28[7]},
      {stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27]},
      {stage2_31[2],stage2_30[7],stage2_29[11],stage2_28[15],stage2_27[23]}
   );
   gpc615_5 gpc2224 (
      {stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47], stage1_27[48]},
      {stage1_28[8]},
      {stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33]},
      {stage2_31[3],stage2_30[8],stage2_29[12],stage2_28[16],stage2_27[24]}
   );
   gpc606_5 gpc2225 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[4],stage2_30[9],stage2_29[13],stage2_28[17]}
   );
   gpc606_5 gpc2226 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[5],stage2_30[10],stage2_29[14],stage2_28[18]}
   );
   gpc606_5 gpc2227 (
      {stage1_28[21], stage1_28[22], stage1_28[23], stage1_28[24], stage1_28[25], stage1_28[26]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[6],stage2_30[11],stage2_29[15],stage2_28[19]}
   );
   gpc606_5 gpc2228 (
      {stage1_28[27], stage1_28[28], stage1_28[29], stage1_28[30], stage1_28[31], stage1_28[32]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[7],stage2_30[12],stage2_29[16],stage2_28[20]}
   );
   gpc606_5 gpc2229 (
      {stage1_28[33], stage1_28[34], stage1_28[35], stage1_28[36], stage1_28[37], stage1_28[38]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[8],stage2_30[13],stage2_29[17],stage2_28[21]}
   );
   gpc606_5 gpc2230 (
      {stage1_28[39], stage1_28[40], stage1_28[41], stage1_28[42], stage1_28[43], stage1_28[44]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[9],stage2_30[14],stage2_29[18],stage2_28[22]}
   );
   gpc606_5 gpc2231 (
      {stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49], stage1_28[50]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[10],stage2_30[15],stage2_29[19],stage2_28[23]}
   );
   gpc606_5 gpc2232 (
      {stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55], stage1_28[56]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[11],stage2_30[16],stage2_29[20],stage2_28[24]}
   );
   gpc606_5 gpc2233 (
      {stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61], stage1_28[62]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[12],stage2_30[17],stage2_29[21],stage2_28[25]}
   );
   gpc606_5 gpc2234 (
      {stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66], stage1_28[67], stage1_28[68]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[13],stage2_30[18],stage2_29[22],stage2_28[26]}
   );
   gpc606_5 gpc2235 (
      {stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[10],stage2_31[14],stage2_30[19],stage2_29[23]}
   );
   gpc606_5 gpc2236 (
      {stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[11],stage2_31[15],stage2_30[20],stage2_29[24]}
   );
   gpc606_5 gpc2237 (
      {stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[12],stage2_31[16],stage2_30[21],stage2_29[25]}
   );
   gpc606_5 gpc2238 (
      {stage1_29[52], stage1_29[53], stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[13],stage2_31[17],stage2_30[22],stage2_29[26]}
   );
   gpc606_5 gpc2239 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[4],stage2_32[14],stage2_31[18],stage2_30[23]}
   );
   gpc606_5 gpc2240 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[5],stage2_32[15],stage2_31[19],stage2_30[24]}
   );
   gpc606_5 gpc2241 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[6],stage2_32[16],stage2_31[20],stage2_30[25]}
   );
   gpc606_5 gpc2242 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[7],stage2_32[17],stage2_31[21],stage2_30[26]}
   );
   gpc615_5 gpc2243 (
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28]},
      {stage1_32[24]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[4],stage2_33[8],stage2_32[18],stage2_31[22]}
   );
   gpc615_5 gpc2244 (
      {stage1_31[29], stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33]},
      {stage1_32[25]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[5],stage2_33[9],stage2_32[19],stage2_31[23]}
   );
   gpc615_5 gpc2245 (
      {stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_32[26]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[6],stage2_33[10],stage2_32[20],stage2_31[24]}
   );
   gpc615_5 gpc2246 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43]},
      {stage1_32[27]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[7],stage2_33[11],stage2_32[21],stage2_31[25]}
   );
   gpc615_5 gpc2247 (
      {stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48]},
      {stage1_32[28]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[8],stage2_33[12],stage2_32[22],stage2_31[26]}
   );
   gpc615_5 gpc2248 (
      {stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage1_32[29]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[9],stage2_33[13],stage2_32[23],stage2_31[27]}
   );
   gpc615_5 gpc2249 (
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58]},
      {stage1_32[30]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[10],stage2_33[14],stage2_32[24],stage2_31[28]}
   );
   gpc615_5 gpc2250 (
      {stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63]},
      {stage1_32[31]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[11],stage2_33[15],stage2_32[25],stage2_31[29]}
   );
   gpc615_5 gpc2251 (
      {stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_32[32]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[12],stage2_33[16],stage2_32[26],stage2_31[30]}
   );
   gpc615_5 gpc2252 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73]},
      {stage1_32[33]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[13],stage2_33[17],stage2_32[27],stage2_31[31]}
   );
   gpc615_5 gpc2253 (
      {stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78]},
      {stage1_32[34]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[14],stage2_33[18],stage2_32[28],stage2_31[32]}
   );
   gpc615_5 gpc2254 (
      {stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_32[35]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[15],stage2_33[19],stage2_32[29],stage2_31[33]}
   );
   gpc615_5 gpc2255 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88]},
      {stage1_32[36]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[16],stage2_33[20],stage2_32[30],stage2_31[34]}
   );
   gpc615_5 gpc2256 (
      {stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93]},
      {stage1_32[37]},
      {stage1_33[78], stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83]},
      {stage2_35[13],stage2_34[17],stage2_33[21],stage2_32[31],stage2_31[35]}
   );
   gpc606_5 gpc2257 (
      {stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[14],stage2_34[18],stage2_33[22],stage2_32[32]}
   );
   gpc606_5 gpc2258 (
      {stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[15],stage2_34[19],stage2_33[23],stage2_32[33]}
   );
   gpc606_5 gpc2259 (
      {stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[16],stage2_34[20],stage2_33[24],stage2_32[34]}
   );
   gpc606_5 gpc2260 (
      {stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[17],stage2_34[21],stage2_33[25],stage2_32[35]}
   );
   gpc606_5 gpc2261 (
      {stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[18],stage2_34[22],stage2_33[26],stage2_32[36]}
   );
   gpc606_5 gpc2262 (
      {stage1_33[84], stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[5],stage2_35[19],stage2_34[23],stage2_33[27]}
   );
   gpc606_5 gpc2263 (
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[1],stage2_36[6],stage2_35[20],stage2_34[24]}
   );
   gpc606_5 gpc2264 (
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[2],stage2_36[7],stage2_35[21],stage2_34[25]}
   );
   gpc606_5 gpc2265 (
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[3],stage2_36[8],stage2_35[22],stage2_34[26]}
   );
   gpc615_5 gpc2266 (
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[4],stage2_36[9],stage2_35[23]}
   );
   gpc615_5 gpc2267 (
      {stage1_35[11], stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15]},
      {stage1_36[19]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[4],stage2_37[5],stage2_36[10],stage2_35[24]}
   );
   gpc615_5 gpc2268 (
      {stage1_35[16], stage1_35[17], stage1_35[18], stage1_35[19], stage1_35[20]},
      {stage1_36[20]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[5],stage2_37[6],stage2_36[11],stage2_35[25]}
   );
   gpc615_5 gpc2269 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[21]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[6],stage2_37[7],stage2_36[12],stage2_35[26]}
   );
   gpc615_5 gpc2270 (
      {stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage1_36[22]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[7],stage2_37[8],stage2_36[13],stage2_35[27]}
   );
   gpc615_5 gpc2271 (
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage1_36[23]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[8],stage2_37[9],stage2_36[14],stage2_35[28]}
   );
   gpc615_5 gpc2272 (
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40]},
      {stage1_36[24]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[9],stage2_37[10],stage2_36[15],stage2_35[29]}
   );
   gpc615_5 gpc2273 (
      {stage1_35[41], stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45]},
      {stage1_36[25]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[10],stage2_37[11],stage2_36[16],stage2_35[30]}
   );
   gpc1343_5 gpc2274 (
      {stage1_36[26], stage1_36[27], stage1_36[28]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51]},
      {stage1_38[0], stage1_38[1], stage1_38[2]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[8],stage2_38[11],stage2_37[12],stage2_36[17]}
   );
   gpc606_5 gpc2275 (
      {stage1_36[29], stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34]},
      {stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8]},
      {stage2_40[1],stage2_39[9],stage2_38[12],stage2_37[13],stage2_36[18]}
   );
   gpc606_5 gpc2276 (
      {stage1_36[35], stage1_36[36], stage1_36[37], stage1_36[38], stage1_36[39], stage1_36[40]},
      {stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14]},
      {stage2_40[2],stage2_39[10],stage2_38[13],stage2_37[14],stage2_36[19]}
   );
   gpc606_5 gpc2277 (
      {stage1_36[41], stage1_36[42], stage1_36[43], stage1_36[44], stage1_36[45], stage1_36[46]},
      {stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage2_40[3],stage2_39[11],stage2_38[14],stage2_37[15],stage2_36[20]}
   );
   gpc615_5 gpc2278 (
      {stage1_36[47], stage1_36[48], stage1_36[49], stage1_36[50], stage1_36[51]},
      {stage1_37[52]},
      {stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26]},
      {stage2_40[4],stage2_39[12],stage2_38[15],stage2_37[16],stage2_36[21]}
   );
   gpc615_5 gpc2279 (
      {stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55], stage1_36[56]},
      {stage1_37[53]},
      {stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32]},
      {stage2_40[5],stage2_39[13],stage2_38[16],stage2_37[17],stage2_36[22]}
   );
   gpc615_5 gpc2280 (
      {stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage1_37[54]},
      {stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38]},
      {stage2_40[6],stage2_39[14],stage2_38[17],stage2_37[18],stage2_36[23]}
   );
   gpc615_5 gpc2281 (
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66]},
      {stage1_37[55]},
      {stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44]},
      {stage2_40[7],stage2_39[15],stage2_38[18],stage2_37[19],stage2_36[24]}
   );
   gpc615_5 gpc2282 (
      {stage1_36[67], stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71]},
      {stage1_37[56]},
      {stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50]},
      {stage2_40[8],stage2_39[16],stage2_38[19],stage2_37[20],stage2_36[25]}
   );
   gpc606_5 gpc2283 (
      {stage1_37[57], stage1_37[58], stage1_37[59], stage1_37[60], stage1_37[61], stage1_37[62]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[9],stage2_39[17],stage2_38[20],stage2_37[21]}
   );
   gpc606_5 gpc2284 (
      {stage1_37[63], stage1_37[64], stage1_37[65], stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[10],stage2_39[18],stage2_38[21],stage2_37[22]}
   );
   gpc606_5 gpc2285 (
      {stage1_37[69], stage1_37[70], stage1_37[71], stage1_37[72], stage1_37[73], stage1_37[74]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[11],stage2_39[19],stage2_38[22],stage2_37[23]}
   );
   gpc606_5 gpc2286 (
      {stage1_37[75], stage1_37[76], stage1_37[77], stage1_37[78], stage1_37[79], stage1_37[80]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[12],stage2_39[20],stage2_38[23],stage2_37[24]}
   );
   gpc606_5 gpc2287 (
      {stage1_37[81], stage1_37[82], stage1_37[83], stage1_37[84], stage1_37[85], stage1_37[86]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[13],stage2_39[21],stage2_38[24],stage2_37[25]}
   );
   gpc606_5 gpc2288 (
      {stage1_37[87], stage1_37[88], stage1_37[89], stage1_37[90], stage1_37[91], stage1_37[92]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[14],stage2_39[22],stage2_38[25],stage2_37[26]}
   );
   gpc606_5 gpc2289 (
      {stage1_37[93], stage1_37[94], stage1_37[95], stage1_37[96], stage1_37[97], stage1_37[98]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[15],stage2_39[23],stage2_38[26],stage2_37[27]}
   );
   gpc606_5 gpc2290 (
      {stage1_37[99], stage1_37[100], stage1_37[101], stage1_37[102], stage1_37[103], stage1_37[104]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[16],stage2_39[24],stage2_38[27],stage2_37[28]}
   );
   gpc606_5 gpc2291 (
      {stage1_37[105], stage1_37[106], stage1_37[107], stage1_37[108], stage1_37[109], stage1_37[110]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[17],stage2_39[25],stage2_38[28],stage2_37[29]}
   );
   gpc606_5 gpc2292 (
      {stage1_37[111], stage1_37[112], stage1_37[113], stage1_37[114], stage1_37[115], stage1_37[116]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[18],stage2_39[26],stage2_38[29],stage2_37[30]}
   );
   gpc615_5 gpc2293 (
      {stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55]},
      {stage1_39[61]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[10],stage2_40[19],stage2_39[27],stage2_38[30]}
   );
   gpc615_5 gpc2294 (
      {stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage1_39[62]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[11],stage2_40[20],stage2_39[28],stage2_38[31]}
   );
   gpc615_5 gpc2295 (
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65]},
      {stage1_39[63]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[12],stage2_40[21],stage2_39[29],stage2_38[32]}
   );
   gpc606_5 gpc2296 (
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[13],stage2_40[22]}
   );
   gpc606_5 gpc2297 (
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[14],stage2_40[23]}
   );
   gpc606_5 gpc2298 (
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[15],stage2_40[24]}
   );
   gpc606_5 gpc2299 (
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[16],stage2_40[25]}
   );
   gpc606_5 gpc2300 (
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[17],stage2_40[26]}
   );
   gpc606_5 gpc2301 (
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[8],stage2_41[18],stage2_40[27]}
   );
   gpc606_5 gpc2302 (
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[9],stage2_41[19],stage2_40[28]}
   );
   gpc606_5 gpc2303 (
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[10],stage2_41[20],stage2_40[29]}
   );
   gpc606_5 gpc2304 (
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[11],stage2_41[21],stage2_40[30]}
   );
   gpc606_5 gpc2305 (
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[9],stage2_43[9],stage2_42[12],stage2_41[22]}
   );
   gpc606_5 gpc2306 (
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[10],stage2_43[10],stage2_42[13],stage2_41[23]}
   );
   gpc606_5 gpc2307 (
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[11],stage2_43[11],stage2_42[14],stage2_41[24]}
   );
   gpc606_5 gpc2308 (
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[12],stage2_43[12],stage2_42[15],stage2_41[25]}
   );
   gpc606_5 gpc2309 (
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[13],stage2_43[13],stage2_42[16],stage2_41[26]}
   );
   gpc606_5 gpc2310 (
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[14],stage2_43[14],stage2_42[17],stage2_41[27]}
   );
   gpc606_5 gpc2311 (
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[15],stage2_43[15],stage2_42[18],stage2_41[28]}
   );
   gpc606_5 gpc2312 (
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[16],stage2_43[16],stage2_42[19],stage2_41[29]}
   );
   gpc606_5 gpc2313 (
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[8],stage2_44[17],stage2_43[17]}
   );
   gpc606_5 gpc2314 (
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[9],stage2_44[18],stage2_43[18]}
   );
   gpc606_5 gpc2315 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[10],stage2_44[19],stage2_43[19]}
   );
   gpc606_5 gpc2316 (
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[3],stage2_45[11],stage2_44[20],stage2_43[20]}
   );
   gpc606_5 gpc2317 (
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[4],stage2_45[12],stage2_44[21],stage2_43[21]}
   );
   gpc606_5 gpc2318 (
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[5],stage2_45[13],stage2_44[22],stage2_43[22]}
   );
   gpc606_5 gpc2319 (
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[6],stage2_45[14],stage2_44[23],stage2_43[23]}
   );
   gpc606_5 gpc2320 (
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[7],stage2_45[15],stage2_44[24],stage2_43[24]}
   );
   gpc606_5 gpc2321 (
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[8],stage2_45[16],stage2_44[25],stage2_43[25]}
   );
   gpc606_5 gpc2322 (
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[9],stage2_45[17],stage2_44[26],stage2_43[26]}
   );
   gpc606_5 gpc2323 (
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[10],stage2_45[18],stage2_44[27],stage2_43[27]}
   );
   gpc615_5 gpc2324 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[66]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[11],stage2_46[11],stage2_45[19],stage2_44[28]}
   );
   gpc615_5 gpc2325 (
      {stage1_44[5], stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9]},
      {stage1_45[67]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[12],stage2_46[12],stage2_45[20],stage2_44[29]}
   );
   gpc606_5 gpc2326 (
      {stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[2],stage2_47[13],stage2_46[13],stage2_45[21]}
   );
   gpc606_5 gpc2327 (
      {stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[3],stage2_47[14],stage2_46[14],stage2_45[22]}
   );
   gpc606_5 gpc2328 (
      {stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[4],stage2_47[15],stage2_46[15],stage2_45[23]}
   );
   gpc606_5 gpc2329 (
      {stage1_45[86], stage1_45[87], stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[5],stage2_47[16],stage2_46[16],stage2_45[24]}
   );
   gpc615_5 gpc2330 (
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16]},
      {stage1_47[24]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[4],stage2_48[6],stage2_47[17],stage2_46[17]}
   );
   gpc615_5 gpc2331 (
      {stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage1_47[25]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[5],stage2_48[7],stage2_47[18],stage2_46[18]}
   );
   gpc615_5 gpc2332 (
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26]},
      {stage1_47[26]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[6],stage2_48[8],stage2_47[19],stage2_46[19]}
   );
   gpc615_5 gpc2333 (
      {stage1_46[27], stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31]},
      {stage1_47[27]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[7],stage2_48[9],stage2_47[20],stage2_46[20]}
   );
   gpc615_5 gpc2334 (
      {stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35], stage1_46[36]},
      {stage1_47[28]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[8],stage2_48[10],stage2_47[21],stage2_46[21]}
   );
   gpc615_5 gpc2335 (
      {stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage1_47[29]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[9],stage2_48[11],stage2_47[22],stage2_46[22]}
   );
   gpc615_5 gpc2336 (
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46]},
      {stage1_47[30]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[10],stage2_48[12],stage2_47[23],stage2_46[23]}
   );
   gpc615_5 gpc2337 (
      {stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage1_47[31]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[11],stage2_48[13],stage2_47[24],stage2_46[24]}
   );
   gpc615_5 gpc2338 (
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56]},
      {stage1_47[32]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[12],stage2_48[14],stage2_47[25],stage2_46[25]}
   );
   gpc606_5 gpc2339 (
      {stage1_47[33], stage1_47[34], stage1_47[35], stage1_47[36], stage1_47[37], stage1_47[38]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[9],stage2_49[13],stage2_48[15],stage2_47[26]}
   );
   gpc606_5 gpc2340 (
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[1],stage2_50[10],stage2_49[14],stage2_48[16]}
   );
   gpc606_5 gpc2341 (
      {stage1_48[60], stage1_48[61], stage1_48[62], stage1_48[63], stage1_48[64], stage1_48[65]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[2],stage2_50[11],stage2_49[15],stage2_48[17]}
   );
   gpc606_5 gpc2342 (
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[2],stage2_51[3],stage2_50[12],stage2_49[16]}
   );
   gpc606_5 gpc2343 (
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[3],stage2_51[4],stage2_50[13],stage2_49[17]}
   );
   gpc606_5 gpc2344 (
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[4],stage2_51[5],stage2_50[14],stage2_49[18]}
   );
   gpc606_5 gpc2345 (
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[5],stage2_51[6],stage2_50[15],stage2_49[19]}
   );
   gpc606_5 gpc2346 (
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[6],stage2_51[7],stage2_50[16],stage2_49[20]}
   );
   gpc606_5 gpc2347 (
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[7],stage2_51[8],stage2_50[17],stage2_49[21]}
   );
   gpc606_5 gpc2348 (
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[8],stage2_51[9],stage2_50[18],stage2_49[22]}
   );
   gpc606_5 gpc2349 (
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[9],stage2_51[10],stage2_50[19],stage2_49[23]}
   );
   gpc606_5 gpc2350 (
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[10],stage2_51[11],stage2_50[20],stage2_49[24]}
   );
   gpc606_5 gpc2351 (
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[11],stage2_51[12],stage2_50[21],stage2_49[25]}
   );
   gpc606_5 gpc2352 (
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage2_53[10],stage2_52[12],stage2_51[13],stage2_50[22],stage2_49[26]}
   );
   gpc606_5 gpc2353 (
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage1_51[66], stage1_51[67], stage1_51[68], stage1_51[69], stage1_51[70], stage1_51[71]},
      {stage2_53[11],stage2_52[13],stage2_51[14],stage2_50[23],stage2_49[27]}
   );
   gpc117_4 gpc2354 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18]},
      {stage1_51[72]},
      {stage1_52[0]},
      {stage2_53[12],stage2_52[14],stage2_51[15],stage2_50[24]}
   );
   gpc606_5 gpc2355 (
      {stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5], stage1_52[6]},
      {stage2_54[0],stage2_53[13],stage2_52[15],stage2_51[16],stage2_50[25]}
   );
   gpc606_5 gpc2356 (
      {stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30]},
      {stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11], stage1_52[12]},
      {stage2_54[1],stage2_53[14],stage2_52[16],stage2_51[17],stage2_50[26]}
   );
   gpc606_5 gpc2357 (
      {stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17], stage1_52[18]},
      {stage2_54[2],stage2_53[15],stage2_52[17],stage2_51[18],stage2_50[27]}
   );
   gpc615_5 gpc2358 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[73]},
      {stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23], stage1_52[24]},
      {stage2_54[3],stage2_53[16],stage2_52[18],stage2_51[19],stage2_50[28]}
   );
   gpc615_5 gpc2359 (
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46]},
      {stage1_51[74]},
      {stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29], stage1_52[30]},
      {stage2_54[4],stage2_53[17],stage2_52[19],stage2_51[20],stage2_50[29]}
   );
   gpc606_5 gpc2360 (
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_53[0], stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage2_55[0],stage2_54[5],stage2_53[18],stage2_52[20],stage2_51[21]}
   );
   gpc606_5 gpc2361 (
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage2_55[1],stage2_54[6],stage2_53[19],stage2_52[21],stage2_51[22]}
   );
   gpc606_5 gpc2362 (
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16], stage1_53[17]},
      {stage2_55[2],stage2_54[7],stage2_53[20],stage2_52[22],stage2_51[23]}
   );
   gpc606_5 gpc2363 (
      {stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[3],stage2_54[8],stage2_53[21],stage2_52[23]}
   );
   gpc606_5 gpc2364 (
      {stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[4],stage2_54[9],stage2_53[22],stage2_52[24]}
   );
   gpc606_5 gpc2365 (
      {stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47], stage1_52[48]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[5],stage2_54[10],stage2_53[23],stage2_52[25]}
   );
   gpc606_5 gpc2366 (
      {stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53], stage1_52[54]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[6],stage2_54[11],stage2_53[24],stage2_52[26]}
   );
   gpc606_5 gpc2367 (
      {stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59], stage1_52[60]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[7],stage2_54[12],stage2_53[25],stage2_52[27]}
   );
   gpc606_5 gpc2368 (
      {stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65], stage1_52[66]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[8],stage2_54[13],stage2_53[26],stage2_52[28]}
   );
   gpc606_5 gpc2369 (
      {stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71], stage1_52[72]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[9],stage2_54[14],stage2_53[27],stage2_52[29]}
   );
   gpc606_5 gpc2370 (
      {stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[7],stage2_55[10],stage2_54[15],stage2_53[28]}
   );
   gpc606_5 gpc2371 (
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[8],stage2_55[11],stage2_54[16],stage2_53[29]}
   );
   gpc606_5 gpc2372 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[9],stage2_55[12],stage2_54[17],stage2_53[30]}
   );
   gpc606_5 gpc2373 (
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[10],stage2_55[13],stage2_54[18],stage2_53[31]}
   );
   gpc606_5 gpc2374 (
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[11],stage2_55[14],stage2_54[19],stage2_53[32]}
   );
   gpc615_5 gpc2375 (
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46]},
      {stage1_55[30]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[5],stage2_56[12],stage2_55[15],stage2_54[20]}
   );
   gpc615_5 gpc2376 (
      {stage1_54[47], stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51]},
      {stage1_55[31]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[6],stage2_56[13],stage2_55[16],stage2_54[21]}
   );
   gpc606_5 gpc2377 (
      {stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[7],stage2_56[14],stage2_55[17]}
   );
   gpc615_5 gpc2378 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[8],stage2_56[15],stage2_55[18]}
   );
   gpc615_5 gpc2379 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[13]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[9],stage2_56[16],stage2_55[19]}
   );
   gpc615_5 gpc2380 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[14]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[10],stage2_56[17],stage2_55[20]}
   );
   gpc615_5 gpc2381 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[15]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[11],stage2_56[18],stage2_55[21]}
   );
   gpc615_5 gpc2382 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[16]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[5],stage2_58[7],stage2_57[12],stage2_56[19],stage2_55[22]}
   );
   gpc615_5 gpc2383 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[17]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[6],stage2_58[8],stage2_57[13],stage2_56[20],stage2_55[23]}
   );
   gpc615_5 gpc2384 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[18]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[7],stage2_58[9],stage2_57[14],stage2_56[21],stage2_55[24]}
   );
   gpc615_5 gpc2385 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[19]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[8],stage2_58[10],stage2_57[15],stage2_56[22],stage2_55[25]}
   );
   gpc615_5 gpc2386 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[20]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[9],stage2_58[11],stage2_57[16],stage2_56[23],stage2_55[26]}
   );
   gpc615_5 gpc2387 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[21]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[10],stage2_58[12],stage2_57[17],stage2_56[24],stage2_55[27]}
   );
   gpc606_5 gpc2388 (
      {stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[11],stage2_58[13],stage2_57[18],stage2_56[25]}
   );
   gpc606_5 gpc2389 (
      {stage1_56[28], stage1_56[29], stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[12],stage2_58[14],stage2_57[19],stage2_56[26]}
   );
   gpc606_5 gpc2390 (
      {stage1_56[34], stage1_56[35], stage1_56[36], stage1_56[37], stage1_56[38], stage1_56[39]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[13],stage2_58[15],stage2_57[20],stage2_56[27]}
   );
   gpc606_5 gpc2391 (
      {stage1_56[40], stage1_56[41], stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45]},
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage2_60[3],stage2_59[14],stage2_58[16],stage2_57[21],stage2_56[28]}
   );
   gpc606_5 gpc2392 (
      {stage1_56[46], stage1_56[47], stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51]},
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage2_60[4],stage2_59[15],stage2_58[17],stage2_57[22],stage2_56[29]}
   );
   gpc606_5 gpc2393 (
      {stage1_56[52], stage1_56[53], stage1_56[54], stage1_56[55], stage1_56[56], stage1_56[57]},
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage2_60[5],stage2_59[16],stage2_58[18],stage2_57[23],stage2_56[30]}
   );
   gpc606_5 gpc2394 (
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[0],stage2_60[6],stage2_59[17],stage2_58[19]}
   );
   gpc606_5 gpc2395 (
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[1],stage2_60[7],stage2_59[18],stage2_58[20]}
   );
   gpc606_5 gpc2396 (
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[2],stage2_60[8],stage2_59[19],stage2_58[21]}
   );
   gpc606_5 gpc2397 (
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[3],stage2_60[9],stage2_59[20],stage2_58[22]}
   );
   gpc615_5 gpc2398 (
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64]},
      {stage1_59[0]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[4],stage2_60[10],stage2_59[21],stage2_58[23]}
   );
   gpc606_5 gpc2399 (
      {stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5], stage1_59[6]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[5],stage2_60[11],stage2_59[22]}
   );
   gpc606_5 gpc2400 (
      {stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11], stage1_59[12]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[6],stage2_60[12],stage2_59[23]}
   );
   gpc606_5 gpc2401 (
      {stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17], stage1_59[18]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[7],stage2_60[13],stage2_59[24]}
   );
   gpc606_5 gpc2402 (
      {stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[8],stage2_60[14],stage2_59[25]}
   );
   gpc606_5 gpc2403 (
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[4],stage2_62[9],stage2_61[9],stage2_60[15]}
   );
   gpc606_5 gpc2404 (
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[5],stage2_62[10],stage2_61[10],stage2_60[16]}
   );
   gpc606_5 gpc2405 (
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[6],stage2_62[11],stage2_61[11],stage2_60[17]}
   );
   gpc606_5 gpc2406 (
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage2_64[3],stage2_63[7],stage2_62[12],stage2_61[12],stage2_60[18]}
   );
   gpc606_5 gpc2407 (
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage2_64[4],stage2_63[8],stage2_62[13],stage2_61[13],stage2_60[19]}
   );
   gpc606_5 gpc2408 (
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage2_64[5],stage2_63[9],stage2_62[14],stage2_61[14],stage2_60[20]}
   );
   gpc606_5 gpc2409 (
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[6],stage2_63[10],stage2_62[15],stage2_61[15]}
   );
   gpc606_5 gpc2410 (
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[7],stage2_63[11],stage2_62[16],stage2_61[16]}
   );
   gpc606_5 gpc2411 (
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[8],stage2_63[12],stage2_62[17],stage2_61[17]}
   );
   gpc2135_5 gpc2412 (
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40]},
      {stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_64[0]},
      {stage1_65[0], stage1_65[1]},
      {stage2_66[0],stage2_65[3],stage2_64[9],stage2_63[13],stage2_62[18]}
   );
   gpc2135_5 gpc2413 (
      {stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[2], stage1_65[3]},
      {stage2_66[1],stage2_65[4],stage2_64[10],stage2_63[14],stage2_62[19]}
   );
   gpc2135_5 gpc2414 (
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50]},
      {stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_64[2]},
      {stage1_65[4], stage1_65[5]},
      {stage2_66[2],stage2_65[5],stage2_64[11],stage2_63[15],stage2_62[20]}
   );
   gpc2135_5 gpc2415 (
      {stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage1_64[3]},
      {stage1_65[6], stage1_65[7]},
      {stage2_66[3],stage2_65[6],stage2_64[12],stage2_63[16],stage2_62[21]}
   );
   gpc2135_5 gpc2416 (
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60]},
      {stage1_63[30], stage1_63[31], stage1_63[32]},
      {stage1_64[4]},
      {stage1_65[8], stage1_65[9]},
      {stage2_66[4],stage2_65[7],stage2_64[13],stage2_63[17],stage2_62[22]}
   );
   gpc2135_5 gpc2417 (
      {stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_64[5]},
      {stage1_65[10], stage1_65[11]},
      {stage2_66[5],stage2_65[8],stage2_64[14],stage2_63[18],stage2_62[23]}
   );
   gpc606_5 gpc2418 (
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71]},
      {stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11]},
      {stage2_66[6],stage2_65[9],stage2_64[15],stage2_63[19],stage2_62[24]}
   );
   gpc606_5 gpc2419 (
      {stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77]},
      {stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17]},
      {stage2_66[7],stage2_65[10],stage2_64[16],stage2_63[20],stage2_62[25]}
   );
   gpc606_5 gpc2420 (
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[0],stage2_66[8],stage2_65[11],stage2_64[17],stage2_63[21]}
   );
   gpc606_5 gpc2421 (
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage1_65[18], stage1_65[19], stage1_65[20], stage1_65[21], stage1_65[22], stage1_65[23]},
      {stage2_67[1],stage2_66[9],stage2_65[12],stage2_64[18],stage2_63[22]}
   );
   gpc1_1 gpc2422 (
      {stage1_0[31]},
      {stage2_0[7]}
   );
   gpc1_1 gpc2423 (
      {stage1_0[32]},
      {stage2_0[8]}
   );
   gpc1_1 gpc2424 (
      {stage1_0[33]},
      {stage2_0[9]}
   );
   gpc1_1 gpc2425 (
      {stage1_1[38]},
      {stage2_1[10]}
   );
   gpc1_1 gpc2426 (
      {stage1_1[39]},
      {stage2_1[11]}
   );
   gpc1_1 gpc2427 (
      {stage1_1[40]},
      {stage2_1[12]}
   );
   gpc1_1 gpc2428 (
      {stage1_1[41]},
      {stage2_1[13]}
   );
   gpc1_1 gpc2429 (
      {stage1_1[42]},
      {stage2_1[14]}
   );
   gpc1_1 gpc2430 (
      {stage1_1[43]},
      {stage2_1[15]}
   );
   gpc1_1 gpc2431 (
      {stage1_1[44]},
      {stage2_1[16]}
   );
   gpc1_1 gpc2432 (
      {stage1_1[45]},
      {stage2_1[17]}
   );
   gpc1_1 gpc2433 (
      {stage1_1[46]},
      {stage2_1[18]}
   );
   gpc1_1 gpc2434 (
      {stage1_2[27]},
      {stage2_2[10]}
   );
   gpc1_1 gpc2435 (
      {stage1_2[28]},
      {stage2_2[11]}
   );
   gpc1_1 gpc2436 (
      {stage1_2[29]},
      {stage2_2[12]}
   );
   gpc1_1 gpc2437 (
      {stage1_2[30]},
      {stage2_2[13]}
   );
   gpc1_1 gpc2438 (
      {stage1_2[31]},
      {stage2_2[14]}
   );
   gpc1_1 gpc2439 (
      {stage1_2[32]},
      {stage2_2[15]}
   );
   gpc1_1 gpc2440 (
      {stage1_2[33]},
      {stage2_2[16]}
   );
   gpc1_1 gpc2441 (
      {stage1_2[34]},
      {stage2_2[17]}
   );
   gpc1_1 gpc2442 (
      {stage1_2[35]},
      {stage2_2[18]}
   );
   gpc1_1 gpc2443 (
      {stage1_2[36]},
      {stage2_2[19]}
   );
   gpc1_1 gpc2444 (
      {stage1_2[37]},
      {stage2_2[20]}
   );
   gpc1_1 gpc2445 (
      {stage1_2[38]},
      {stage2_2[21]}
   );
   gpc1_1 gpc2446 (
      {stage1_2[39]},
      {stage2_2[22]}
   );
   gpc1_1 gpc2447 (
      {stage1_2[40]},
      {stage2_2[23]}
   );
   gpc1_1 gpc2448 (
      {stage1_2[41]},
      {stage2_2[24]}
   );
   gpc1_1 gpc2449 (
      {stage1_2[42]},
      {stage2_2[25]}
   );
   gpc1_1 gpc2450 (
      {stage1_2[43]},
      {stage2_2[26]}
   );
   gpc1_1 gpc2451 (
      {stage1_2[44]},
      {stage2_2[27]}
   );
   gpc1_1 gpc2452 (
      {stage1_2[45]},
      {stage2_2[28]}
   );
   gpc1_1 gpc2453 (
      {stage1_2[46]},
      {stage2_2[29]}
   );
   gpc1_1 gpc2454 (
      {stage1_2[47]},
      {stage2_2[30]}
   );
   gpc1_1 gpc2455 (
      {stage1_2[48]},
      {stage2_2[31]}
   );
   gpc1_1 gpc2456 (
      {stage1_2[49]},
      {stage2_2[32]}
   );
   gpc1_1 gpc2457 (
      {stage1_2[50]},
      {stage2_2[33]}
   );
   gpc1_1 gpc2458 (
      {stage1_2[51]},
      {stage2_2[34]}
   );
   gpc1_1 gpc2459 (
      {stage1_2[52]},
      {stage2_2[35]}
   );
   gpc1_1 gpc2460 (
      {stage1_2[53]},
      {stage2_2[36]}
   );
   gpc1_1 gpc2461 (
      {stage1_2[54]},
      {stage2_2[37]}
   );
   gpc1_1 gpc2462 (
      {stage1_4[66]},
      {stage2_4[31]}
   );
   gpc1_1 gpc2463 (
      {stage1_4[67]},
      {stage2_4[32]}
   );
   gpc1_1 gpc2464 (
      {stage1_4[68]},
      {stage2_4[33]}
   );
   gpc1_1 gpc2465 (
      {stage1_4[69]},
      {stage2_4[34]}
   );
   gpc1_1 gpc2466 (
      {stage1_4[70]},
      {stage2_4[35]}
   );
   gpc1_1 gpc2467 (
      {stage1_4[71]},
      {stage2_4[36]}
   );
   gpc1_1 gpc2468 (
      {stage1_4[72]},
      {stage2_4[37]}
   );
   gpc1_1 gpc2469 (
      {stage1_4[73]},
      {stage2_4[38]}
   );
   gpc1_1 gpc2470 (
      {stage1_4[74]},
      {stage2_4[39]}
   );
   gpc1_1 gpc2471 (
      {stage1_4[75]},
      {stage2_4[40]}
   );
   gpc1_1 gpc2472 (
      {stage1_4[76]},
      {stage2_4[41]}
   );
   gpc1_1 gpc2473 (
      {stage1_4[77]},
      {stage2_4[42]}
   );
   gpc1_1 gpc2474 (
      {stage1_4[78]},
      {stage2_4[43]}
   );
   gpc1_1 gpc2475 (
      {stage1_4[79]},
      {stage2_4[44]}
   );
   gpc1_1 gpc2476 (
      {stage1_4[80]},
      {stage2_4[45]}
   );
   gpc1_1 gpc2477 (
      {stage1_4[81]},
      {stage2_4[46]}
   );
   gpc1_1 gpc2478 (
      {stage1_4[82]},
      {stage2_4[47]}
   );
   gpc1_1 gpc2479 (
      {stage1_5[109]},
      {stage2_5[30]}
   );
   gpc1_1 gpc2480 (
      {stage1_5[110]},
      {stage2_5[31]}
   );
   gpc1_1 gpc2481 (
      {stage1_5[111]},
      {stage2_5[32]}
   );
   gpc1_1 gpc2482 (
      {stage1_5[112]},
      {stage2_5[33]}
   );
   gpc1_1 gpc2483 (
      {stage1_5[113]},
      {stage2_5[34]}
   );
   gpc1_1 gpc2484 (
      {stage1_5[114]},
      {stage2_5[35]}
   );
   gpc1_1 gpc2485 (
      {stage1_7[64]},
      {stage2_7[34]}
   );
   gpc1_1 gpc2486 (
      {stage1_7[65]},
      {stage2_7[35]}
   );
   gpc1_1 gpc2487 (
      {stage1_7[66]},
      {stage2_7[36]}
   );
   gpc1_1 gpc2488 (
      {stage1_7[67]},
      {stage2_7[37]}
   );
   gpc1_1 gpc2489 (
      {stage1_7[68]},
      {stage2_7[38]}
   );
   gpc1_1 gpc2490 (
      {stage1_7[69]},
      {stage2_7[39]}
   );
   gpc1_1 gpc2491 (
      {stage1_7[70]},
      {stage2_7[40]}
   );
   gpc1_1 gpc2492 (
      {stage1_8[46]},
      {stage2_8[26]}
   );
   gpc1_1 gpc2493 (
      {stage1_8[47]},
      {stage2_8[27]}
   );
   gpc1_1 gpc2494 (
      {stage1_8[48]},
      {stage2_8[28]}
   );
   gpc1_1 gpc2495 (
      {stage1_8[49]},
      {stage2_8[29]}
   );
   gpc1_1 gpc2496 (
      {stage1_8[50]},
      {stage2_8[30]}
   );
   gpc1_1 gpc2497 (
      {stage1_8[51]},
      {stage2_8[31]}
   );
   gpc1_1 gpc2498 (
      {stage1_8[52]},
      {stage2_8[32]}
   );
   gpc1_1 gpc2499 (
      {stage1_8[53]},
      {stage2_8[33]}
   );
   gpc1_1 gpc2500 (
      {stage1_8[54]},
      {stage2_8[34]}
   );
   gpc1_1 gpc2501 (
      {stage1_8[55]},
      {stage2_8[35]}
   );
   gpc1_1 gpc2502 (
      {stage1_8[56]},
      {stage2_8[36]}
   );
   gpc1_1 gpc2503 (
      {stage1_8[57]},
      {stage2_8[37]}
   );
   gpc1_1 gpc2504 (
      {stage1_8[58]},
      {stage2_8[38]}
   );
   gpc1_1 gpc2505 (
      {stage1_8[59]},
      {stage2_8[39]}
   );
   gpc1_1 gpc2506 (
      {stage1_8[60]},
      {stage2_8[40]}
   );
   gpc1_1 gpc2507 (
      {stage1_8[61]},
      {stage2_8[41]}
   );
   gpc1_1 gpc2508 (
      {stage1_8[62]},
      {stage2_8[42]}
   );
   gpc1_1 gpc2509 (
      {stage1_8[63]},
      {stage2_8[43]}
   );
   gpc1_1 gpc2510 (
      {stage1_8[64]},
      {stage2_8[44]}
   );
   gpc1_1 gpc2511 (
      {stage1_8[65]},
      {stage2_8[45]}
   );
   gpc1_1 gpc2512 (
      {stage1_8[66]},
      {stage2_8[46]}
   );
   gpc1_1 gpc2513 (
      {stage1_8[67]},
      {stage2_8[47]}
   );
   gpc1_1 gpc2514 (
      {stage1_8[68]},
      {stage2_8[48]}
   );
   gpc1_1 gpc2515 (
      {stage1_8[69]},
      {stage2_8[49]}
   );
   gpc1_1 gpc2516 (
      {stage1_8[70]},
      {stage2_8[50]}
   );
   gpc1_1 gpc2517 (
      {stage1_8[71]},
      {stage2_8[51]}
   );
   gpc1_1 gpc2518 (
      {stage1_8[72]},
      {stage2_8[52]}
   );
   gpc1_1 gpc2519 (
      {stage1_8[73]},
      {stage2_8[53]}
   );
   gpc1_1 gpc2520 (
      {stage1_8[74]},
      {stage2_8[54]}
   );
   gpc1_1 gpc2521 (
      {stage1_8[75]},
      {stage2_8[55]}
   );
   gpc1_1 gpc2522 (
      {stage1_8[76]},
      {stage2_8[56]}
   );
   gpc1_1 gpc2523 (
      {stage1_8[77]},
      {stage2_8[57]}
   );
   gpc1_1 gpc2524 (
      {stage1_8[78]},
      {stage2_8[58]}
   );
   gpc1_1 gpc2525 (
      {stage1_8[79]},
      {stage2_8[59]}
   );
   gpc1_1 gpc2526 (
      {stage1_8[80]},
      {stage2_8[60]}
   );
   gpc1_1 gpc2527 (
      {stage1_9[54]},
      {stage2_9[22]}
   );
   gpc1_1 gpc2528 (
      {stage1_9[55]},
      {stage2_9[23]}
   );
   gpc1_1 gpc2529 (
      {stage1_9[56]},
      {stage2_9[24]}
   );
   gpc1_1 gpc2530 (
      {stage1_9[57]},
      {stage2_9[25]}
   );
   gpc1_1 gpc2531 (
      {stage1_10[79]},
      {stage2_10[25]}
   );
   gpc1_1 gpc2532 (
      {stage1_10[80]},
      {stage2_10[26]}
   );
   gpc1_1 gpc2533 (
      {stage1_10[81]},
      {stage2_10[27]}
   );
   gpc1_1 gpc2534 (
      {stage1_10[82]},
      {stage2_10[28]}
   );
   gpc1_1 gpc2535 (
      {stage1_10[83]},
      {stage2_10[29]}
   );
   gpc1_1 gpc2536 (
      {stage1_10[84]},
      {stage2_10[30]}
   );
   gpc1_1 gpc2537 (
      {stage1_10[85]},
      {stage2_10[31]}
   );
   gpc1_1 gpc2538 (
      {stage1_10[86]},
      {stage2_10[32]}
   );
   gpc1_1 gpc2539 (
      {stage1_10[87]},
      {stage2_10[33]}
   );
   gpc1_1 gpc2540 (
      {stage1_10[88]},
      {stage2_10[34]}
   );
   gpc1_1 gpc2541 (
      {stage1_10[89]},
      {stage2_10[35]}
   );
   gpc1_1 gpc2542 (
      {stage1_10[90]},
      {stage2_10[36]}
   );
   gpc1_1 gpc2543 (
      {stage1_10[91]},
      {stage2_10[37]}
   );
   gpc1_1 gpc2544 (
      {stage1_10[92]},
      {stage2_10[38]}
   );
   gpc1_1 gpc2545 (
      {stage1_10[93]},
      {stage2_10[39]}
   );
   gpc1_1 gpc2546 (
      {stage1_10[94]},
      {stage2_10[40]}
   );
   gpc1_1 gpc2547 (
      {stage1_11[74]},
      {stage2_11[32]}
   );
   gpc1_1 gpc2548 (
      {stage1_11[75]},
      {stage2_11[33]}
   );
   gpc1_1 gpc2549 (
      {stage1_11[76]},
      {stage2_11[34]}
   );
   gpc1_1 gpc2550 (
      {stage1_11[77]},
      {stage2_11[35]}
   );
   gpc1_1 gpc2551 (
      {stage1_11[78]},
      {stage2_11[36]}
   );
   gpc1_1 gpc2552 (
      {stage1_11[79]},
      {stage2_11[37]}
   );
   gpc1_1 gpc2553 (
      {stage1_11[80]},
      {stage2_11[38]}
   );
   gpc1_1 gpc2554 (
      {stage1_12[63]},
      {stage2_12[27]}
   );
   gpc1_1 gpc2555 (
      {stage1_12[64]},
      {stage2_12[28]}
   );
   gpc1_1 gpc2556 (
      {stage1_12[65]},
      {stage2_12[29]}
   );
   gpc1_1 gpc2557 (
      {stage1_12[66]},
      {stage2_12[30]}
   );
   gpc1_1 gpc2558 (
      {stage1_13[66]},
      {stage2_13[24]}
   );
   gpc1_1 gpc2559 (
      {stage1_13[67]},
      {stage2_13[25]}
   );
   gpc1_1 gpc2560 (
      {stage1_13[68]},
      {stage2_13[26]}
   );
   gpc1_1 gpc2561 (
      {stage1_13[69]},
      {stage2_13[27]}
   );
   gpc1_1 gpc2562 (
      {stage1_13[70]},
      {stage2_13[28]}
   );
   gpc1_1 gpc2563 (
      {stage1_13[71]},
      {stage2_13[29]}
   );
   gpc1_1 gpc2564 (
      {stage1_13[72]},
      {stage2_13[30]}
   );
   gpc1_1 gpc2565 (
      {stage1_13[73]},
      {stage2_13[31]}
   );
   gpc1_1 gpc2566 (
      {stage1_13[74]},
      {stage2_13[32]}
   );
   gpc1_1 gpc2567 (
      {stage1_13[75]},
      {stage2_13[33]}
   );
   gpc1_1 gpc2568 (
      {stage1_13[76]},
      {stage2_13[34]}
   );
   gpc1_1 gpc2569 (
      {stage1_13[77]},
      {stage2_13[35]}
   );
   gpc1_1 gpc2570 (
      {stage1_13[78]},
      {stage2_13[36]}
   );
   gpc1_1 gpc2571 (
      {stage1_13[79]},
      {stage2_13[37]}
   );
   gpc1_1 gpc2572 (
      {stage1_13[80]},
      {stage2_13[38]}
   );
   gpc1_1 gpc2573 (
      {stage1_13[81]},
      {stage2_13[39]}
   );
   gpc1_1 gpc2574 (
      {stage1_13[82]},
      {stage2_13[40]}
   );
   gpc1_1 gpc2575 (
      {stage1_13[83]},
      {stage2_13[41]}
   );
   gpc1_1 gpc2576 (
      {stage1_13[84]},
      {stage2_13[42]}
   );
   gpc1_1 gpc2577 (
      {stage1_13[85]},
      {stage2_13[43]}
   );
   gpc1_1 gpc2578 (
      {stage1_13[86]},
      {stage2_13[44]}
   );
   gpc1_1 gpc2579 (
      {stage1_14[10]},
      {stage2_14[22]}
   );
   gpc1_1 gpc2580 (
      {stage1_14[11]},
      {stage2_14[23]}
   );
   gpc1_1 gpc2581 (
      {stage1_14[12]},
      {stage2_14[24]}
   );
   gpc1_1 gpc2582 (
      {stage1_14[13]},
      {stage2_14[25]}
   );
   gpc1_1 gpc2583 (
      {stage1_14[14]},
      {stage2_14[26]}
   );
   gpc1_1 gpc2584 (
      {stage1_14[15]},
      {stage2_14[27]}
   );
   gpc1_1 gpc2585 (
      {stage1_14[16]},
      {stage2_14[28]}
   );
   gpc1_1 gpc2586 (
      {stage1_14[17]},
      {stage2_14[29]}
   );
   gpc1_1 gpc2587 (
      {stage1_14[18]},
      {stage2_14[30]}
   );
   gpc1_1 gpc2588 (
      {stage1_14[19]},
      {stage2_14[31]}
   );
   gpc1_1 gpc2589 (
      {stage1_14[20]},
      {stage2_14[32]}
   );
   gpc1_1 gpc2590 (
      {stage1_14[21]},
      {stage2_14[33]}
   );
   gpc1_1 gpc2591 (
      {stage1_14[22]},
      {stage2_14[34]}
   );
   gpc1_1 gpc2592 (
      {stage1_14[23]},
      {stage2_14[35]}
   );
   gpc1_1 gpc2593 (
      {stage1_14[24]},
      {stage2_14[36]}
   );
   gpc1_1 gpc2594 (
      {stage1_14[25]},
      {stage2_14[37]}
   );
   gpc1_1 gpc2595 (
      {stage1_14[26]},
      {stage2_14[38]}
   );
   gpc1_1 gpc2596 (
      {stage1_14[27]},
      {stage2_14[39]}
   );
   gpc1_1 gpc2597 (
      {stage1_14[28]},
      {stage2_14[40]}
   );
   gpc1_1 gpc2598 (
      {stage1_14[29]},
      {stage2_14[41]}
   );
   gpc1_1 gpc2599 (
      {stage1_14[30]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2600 (
      {stage1_14[31]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2601 (
      {stage1_14[32]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2602 (
      {stage1_14[33]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2603 (
      {stage1_14[34]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2604 (
      {stage1_14[35]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2605 (
      {stage1_14[36]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2606 (
      {stage1_14[37]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2607 (
      {stage1_14[38]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2608 (
      {stage1_14[39]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2609 (
      {stage1_14[40]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2610 (
      {stage1_14[41]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2611 (
      {stage1_14[42]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2612 (
      {stage1_14[43]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2613 (
      {stage1_14[44]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2614 (
      {stage1_14[45]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2615 (
      {stage1_14[46]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2616 (
      {stage1_14[47]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2617 (
      {stage1_14[48]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2618 (
      {stage1_14[49]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2619 (
      {stage1_14[50]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2620 (
      {stage1_14[51]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2621 (
      {stage1_14[52]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2622 (
      {stage1_14[53]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2623 (
      {stage1_14[54]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2624 (
      {stage1_14[55]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2625 (
      {stage1_14[56]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2626 (
      {stage1_14[57]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2627 (
      {stage1_14[58]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2628 (
      {stage1_14[59]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2629 (
      {stage1_14[60]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2630 (
      {stage1_14[61]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2631 (
      {stage1_15[86]},
      {stage2_15[25]}
   );
   gpc1_1 gpc2632 (
      {stage1_15[87]},
      {stage2_15[26]}
   );
   gpc1_1 gpc2633 (
      {stage1_15[88]},
      {stage2_15[27]}
   );
   gpc1_1 gpc2634 (
      {stage1_15[89]},
      {stage2_15[28]}
   );
   gpc1_1 gpc2635 (
      {stage1_15[90]},
      {stage2_15[29]}
   );
   gpc1_1 gpc2636 (
      {stage1_15[91]},
      {stage2_15[30]}
   );
   gpc1_1 gpc2637 (
      {stage1_15[92]},
      {stage2_15[31]}
   );
   gpc1_1 gpc2638 (
      {stage1_15[93]},
      {stage2_15[32]}
   );
   gpc1_1 gpc2639 (
      {stage1_15[94]},
      {stage2_15[33]}
   );
   gpc1_1 gpc2640 (
      {stage1_15[95]},
      {stage2_15[34]}
   );
   gpc1_1 gpc2641 (
      {stage1_15[96]},
      {stage2_15[35]}
   );
   gpc1_1 gpc2642 (
      {stage1_15[97]},
      {stage2_15[36]}
   );
   gpc1_1 gpc2643 (
      {stage1_16[42]},
      {stage2_16[21]}
   );
   gpc1_1 gpc2644 (
      {stage1_16[43]},
      {stage2_16[22]}
   );
   gpc1_1 gpc2645 (
      {stage1_16[44]},
      {stage2_16[23]}
   );
   gpc1_1 gpc2646 (
      {stage1_16[45]},
      {stage2_16[24]}
   );
   gpc1_1 gpc2647 (
      {stage1_16[46]},
      {stage2_16[25]}
   );
   gpc1_1 gpc2648 (
      {stage1_16[47]},
      {stage2_16[26]}
   );
   gpc1_1 gpc2649 (
      {stage1_16[48]},
      {stage2_16[27]}
   );
   gpc1_1 gpc2650 (
      {stage1_16[49]},
      {stage2_16[28]}
   );
   gpc1_1 gpc2651 (
      {stage1_16[50]},
      {stage2_16[29]}
   );
   gpc1_1 gpc2652 (
      {stage1_16[51]},
      {stage2_16[30]}
   );
   gpc1_1 gpc2653 (
      {stage1_16[52]},
      {stage2_16[31]}
   );
   gpc1_1 gpc2654 (
      {stage1_16[53]},
      {stage2_16[32]}
   );
   gpc1_1 gpc2655 (
      {stage1_16[54]},
      {stage2_16[33]}
   );
   gpc1_1 gpc2656 (
      {stage1_16[55]},
      {stage2_16[34]}
   );
   gpc1_1 gpc2657 (
      {stage1_16[56]},
      {stage2_16[35]}
   );
   gpc1_1 gpc2658 (
      {stage1_16[57]},
      {stage2_16[36]}
   );
   gpc1_1 gpc2659 (
      {stage1_16[58]},
      {stage2_16[37]}
   );
   gpc1_1 gpc2660 (
      {stage1_16[59]},
      {stage2_16[38]}
   );
   gpc1_1 gpc2661 (
      {stage1_16[60]},
      {stage2_16[39]}
   );
   gpc1_1 gpc2662 (
      {stage1_16[61]},
      {stage2_16[40]}
   );
   gpc1_1 gpc2663 (
      {stage1_16[62]},
      {stage2_16[41]}
   );
   gpc1_1 gpc2664 (
      {stage1_16[63]},
      {stage2_16[42]}
   );
   gpc1_1 gpc2665 (
      {stage1_16[64]},
      {stage2_16[43]}
   );
   gpc1_1 gpc2666 (
      {stage1_16[65]},
      {stage2_16[44]}
   );
   gpc1_1 gpc2667 (
      {stage1_16[66]},
      {stage2_16[45]}
   );
   gpc1_1 gpc2668 (
      {stage1_16[67]},
      {stage2_16[46]}
   );
   gpc1_1 gpc2669 (
      {stage1_17[100]},
      {stage2_17[26]}
   );
   gpc1_1 gpc2670 (
      {stage1_17[101]},
      {stage2_17[27]}
   );
   gpc1_1 gpc2671 (
      {stage1_17[102]},
      {stage2_17[28]}
   );
   gpc1_1 gpc2672 (
      {stage1_17[103]},
      {stage2_17[29]}
   );
   gpc1_1 gpc2673 (
      {stage1_17[104]},
      {stage2_17[30]}
   );
   gpc1_1 gpc2674 (
      {stage1_17[105]},
      {stage2_17[31]}
   );
   gpc1_1 gpc2675 (
      {stage1_17[106]},
      {stage2_17[32]}
   );
   gpc1_1 gpc2676 (
      {stage1_17[107]},
      {stage2_17[33]}
   );
   gpc1_1 gpc2677 (
      {stage1_17[108]},
      {stage2_17[34]}
   );
   gpc1_1 gpc2678 (
      {stage1_17[109]},
      {stage2_17[35]}
   );
   gpc1_1 gpc2679 (
      {stage1_17[110]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2680 (
      {stage1_17[111]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2681 (
      {stage1_17[112]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2682 (
      {stage1_17[113]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2683 (
      {stage1_18[47]},
      {stage2_18[27]}
   );
   gpc1_1 gpc2684 (
      {stage1_18[48]},
      {stage2_18[28]}
   );
   gpc1_1 gpc2685 (
      {stage1_18[49]},
      {stage2_18[29]}
   );
   gpc1_1 gpc2686 (
      {stage1_18[50]},
      {stage2_18[30]}
   );
   gpc1_1 gpc2687 (
      {stage1_18[51]},
      {stage2_18[31]}
   );
   gpc1_1 gpc2688 (
      {stage1_18[52]},
      {stage2_18[32]}
   );
   gpc1_1 gpc2689 (
      {stage1_18[53]},
      {stage2_18[33]}
   );
   gpc1_1 gpc2690 (
      {stage1_18[54]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2691 (
      {stage1_18[55]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2692 (
      {stage1_18[56]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2693 (
      {stage1_18[57]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2694 (
      {stage1_18[58]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2695 (
      {stage1_18[59]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2696 (
      {stage1_18[60]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2697 (
      {stage1_18[61]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2698 (
      {stage1_18[62]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2699 (
      {stage1_19[48]},
      {stage2_19[28]}
   );
   gpc1_1 gpc2700 (
      {stage1_19[49]},
      {stage2_19[29]}
   );
   gpc1_1 gpc2701 (
      {stage1_19[50]},
      {stage2_19[30]}
   );
   gpc1_1 gpc2702 (
      {stage1_19[51]},
      {stage2_19[31]}
   );
   gpc1_1 gpc2703 (
      {stage1_19[52]},
      {stage2_19[32]}
   );
   gpc1_1 gpc2704 (
      {stage1_19[53]},
      {stage2_19[33]}
   );
   gpc1_1 gpc2705 (
      {stage1_19[54]},
      {stage2_19[34]}
   );
   gpc1_1 gpc2706 (
      {stage1_19[55]},
      {stage2_19[35]}
   );
   gpc1_1 gpc2707 (
      {stage1_19[56]},
      {stage2_19[36]}
   );
   gpc1_1 gpc2708 (
      {stage1_19[57]},
      {stage2_19[37]}
   );
   gpc1_1 gpc2709 (
      {stage1_19[58]},
      {stage2_19[38]}
   );
   gpc1_1 gpc2710 (
      {stage1_19[59]},
      {stage2_19[39]}
   );
   gpc1_1 gpc2711 (
      {stage1_19[60]},
      {stage2_19[40]}
   );
   gpc1_1 gpc2712 (
      {stage1_19[61]},
      {stage2_19[41]}
   );
   gpc1_1 gpc2713 (
      {stage1_19[62]},
      {stage2_19[42]}
   );
   gpc1_1 gpc2714 (
      {stage1_19[63]},
      {stage2_19[43]}
   );
   gpc1_1 gpc2715 (
      {stage1_19[64]},
      {stage2_19[44]}
   );
   gpc1_1 gpc2716 (
      {stage1_19[65]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2717 (
      {stage1_19[66]},
      {stage2_19[46]}
   );
   gpc1_1 gpc2718 (
      {stage1_19[67]},
      {stage2_19[47]}
   );
   gpc1_1 gpc2719 (
      {stage1_19[68]},
      {stage2_19[48]}
   );
   gpc1_1 gpc2720 (
      {stage1_19[69]},
      {stage2_19[49]}
   );
   gpc1_1 gpc2721 (
      {stage1_19[70]},
      {stage2_19[50]}
   );
   gpc1_1 gpc2722 (
      {stage1_20[27]},
      {stage2_20[17]}
   );
   gpc1_1 gpc2723 (
      {stage1_20[28]},
      {stage2_20[18]}
   );
   gpc1_1 gpc2724 (
      {stage1_20[29]},
      {stage2_20[19]}
   );
   gpc1_1 gpc2725 (
      {stage1_20[30]},
      {stage2_20[20]}
   );
   gpc1_1 gpc2726 (
      {stage1_20[31]},
      {stage2_20[21]}
   );
   gpc1_1 gpc2727 (
      {stage1_20[32]},
      {stage2_20[22]}
   );
   gpc1_1 gpc2728 (
      {stage1_20[33]},
      {stage2_20[23]}
   );
   gpc1_1 gpc2729 (
      {stage1_20[34]},
      {stage2_20[24]}
   );
   gpc1_1 gpc2730 (
      {stage1_20[35]},
      {stage2_20[25]}
   );
   gpc1_1 gpc2731 (
      {stage1_20[36]},
      {stage2_20[26]}
   );
   gpc1_1 gpc2732 (
      {stage1_20[37]},
      {stage2_20[27]}
   );
   gpc1_1 gpc2733 (
      {stage1_20[38]},
      {stage2_20[28]}
   );
   gpc1_1 gpc2734 (
      {stage1_20[39]},
      {stage2_20[29]}
   );
   gpc1_1 gpc2735 (
      {stage1_20[40]},
      {stage2_20[30]}
   );
   gpc1_1 gpc2736 (
      {stage1_20[41]},
      {stage2_20[31]}
   );
   gpc1_1 gpc2737 (
      {stage1_20[42]},
      {stage2_20[32]}
   );
   gpc1_1 gpc2738 (
      {stage1_20[43]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2739 (
      {stage1_20[44]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2740 (
      {stage1_20[45]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2741 (
      {stage1_20[46]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2742 (
      {stage1_20[47]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2743 (
      {stage1_20[48]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2744 (
      {stage1_20[49]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2745 (
      {stage1_20[50]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2746 (
      {stage1_20[51]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2747 (
      {stage1_20[52]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2748 (
      {stage1_20[53]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2749 (
      {stage1_20[54]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2750 (
      {stage1_20[55]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2751 (
      {stage1_20[56]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2752 (
      {stage1_20[57]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2753 (
      {stage1_20[58]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2754 (
      {stage1_20[59]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2755 (
      {stage1_20[60]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2756 (
      {stage1_20[61]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2757 (
      {stage1_20[62]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2758 (
      {stage1_20[63]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2759 (
      {stage1_20[64]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2760 (
      {stage1_20[65]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2761 (
      {stage1_20[66]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2762 (
      {stage1_20[67]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2763 (
      {stage1_21[48]},
      {stage2_21[17]}
   );
   gpc1_1 gpc2764 (
      {stage1_21[49]},
      {stage2_21[18]}
   );
   gpc1_1 gpc2765 (
      {stage1_21[50]},
      {stage2_21[19]}
   );
   gpc1_1 gpc2766 (
      {stage1_21[51]},
      {stage2_21[20]}
   );
   gpc1_1 gpc2767 (
      {stage1_21[52]},
      {stage2_21[21]}
   );
   gpc1_1 gpc2768 (
      {stage1_21[53]},
      {stage2_21[22]}
   );
   gpc1_1 gpc2769 (
      {stage1_21[54]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2770 (
      {stage1_21[55]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2771 (
      {stage1_21[56]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2772 (
      {stage1_21[57]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2773 (
      {stage1_21[58]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2774 (
      {stage1_21[59]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2775 (
      {stage1_21[60]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2776 (
      {stage1_21[61]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2777 (
      {stage1_21[62]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2778 (
      {stage1_21[63]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2779 (
      {stage1_21[64]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2780 (
      {stage1_21[65]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2781 (
      {stage1_21[66]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2782 (
      {stage1_21[67]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2783 (
      {stage1_21[68]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2784 (
      {stage1_21[69]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2785 (
      {stage1_21[70]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2786 (
      {stage1_22[62]},
      {stage2_22[26]}
   );
   gpc1_1 gpc2787 (
      {stage1_22[63]},
      {stage2_22[27]}
   );
   gpc1_1 gpc2788 (
      {stage1_22[64]},
      {stage2_22[28]}
   );
   gpc1_1 gpc2789 (
      {stage1_22[65]},
      {stage2_22[29]}
   );
   gpc1_1 gpc2790 (
      {stage1_22[66]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2791 (
      {stage1_23[127]},
      {stage2_23[31]}
   );
   gpc1_1 gpc2792 (
      {stage1_23[128]},
      {stage2_23[32]}
   );
   gpc1_1 gpc2793 (
      {stage1_23[129]},
      {stage2_23[33]}
   );
   gpc1_1 gpc2794 (
      {stage1_23[130]},
      {stage2_23[34]}
   );
   gpc1_1 gpc2795 (
      {stage1_23[131]},
      {stage2_23[35]}
   );
   gpc1_1 gpc2796 (
      {stage1_23[132]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2797 (
      {stage1_23[133]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2798 (
      {stage1_23[134]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2799 (
      {stage1_23[135]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2800 (
      {stage1_23[136]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2801 (
      {stage1_23[137]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2802 (
      {stage1_23[138]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2803 (
      {stage1_23[139]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2804 (
      {stage1_23[140]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2805 (
      {stage1_23[141]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2806 (
      {stage1_23[142]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2807 (
      {stage1_24[69]},
      {stage2_24[32]}
   );
   gpc1_1 gpc2808 (
      {stage1_24[70]},
      {stage2_24[33]}
   );
   gpc1_1 gpc2809 (
      {stage1_24[71]},
      {stage2_24[34]}
   );
   gpc1_1 gpc2810 (
      {stage1_24[72]},
      {stage2_24[35]}
   );
   gpc1_1 gpc2811 (
      {stage1_24[73]},
      {stage2_24[36]}
   );
   gpc1_1 gpc2812 (
      {stage1_24[74]},
      {stage2_24[37]}
   );
   gpc1_1 gpc2813 (
      {stage1_24[75]},
      {stage2_24[38]}
   );
   gpc1_1 gpc2814 (
      {stage1_24[76]},
      {stage2_24[39]}
   );
   gpc1_1 gpc2815 (
      {stage1_24[77]},
      {stage2_24[40]}
   );
   gpc1_1 gpc2816 (
      {stage1_24[78]},
      {stage2_24[41]}
   );
   gpc1_1 gpc2817 (
      {stage1_24[79]},
      {stage2_24[42]}
   );
   gpc1_1 gpc2818 (
      {stage1_24[80]},
      {stage2_24[43]}
   );
   gpc1_1 gpc2819 (
      {stage1_24[81]},
      {stage2_24[44]}
   );
   gpc1_1 gpc2820 (
      {stage1_24[82]},
      {stage2_24[45]}
   );
   gpc1_1 gpc2821 (
      {stage1_25[83]},
      {stage2_25[35]}
   );
   gpc1_1 gpc2822 (
      {stage1_25[84]},
      {stage2_25[36]}
   );
   gpc1_1 gpc2823 (
      {stage1_26[54]},
      {stage2_26[35]}
   );
   gpc1_1 gpc2824 (
      {stage1_26[55]},
      {stage2_26[36]}
   );
   gpc1_1 gpc2825 (
      {stage1_26[56]},
      {stage2_26[37]}
   );
   gpc1_1 gpc2826 (
      {stage1_26[57]},
      {stage2_26[38]}
   );
   gpc1_1 gpc2827 (
      {stage1_26[58]},
      {stage2_26[39]}
   );
   gpc1_1 gpc2828 (
      {stage1_26[59]},
      {stage2_26[40]}
   );
   gpc1_1 gpc2829 (
      {stage1_26[60]},
      {stage2_26[41]}
   );
   gpc1_1 gpc2830 (
      {stage1_26[61]},
      {stage2_26[42]}
   );
   gpc1_1 gpc2831 (
      {stage1_26[62]},
      {stage2_26[43]}
   );
   gpc1_1 gpc2832 (
      {stage1_26[63]},
      {stage2_26[44]}
   );
   gpc1_1 gpc2833 (
      {stage1_26[64]},
      {stage2_26[45]}
   );
   gpc1_1 gpc2834 (
      {stage1_26[65]},
      {stage2_26[46]}
   );
   gpc1_1 gpc2835 (
      {stage1_26[66]},
      {stage2_26[47]}
   );
   gpc1_1 gpc2836 (
      {stage1_26[67]},
      {stage2_26[48]}
   );
   gpc1_1 gpc2837 (
      {stage1_26[68]},
      {stage2_26[49]}
   );
   gpc1_1 gpc2838 (
      {stage1_26[69]},
      {stage2_26[50]}
   );
   gpc1_1 gpc2839 (
      {stage1_26[70]},
      {stage2_26[51]}
   );
   gpc1_1 gpc2840 (
      {stage1_26[71]},
      {stage2_26[52]}
   );
   gpc1_1 gpc2841 (
      {stage1_27[49]},
      {stage2_27[25]}
   );
   gpc1_1 gpc2842 (
      {stage1_27[50]},
      {stage2_27[26]}
   );
   gpc1_1 gpc2843 (
      {stage1_27[51]},
      {stage2_27[27]}
   );
   gpc1_1 gpc2844 (
      {stage1_27[52]},
      {stage2_27[28]}
   );
   gpc1_1 gpc2845 (
      {stage1_27[53]},
      {stage2_27[29]}
   );
   gpc1_1 gpc2846 (
      {stage1_27[54]},
      {stage2_27[30]}
   );
   gpc1_1 gpc2847 (
      {stage1_27[55]},
      {stage2_27[31]}
   );
   gpc1_1 gpc2848 (
      {stage1_27[56]},
      {stage2_27[32]}
   );
   gpc1_1 gpc2849 (
      {stage1_27[57]},
      {stage2_27[33]}
   );
   gpc1_1 gpc2850 (
      {stage1_27[58]},
      {stage2_27[34]}
   );
   gpc1_1 gpc2851 (
      {stage1_27[59]},
      {stage2_27[35]}
   );
   gpc1_1 gpc2852 (
      {stage1_27[60]},
      {stage2_27[36]}
   );
   gpc1_1 gpc2853 (
      {stage1_27[61]},
      {stage2_27[37]}
   );
   gpc1_1 gpc2854 (
      {stage1_27[62]},
      {stage2_27[38]}
   );
   gpc1_1 gpc2855 (
      {stage1_27[63]},
      {stage2_27[39]}
   );
   gpc1_1 gpc2856 (
      {stage1_27[64]},
      {stage2_27[40]}
   );
   gpc1_1 gpc2857 (
      {stage1_27[65]},
      {stage2_27[41]}
   );
   gpc1_1 gpc2858 (
      {stage1_27[66]},
      {stage2_27[42]}
   );
   gpc1_1 gpc2859 (
      {stage1_27[67]},
      {stage2_27[43]}
   );
   gpc1_1 gpc2860 (
      {stage1_27[68]},
      {stage2_27[44]}
   );
   gpc1_1 gpc2861 (
      {stage1_27[69]},
      {stage2_27[45]}
   );
   gpc1_1 gpc2862 (
      {stage1_27[70]},
      {stage2_27[46]}
   );
   gpc1_1 gpc2863 (
      {stage1_27[71]},
      {stage2_27[47]}
   );
   gpc1_1 gpc2864 (
      {stage1_27[72]},
      {stage2_27[48]}
   );
   gpc1_1 gpc2865 (
      {stage1_27[73]},
      {stage2_27[49]}
   );
   gpc1_1 gpc2866 (
      {stage1_28[69]},
      {stage2_28[27]}
   );
   gpc1_1 gpc2867 (
      {stage1_28[70]},
      {stage2_28[28]}
   );
   gpc1_1 gpc2868 (
      {stage1_28[71]},
      {stage2_28[29]}
   );
   gpc1_1 gpc2869 (
      {stage1_28[72]},
      {stage2_28[30]}
   );
   gpc1_1 gpc2870 (
      {stage1_28[73]},
      {stage2_28[31]}
   );
   gpc1_1 gpc2871 (
      {stage1_28[74]},
      {stage2_28[32]}
   );
   gpc1_1 gpc2872 (
      {stage1_28[75]},
      {stage2_28[33]}
   );
   gpc1_1 gpc2873 (
      {stage1_28[76]},
      {stage2_28[34]}
   );
   gpc1_1 gpc2874 (
      {stage1_29[58]},
      {stage2_29[27]}
   );
   gpc1_1 gpc2875 (
      {stage1_29[59]},
      {stage2_29[28]}
   );
   gpc1_1 gpc2876 (
      {stage1_29[60]},
      {stage2_29[29]}
   );
   gpc1_1 gpc2877 (
      {stage1_29[61]},
      {stage2_29[30]}
   );
   gpc1_1 gpc2878 (
      {stage1_29[62]},
      {stage2_29[31]}
   );
   gpc1_1 gpc2879 (
      {stage1_29[63]},
      {stage2_29[32]}
   );
   gpc1_1 gpc2880 (
      {stage1_29[64]},
      {stage2_29[33]}
   );
   gpc1_1 gpc2881 (
      {stage1_29[65]},
      {stage2_29[34]}
   );
   gpc1_1 gpc2882 (
      {stage1_29[66]},
      {stage2_29[35]}
   );
   gpc1_1 gpc2883 (
      {stage1_29[67]},
      {stage2_29[36]}
   );
   gpc1_1 gpc2884 (
      {stage1_29[68]},
      {stage2_29[37]}
   );
   gpc1_1 gpc2885 (
      {stage1_29[69]},
      {stage2_29[38]}
   );
   gpc1_1 gpc2886 (
      {stage1_29[70]},
      {stage2_29[39]}
   );
   gpc1_1 gpc2887 (
      {stage1_29[71]},
      {stage2_29[40]}
   );
   gpc1_1 gpc2888 (
      {stage1_29[72]},
      {stage2_29[41]}
   );
   gpc1_1 gpc2889 (
      {stage1_29[73]},
      {stage2_29[42]}
   );
   gpc1_1 gpc2890 (
      {stage1_29[74]},
      {stage2_29[43]}
   );
   gpc1_1 gpc2891 (
      {stage1_29[75]},
      {stage2_29[44]}
   );
   gpc1_1 gpc2892 (
      {stage1_29[76]},
      {stage2_29[45]}
   );
   gpc1_1 gpc2893 (
      {stage1_29[77]},
      {stage2_29[46]}
   );
   gpc1_1 gpc2894 (
      {stage1_29[78]},
      {stage2_29[47]}
   );
   gpc1_1 gpc2895 (
      {stage1_29[79]},
      {stage2_29[48]}
   );
   gpc1_1 gpc2896 (
      {stage1_29[80]},
      {stage2_29[49]}
   );
   gpc1_1 gpc2897 (
      {stage1_30[84]},
      {stage2_30[27]}
   );
   gpc1_1 gpc2898 (
      {stage1_30[85]},
      {stage2_30[28]}
   );
   gpc1_1 gpc2899 (
      {stage1_30[86]},
      {stage2_30[29]}
   );
   gpc1_1 gpc2900 (
      {stage1_30[87]},
      {stage2_30[30]}
   );
   gpc1_1 gpc2901 (
      {stage1_30[88]},
      {stage2_30[31]}
   );
   gpc1_1 gpc2902 (
      {stage1_30[89]},
      {stage2_30[32]}
   );
   gpc1_1 gpc2903 (
      {stage1_30[90]},
      {stage2_30[33]}
   );
   gpc1_1 gpc2904 (
      {stage1_30[91]},
      {stage2_30[34]}
   );
   gpc1_1 gpc2905 (
      {stage1_30[92]},
      {stage2_30[35]}
   );
   gpc1_1 gpc2906 (
      {stage1_30[93]},
      {stage2_30[36]}
   );
   gpc1_1 gpc2907 (
      {stage1_30[94]},
      {stage2_30[37]}
   );
   gpc1_1 gpc2908 (
      {stage1_30[95]},
      {stage2_30[38]}
   );
   gpc1_1 gpc2909 (
      {stage1_30[96]},
      {stage2_30[39]}
   );
   gpc1_1 gpc2910 (
      {stage1_30[97]},
      {stage2_30[40]}
   );
   gpc1_1 gpc2911 (
      {stage1_30[98]},
      {stage2_30[41]}
   );
   gpc1_1 gpc2912 (
      {stage1_30[99]},
      {stage2_30[42]}
   );
   gpc1_1 gpc2913 (
      {stage1_30[100]},
      {stage2_30[43]}
   );
   gpc1_1 gpc2914 (
      {stage1_30[101]},
      {stage2_30[44]}
   );
   gpc1_1 gpc2915 (
      {stage1_30[102]},
      {stage2_30[45]}
   );
   gpc1_1 gpc2916 (
      {stage1_30[103]},
      {stage2_30[46]}
   );
   gpc1_1 gpc2917 (
      {stage1_30[104]},
      {stage2_30[47]}
   );
   gpc1_1 gpc2918 (
      {stage1_30[105]},
      {stage2_30[48]}
   );
   gpc1_1 gpc2919 (
      {stage1_30[106]},
      {stage2_30[49]}
   );
   gpc1_1 gpc2920 (
      {stage1_31[94]},
      {stage2_31[36]}
   );
   gpc1_1 gpc2921 (
      {stage1_31[95]},
      {stage2_31[37]}
   );
   gpc1_1 gpc2922 (
      {stage1_31[96]},
      {stage2_31[38]}
   );
   gpc1_1 gpc2923 (
      {stage1_32[68]},
      {stage2_32[37]}
   );
   gpc1_1 gpc2924 (
      {stage1_32[69]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2925 (
      {stage1_32[70]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2926 (
      {stage1_32[71]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2927 (
      {stage1_32[72]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2928 (
      {stage1_32[73]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2929 (
      {stage1_32[74]},
      {stage2_32[43]}
   );
   gpc1_1 gpc2930 (
      {stage1_32[75]},
      {stage2_32[44]}
   );
   gpc1_1 gpc2931 (
      {stage1_32[76]},
      {stage2_32[45]}
   );
   gpc1_1 gpc2932 (
      {stage1_32[77]},
      {stage2_32[46]}
   );
   gpc1_1 gpc2933 (
      {stage1_32[78]},
      {stage2_32[47]}
   );
   gpc1_1 gpc2934 (
      {stage1_32[79]},
      {stage2_32[48]}
   );
   gpc1_1 gpc2935 (
      {stage1_32[80]},
      {stage2_32[49]}
   );
   gpc1_1 gpc2936 (
      {stage1_32[81]},
      {stage2_32[50]}
   );
   gpc1_1 gpc2937 (
      {stage1_32[82]},
      {stage2_32[51]}
   );
   gpc1_1 gpc2938 (
      {stage1_32[83]},
      {stage2_32[52]}
   );
   gpc1_1 gpc2939 (
      {stage1_32[84]},
      {stage2_32[53]}
   );
   gpc1_1 gpc2940 (
      {stage1_32[85]},
      {stage2_32[54]}
   );
   gpc1_1 gpc2941 (
      {stage1_32[86]},
      {stage2_32[55]}
   );
   gpc1_1 gpc2942 (
      {stage1_34[48]},
      {stage2_34[27]}
   );
   gpc1_1 gpc2943 (
      {stage1_34[49]},
      {stage2_34[28]}
   );
   gpc1_1 gpc2944 (
      {stage1_34[50]},
      {stage2_34[29]}
   );
   gpc1_1 gpc2945 (
      {stage1_34[51]},
      {stage2_34[30]}
   );
   gpc1_1 gpc2946 (
      {stage1_34[52]},
      {stage2_34[31]}
   );
   gpc1_1 gpc2947 (
      {stage1_34[53]},
      {stage2_34[32]}
   );
   gpc1_1 gpc2948 (
      {stage1_34[54]},
      {stage2_34[33]}
   );
   gpc1_1 gpc2949 (
      {stage1_34[55]},
      {stage2_34[34]}
   );
   gpc1_1 gpc2950 (
      {stage1_35[46]},
      {stage2_35[31]}
   );
   gpc1_1 gpc2951 (
      {stage1_35[47]},
      {stage2_35[32]}
   );
   gpc1_1 gpc2952 (
      {stage1_35[48]},
      {stage2_35[33]}
   );
   gpc1_1 gpc2953 (
      {stage1_35[49]},
      {stage2_35[34]}
   );
   gpc1_1 gpc2954 (
      {stage1_35[50]},
      {stage2_35[35]}
   );
   gpc1_1 gpc2955 (
      {stage1_35[51]},
      {stage2_35[36]}
   );
   gpc1_1 gpc2956 (
      {stage1_35[52]},
      {stage2_35[37]}
   );
   gpc1_1 gpc2957 (
      {stage1_35[53]},
      {stage2_35[38]}
   );
   gpc1_1 gpc2958 (
      {stage1_35[54]},
      {stage2_35[39]}
   );
   gpc1_1 gpc2959 (
      {stage1_35[55]},
      {stage2_35[40]}
   );
   gpc1_1 gpc2960 (
      {stage1_35[56]},
      {stage2_35[41]}
   );
   gpc1_1 gpc2961 (
      {stage1_35[57]},
      {stage2_35[42]}
   );
   gpc1_1 gpc2962 (
      {stage1_35[58]},
      {stage2_35[43]}
   );
   gpc1_1 gpc2963 (
      {stage1_35[59]},
      {stage2_35[44]}
   );
   gpc1_1 gpc2964 (
      {stage1_36[72]},
      {stage2_36[26]}
   );
   gpc1_1 gpc2965 (
      {stage1_36[73]},
      {stage2_36[27]}
   );
   gpc1_1 gpc2966 (
      {stage1_36[74]},
      {stage2_36[28]}
   );
   gpc1_1 gpc2967 (
      {stage1_36[75]},
      {stage2_36[29]}
   );
   gpc1_1 gpc2968 (
      {stage1_36[76]},
      {stage2_36[30]}
   );
   gpc1_1 gpc2969 (
      {stage1_36[77]},
      {stage2_36[31]}
   );
   gpc1_1 gpc2970 (
      {stage1_36[78]},
      {stage2_36[32]}
   );
   gpc1_1 gpc2971 (
      {stage1_36[79]},
      {stage2_36[33]}
   );
   gpc1_1 gpc2972 (
      {stage1_36[80]},
      {stage2_36[34]}
   );
   gpc1_1 gpc2973 (
      {stage1_36[81]},
      {stage2_36[35]}
   );
   gpc1_1 gpc2974 (
      {stage1_36[82]},
      {stage2_36[36]}
   );
   gpc1_1 gpc2975 (
      {stage1_37[117]},
      {stage2_37[31]}
   );
   gpc1_1 gpc2976 (
      {stage1_37[118]},
      {stage2_37[32]}
   );
   gpc1_1 gpc2977 (
      {stage1_37[119]},
      {stage2_37[33]}
   );
   gpc1_1 gpc2978 (
      {stage1_37[120]},
      {stage2_37[34]}
   );
   gpc1_1 gpc2979 (
      {stage1_37[121]},
      {stage2_37[35]}
   );
   gpc1_1 gpc2980 (
      {stage1_37[122]},
      {stage2_37[36]}
   );
   gpc1_1 gpc2981 (
      {stage1_37[123]},
      {stage2_37[37]}
   );
   gpc1_1 gpc2982 (
      {stage1_37[124]},
      {stage2_37[38]}
   );
   gpc1_1 gpc2983 (
      {stage1_37[125]},
      {stage2_37[39]}
   );
   gpc1_1 gpc2984 (
      {stage1_37[126]},
      {stage2_37[40]}
   );
   gpc1_1 gpc2985 (
      {stage1_37[127]},
      {stage2_37[41]}
   );
   gpc1_1 gpc2986 (
      {stage1_39[64]},
      {stage2_39[30]}
   );
   gpc1_1 gpc2987 (
      {stage1_39[65]},
      {stage2_39[31]}
   );
   gpc1_1 gpc2988 (
      {stage1_39[66]},
      {stage2_39[32]}
   );
   gpc1_1 gpc2989 (
      {stage1_39[67]},
      {stage2_39[33]}
   );
   gpc1_1 gpc2990 (
      {stage1_40[72]},
      {stage2_40[31]}
   );
   gpc1_1 gpc2991 (
      {stage1_40[73]},
      {stage2_40[32]}
   );
   gpc1_1 gpc2992 (
      {stage1_40[74]},
      {stage2_40[33]}
   );
   gpc1_1 gpc2993 (
      {stage1_40[75]},
      {stage2_40[34]}
   );
   gpc1_1 gpc2994 (
      {stage1_40[76]},
      {stage2_40[35]}
   );
   gpc1_1 gpc2995 (
      {stage1_40[77]},
      {stage2_40[36]}
   );
   gpc1_1 gpc2996 (
      {stage1_40[78]},
      {stage2_40[37]}
   );
   gpc1_1 gpc2997 (
      {stage1_40[79]},
      {stage2_40[38]}
   );
   gpc1_1 gpc2998 (
      {stage1_40[80]},
      {stage2_40[39]}
   );
   gpc1_1 gpc2999 (
      {stage1_40[81]},
      {stage2_40[40]}
   );
   gpc1_1 gpc3000 (
      {stage1_41[48]},
      {stage2_41[30]}
   );
   gpc1_1 gpc3001 (
      {stage1_41[49]},
      {stage2_41[31]}
   );
   gpc1_1 gpc3002 (
      {stage1_41[50]},
      {stage2_41[32]}
   );
   gpc1_1 gpc3003 (
      {stage1_41[51]},
      {stage2_41[33]}
   );
   gpc1_1 gpc3004 (
      {stage1_41[52]},
      {stage2_41[34]}
   );
   gpc1_1 gpc3005 (
      {stage1_41[53]},
      {stage2_41[35]}
   );
   gpc1_1 gpc3006 (
      {stage1_41[54]},
      {stage2_41[36]}
   );
   gpc1_1 gpc3007 (
      {stage1_41[55]},
      {stage2_41[37]}
   );
   gpc1_1 gpc3008 (
      {stage1_41[56]},
      {stage2_41[38]}
   );
   gpc1_1 gpc3009 (
      {stage1_41[57]},
      {stage2_41[39]}
   );
   gpc1_1 gpc3010 (
      {stage1_41[58]},
      {stage2_41[40]}
   );
   gpc1_1 gpc3011 (
      {stage1_41[59]},
      {stage2_41[41]}
   );
   gpc1_1 gpc3012 (
      {stage1_41[60]},
      {stage2_41[42]}
   );
   gpc1_1 gpc3013 (
      {stage1_41[61]},
      {stage2_41[43]}
   );
   gpc1_1 gpc3014 (
      {stage1_41[62]},
      {stage2_41[44]}
   );
   gpc1_1 gpc3015 (
      {stage1_41[63]},
      {stage2_41[45]}
   );
   gpc1_1 gpc3016 (
      {stage1_41[64]},
      {stage2_41[46]}
   );
   gpc1_1 gpc3017 (
      {stage1_41[65]},
      {stage2_41[47]}
   );
   gpc1_1 gpc3018 (
      {stage1_41[66]},
      {stage2_41[48]}
   );
   gpc1_1 gpc3019 (
      {stage1_41[67]},
      {stage2_41[49]}
   );
   gpc1_1 gpc3020 (
      {stage1_41[68]},
      {stage2_41[50]}
   );
   gpc1_1 gpc3021 (
      {stage1_41[69]},
      {stage2_41[51]}
   );
   gpc1_1 gpc3022 (
      {stage1_41[70]},
      {stage2_41[52]}
   );
   gpc1_1 gpc3023 (
      {stage1_41[71]},
      {stage2_41[53]}
   );
   gpc1_1 gpc3024 (
      {stage1_41[72]},
      {stage2_41[54]}
   );
   gpc1_1 gpc3025 (
      {stage1_41[73]},
      {stage2_41[55]}
   );
   gpc1_1 gpc3026 (
      {stage1_42[54]},
      {stage2_42[20]}
   );
   gpc1_1 gpc3027 (
      {stage1_42[55]},
      {stage2_42[21]}
   );
   gpc1_1 gpc3028 (
      {stage1_42[56]},
      {stage2_42[22]}
   );
   gpc1_1 gpc3029 (
      {stage1_42[57]},
      {stage2_42[23]}
   );
   gpc1_1 gpc3030 (
      {stage1_42[58]},
      {stage2_42[24]}
   );
   gpc1_1 gpc3031 (
      {stage1_42[59]},
      {stage2_42[25]}
   );
   gpc1_1 gpc3032 (
      {stage1_42[60]},
      {stage2_42[26]}
   );
   gpc1_1 gpc3033 (
      {stage1_42[61]},
      {stage2_42[27]}
   );
   gpc1_1 gpc3034 (
      {stage1_42[62]},
      {stage2_42[28]}
   );
   gpc1_1 gpc3035 (
      {stage1_42[63]},
      {stage2_42[29]}
   );
   gpc1_1 gpc3036 (
      {stage1_42[64]},
      {stage2_42[30]}
   );
   gpc1_1 gpc3037 (
      {stage1_42[65]},
      {stage2_42[31]}
   );
   gpc1_1 gpc3038 (
      {stage1_42[66]},
      {stage2_42[32]}
   );
   gpc1_1 gpc3039 (
      {stage1_42[67]},
      {stage2_42[33]}
   );
   gpc1_1 gpc3040 (
      {stage1_42[68]},
      {stage2_42[34]}
   );
   gpc1_1 gpc3041 (
      {stage1_42[69]},
      {stage2_42[35]}
   );
   gpc1_1 gpc3042 (
      {stage1_42[70]},
      {stage2_42[36]}
   );
   gpc1_1 gpc3043 (
      {stage1_42[71]},
      {stage2_42[37]}
   );
   gpc1_1 gpc3044 (
      {stage1_42[72]},
      {stage2_42[38]}
   );
   gpc1_1 gpc3045 (
      {stage1_42[73]},
      {stage2_42[39]}
   );
   gpc1_1 gpc3046 (
      {stage1_42[74]},
      {stage2_42[40]}
   );
   gpc1_1 gpc3047 (
      {stage1_42[75]},
      {stage2_42[41]}
   );
   gpc1_1 gpc3048 (
      {stage1_42[76]},
      {stage2_42[42]}
   );
   gpc1_1 gpc3049 (
      {stage1_42[77]},
      {stage2_42[43]}
   );
   gpc1_1 gpc3050 (
      {stage1_42[78]},
      {stage2_42[44]}
   );
   gpc1_1 gpc3051 (
      {stage1_42[79]},
      {stage2_42[45]}
   );
   gpc1_1 gpc3052 (
      {stage1_42[80]},
      {stage2_42[46]}
   );
   gpc1_1 gpc3053 (
      {stage1_42[81]},
      {stage2_42[47]}
   );
   gpc1_1 gpc3054 (
      {stage1_42[82]},
      {stage2_42[48]}
   );
   gpc1_1 gpc3055 (
      {stage1_42[83]},
      {stage2_42[49]}
   );
   gpc1_1 gpc3056 (
      {stage1_42[84]},
      {stage2_42[50]}
   );
   gpc1_1 gpc3057 (
      {stage1_42[85]},
      {stage2_42[51]}
   );
   gpc1_1 gpc3058 (
      {stage1_42[86]},
      {stage2_42[52]}
   );
   gpc1_1 gpc3059 (
      {stage1_42[87]},
      {stage2_42[53]}
   );
   gpc1_1 gpc3060 (
      {stage1_42[88]},
      {stage2_42[54]}
   );
   gpc1_1 gpc3061 (
      {stage1_42[89]},
      {stage2_42[55]}
   );
   gpc1_1 gpc3062 (
      {stage1_42[90]},
      {stage2_42[56]}
   );
   gpc1_1 gpc3063 (
      {stage1_42[91]},
      {stage2_42[57]}
   );
   gpc1_1 gpc3064 (
      {stage1_42[92]},
      {stage2_42[58]}
   );
   gpc1_1 gpc3065 (
      {stage1_42[93]},
      {stage2_42[59]}
   );
   gpc1_1 gpc3066 (
      {stage1_42[94]},
      {stage2_42[60]}
   );
   gpc1_1 gpc3067 (
      {stage1_42[95]},
      {stage2_42[61]}
   );
   gpc1_1 gpc3068 (
      {stage1_43[114]},
      {stage2_43[28]}
   );
   gpc1_1 gpc3069 (
      {stage1_43[115]},
      {stage2_43[29]}
   );
   gpc1_1 gpc3070 (
      {stage1_43[116]},
      {stage2_43[30]}
   );
   gpc1_1 gpc3071 (
      {stage1_43[117]},
      {stage2_43[31]}
   );
   gpc1_1 gpc3072 (
      {stage1_43[118]},
      {stage2_43[32]}
   );
   gpc1_1 gpc3073 (
      {stage1_43[119]},
      {stage2_43[33]}
   );
   gpc1_1 gpc3074 (
      {stage1_43[120]},
      {stage2_43[34]}
   );
   gpc1_1 gpc3075 (
      {stage1_43[121]},
      {stage2_43[35]}
   );
   gpc1_1 gpc3076 (
      {stage1_43[122]},
      {stage2_43[36]}
   );
   gpc1_1 gpc3077 (
      {stage1_43[123]},
      {stage2_43[37]}
   );
   gpc1_1 gpc3078 (
      {stage1_43[124]},
      {stage2_43[38]}
   );
   gpc1_1 gpc3079 (
      {stage1_43[125]},
      {stage2_43[39]}
   );
   gpc1_1 gpc3080 (
      {stage1_43[126]},
      {stage2_43[40]}
   );
   gpc1_1 gpc3081 (
      {stage1_43[127]},
      {stage2_43[41]}
   );
   gpc1_1 gpc3082 (
      {stage1_43[128]},
      {stage2_43[42]}
   );
   gpc1_1 gpc3083 (
      {stage1_43[129]},
      {stage2_43[43]}
   );
   gpc1_1 gpc3084 (
      {stage1_43[130]},
      {stage2_43[44]}
   );
   gpc1_1 gpc3085 (
      {stage1_43[131]},
      {stage2_43[45]}
   );
   gpc1_1 gpc3086 (
      {stage1_43[132]},
      {stage2_43[46]}
   );
   gpc1_1 gpc3087 (
      {stage1_43[133]},
      {stage2_43[47]}
   );
   gpc1_1 gpc3088 (
      {stage1_43[134]},
      {stage2_43[48]}
   );
   gpc1_1 gpc3089 (
      {stage1_43[135]},
      {stage2_43[49]}
   );
   gpc1_1 gpc3090 (
      {stage1_43[136]},
      {stage2_43[50]}
   );
   gpc1_1 gpc3091 (
      {stage1_43[137]},
      {stage2_43[51]}
   );
   gpc1_1 gpc3092 (
      {stage1_44[10]},
      {stage2_44[30]}
   );
   gpc1_1 gpc3093 (
      {stage1_44[11]},
      {stage2_44[31]}
   );
   gpc1_1 gpc3094 (
      {stage1_44[12]},
      {stage2_44[32]}
   );
   gpc1_1 gpc3095 (
      {stage1_44[13]},
      {stage2_44[33]}
   );
   gpc1_1 gpc3096 (
      {stage1_44[14]},
      {stage2_44[34]}
   );
   gpc1_1 gpc3097 (
      {stage1_44[15]},
      {stage2_44[35]}
   );
   gpc1_1 gpc3098 (
      {stage1_44[16]},
      {stage2_44[36]}
   );
   gpc1_1 gpc3099 (
      {stage1_44[17]},
      {stage2_44[37]}
   );
   gpc1_1 gpc3100 (
      {stage1_44[18]},
      {stage2_44[38]}
   );
   gpc1_1 gpc3101 (
      {stage1_44[19]},
      {stage2_44[39]}
   );
   gpc1_1 gpc3102 (
      {stage1_44[20]},
      {stage2_44[40]}
   );
   gpc1_1 gpc3103 (
      {stage1_44[21]},
      {stage2_44[41]}
   );
   gpc1_1 gpc3104 (
      {stage1_44[22]},
      {stage2_44[42]}
   );
   gpc1_1 gpc3105 (
      {stage1_44[23]},
      {stage2_44[43]}
   );
   gpc1_1 gpc3106 (
      {stage1_44[24]},
      {stage2_44[44]}
   );
   gpc1_1 gpc3107 (
      {stage1_44[25]},
      {stage2_44[45]}
   );
   gpc1_1 gpc3108 (
      {stage1_44[26]},
      {stage2_44[46]}
   );
   gpc1_1 gpc3109 (
      {stage1_44[27]},
      {stage2_44[47]}
   );
   gpc1_1 gpc3110 (
      {stage1_44[28]},
      {stage2_44[48]}
   );
   gpc1_1 gpc3111 (
      {stage1_44[29]},
      {stage2_44[49]}
   );
   gpc1_1 gpc3112 (
      {stage1_44[30]},
      {stage2_44[50]}
   );
   gpc1_1 gpc3113 (
      {stage1_44[31]},
      {stage2_44[51]}
   );
   gpc1_1 gpc3114 (
      {stage1_44[32]},
      {stage2_44[52]}
   );
   gpc1_1 gpc3115 (
      {stage1_44[33]},
      {stage2_44[53]}
   );
   gpc1_1 gpc3116 (
      {stage1_44[34]},
      {stage2_44[54]}
   );
   gpc1_1 gpc3117 (
      {stage1_44[35]},
      {stage2_44[55]}
   );
   gpc1_1 gpc3118 (
      {stage1_44[36]},
      {stage2_44[56]}
   );
   gpc1_1 gpc3119 (
      {stage1_44[37]},
      {stage2_44[57]}
   );
   gpc1_1 gpc3120 (
      {stage1_44[38]},
      {stage2_44[58]}
   );
   gpc1_1 gpc3121 (
      {stage1_44[39]},
      {stage2_44[59]}
   );
   gpc1_1 gpc3122 (
      {stage1_44[40]},
      {stage2_44[60]}
   );
   gpc1_1 gpc3123 (
      {stage1_44[41]},
      {stage2_44[61]}
   );
   gpc1_1 gpc3124 (
      {stage1_44[42]},
      {stage2_44[62]}
   );
   gpc1_1 gpc3125 (
      {stage1_44[43]},
      {stage2_44[63]}
   );
   gpc1_1 gpc3126 (
      {stage1_44[44]},
      {stage2_44[64]}
   );
   gpc1_1 gpc3127 (
      {stage1_44[45]},
      {stage2_44[65]}
   );
   gpc1_1 gpc3128 (
      {stage1_45[92]},
      {stage2_45[25]}
   );
   gpc1_1 gpc3129 (
      {stage1_46[57]},
      {stage2_46[26]}
   );
   gpc1_1 gpc3130 (
      {stage1_46[58]},
      {stage2_46[27]}
   );
   gpc1_1 gpc3131 (
      {stage1_46[59]},
      {stage2_46[28]}
   );
   gpc1_1 gpc3132 (
      {stage1_46[60]},
      {stage2_46[29]}
   );
   gpc1_1 gpc3133 (
      {stage1_46[61]},
      {stage2_46[30]}
   );
   gpc1_1 gpc3134 (
      {stage1_46[62]},
      {stage2_46[31]}
   );
   gpc1_1 gpc3135 (
      {stage1_46[63]},
      {stage2_46[32]}
   );
   gpc1_1 gpc3136 (
      {stage1_47[39]},
      {stage2_47[27]}
   );
   gpc1_1 gpc3137 (
      {stage1_47[40]},
      {stage2_47[28]}
   );
   gpc1_1 gpc3138 (
      {stage1_47[41]},
      {stage2_47[29]}
   );
   gpc1_1 gpc3139 (
      {stage1_47[42]},
      {stage2_47[30]}
   );
   gpc1_1 gpc3140 (
      {stage1_47[43]},
      {stage2_47[31]}
   );
   gpc1_1 gpc3141 (
      {stage1_47[44]},
      {stage2_47[32]}
   );
   gpc1_1 gpc3142 (
      {stage1_47[45]},
      {stage2_47[33]}
   );
   gpc1_1 gpc3143 (
      {stage1_47[46]},
      {stage2_47[34]}
   );
   gpc1_1 gpc3144 (
      {stage1_47[47]},
      {stage2_47[35]}
   );
   gpc1_1 gpc3145 (
      {stage1_47[48]},
      {stage2_47[36]}
   );
   gpc1_1 gpc3146 (
      {stage1_47[49]},
      {stage2_47[37]}
   );
   gpc1_1 gpc3147 (
      {stage1_47[50]},
      {stage2_47[38]}
   );
   gpc1_1 gpc3148 (
      {stage1_47[51]},
      {stage2_47[39]}
   );
   gpc1_1 gpc3149 (
      {stage1_47[52]},
      {stage2_47[40]}
   );
   gpc1_1 gpc3150 (
      {stage1_47[53]},
      {stage2_47[41]}
   );
   gpc1_1 gpc3151 (
      {stage1_47[54]},
      {stage2_47[42]}
   );
   gpc1_1 gpc3152 (
      {stage1_47[55]},
      {stage2_47[43]}
   );
   gpc1_1 gpc3153 (
      {stage1_47[56]},
      {stage2_47[44]}
   );
   gpc1_1 gpc3154 (
      {stage1_47[57]},
      {stage2_47[45]}
   );
   gpc1_1 gpc3155 (
      {stage1_48[66]},
      {stage2_48[18]}
   );
   gpc1_1 gpc3156 (
      {stage1_48[67]},
      {stage2_48[19]}
   );
   gpc1_1 gpc3157 (
      {stage1_48[68]},
      {stage2_48[20]}
   );
   gpc1_1 gpc3158 (
      {stage1_48[69]},
      {stage2_48[21]}
   );
   gpc1_1 gpc3159 (
      {stage1_48[70]},
      {stage2_48[22]}
   );
   gpc1_1 gpc3160 (
      {stage1_48[71]},
      {stage2_48[23]}
   );
   gpc1_1 gpc3161 (
      {stage1_49[78]},
      {stage2_49[28]}
   );
   gpc1_1 gpc3162 (
      {stage1_49[79]},
      {stage2_49[29]}
   );
   gpc1_1 gpc3163 (
      {stage1_49[80]},
      {stage2_49[30]}
   );
   gpc1_1 gpc3164 (
      {stage1_49[81]},
      {stage2_49[31]}
   );
   gpc1_1 gpc3165 (
      {stage1_49[82]},
      {stage2_49[32]}
   );
   gpc1_1 gpc3166 (
      {stage1_49[83]},
      {stage2_49[33]}
   );
   gpc1_1 gpc3167 (
      {stage1_49[84]},
      {stage2_49[34]}
   );
   gpc1_1 gpc3168 (
      {stage1_49[85]},
      {stage2_49[35]}
   );
   gpc1_1 gpc3169 (
      {stage1_49[86]},
      {stage2_49[36]}
   );
   gpc1_1 gpc3170 (
      {stage1_50[47]},
      {stage2_50[30]}
   );
   gpc1_1 gpc3171 (
      {stage1_50[48]},
      {stage2_50[31]}
   );
   gpc1_1 gpc3172 (
      {stage1_50[49]},
      {stage2_50[32]}
   );
   gpc1_1 gpc3173 (
      {stage1_50[50]},
      {stage2_50[33]}
   );
   gpc1_1 gpc3174 (
      {stage1_50[51]},
      {stage2_50[34]}
   );
   gpc1_1 gpc3175 (
      {stage1_50[52]},
      {stage2_50[35]}
   );
   gpc1_1 gpc3176 (
      {stage1_50[53]},
      {stage2_50[36]}
   );
   gpc1_1 gpc3177 (
      {stage1_50[54]},
      {stage2_50[37]}
   );
   gpc1_1 gpc3178 (
      {stage1_50[55]},
      {stage2_50[38]}
   );
   gpc1_1 gpc3179 (
      {stage1_50[56]},
      {stage2_50[39]}
   );
   gpc1_1 gpc3180 (
      {stage1_50[57]},
      {stage2_50[40]}
   );
   gpc1_1 gpc3181 (
      {stage1_51[93]},
      {stage2_51[24]}
   );
   gpc1_1 gpc3182 (
      {stage1_52[73]},
      {stage2_52[30]}
   );
   gpc1_1 gpc3183 (
      {stage1_52[74]},
      {stage2_52[31]}
   );
   gpc1_1 gpc3184 (
      {stage1_52[75]},
      {stage2_52[32]}
   );
   gpc1_1 gpc3185 (
      {stage1_52[76]},
      {stage2_52[33]}
   );
   gpc1_1 gpc3186 (
      {stage1_53[48]},
      {stage2_53[33]}
   );
   gpc1_1 gpc3187 (
      {stage1_53[49]},
      {stage2_53[34]}
   );
   gpc1_1 gpc3188 (
      {stage1_53[50]},
      {stage2_53[35]}
   );
   gpc1_1 gpc3189 (
      {stage1_53[51]},
      {stage2_53[36]}
   );
   gpc1_1 gpc3190 (
      {stage1_53[52]},
      {stage2_53[37]}
   );
   gpc1_1 gpc3191 (
      {stage1_53[53]},
      {stage2_53[38]}
   );
   gpc1_1 gpc3192 (
      {stage1_53[54]},
      {stage2_53[39]}
   );
   gpc1_1 gpc3193 (
      {stage1_53[55]},
      {stage2_53[40]}
   );
   gpc1_1 gpc3194 (
      {stage1_53[56]},
      {stage2_53[41]}
   );
   gpc1_1 gpc3195 (
      {stage1_53[57]},
      {stage2_53[42]}
   );
   gpc1_1 gpc3196 (
      {stage1_53[58]},
      {stage2_53[43]}
   );
   gpc1_1 gpc3197 (
      {stage1_53[59]},
      {stage2_53[44]}
   );
   gpc1_1 gpc3198 (
      {stage1_53[60]},
      {stage2_53[45]}
   );
   gpc1_1 gpc3199 (
      {stage1_53[61]},
      {stage2_53[46]}
   );
   gpc1_1 gpc3200 (
      {stage1_53[62]},
      {stage2_53[47]}
   );
   gpc1_1 gpc3201 (
      {stage1_53[63]},
      {stage2_53[48]}
   );
   gpc1_1 gpc3202 (
      {stage1_53[64]},
      {stage2_53[49]}
   );
   gpc1_1 gpc3203 (
      {stage1_53[65]},
      {stage2_53[50]}
   );
   gpc1_1 gpc3204 (
      {stage1_54[52]},
      {stage2_54[22]}
   );
   gpc1_1 gpc3205 (
      {stage1_54[53]},
      {stage2_54[23]}
   );
   gpc1_1 gpc3206 (
      {stage1_54[54]},
      {stage2_54[24]}
   );
   gpc1_1 gpc3207 (
      {stage1_54[55]},
      {stage2_54[25]}
   );
   gpc1_1 gpc3208 (
      {stage1_54[56]},
      {stage2_54[26]}
   );
   gpc1_1 gpc3209 (
      {stage1_54[57]},
      {stage2_54[27]}
   );
   gpc1_1 gpc3210 (
      {stage1_55[88]},
      {stage2_55[28]}
   );
   gpc1_1 gpc3211 (
      {stage1_55[89]},
      {stage2_55[29]}
   );
   gpc1_1 gpc3212 (
      {stage1_55[90]},
      {stage2_55[30]}
   );
   gpc1_1 gpc3213 (
      {stage1_55[91]},
      {stage2_55[31]}
   );
   gpc1_1 gpc3214 (
      {stage1_55[92]},
      {stage2_55[32]}
   );
   gpc1_1 gpc3215 (
      {stage1_55[93]},
      {stage2_55[33]}
   );
   gpc1_1 gpc3216 (
      {stage1_55[94]},
      {stage2_55[34]}
   );
   gpc1_1 gpc3217 (
      {stage1_55[95]},
      {stage2_55[35]}
   );
   gpc1_1 gpc3218 (
      {stage1_55[96]},
      {stage2_55[36]}
   );
   gpc1_1 gpc3219 (
      {stage1_55[97]},
      {stage2_55[37]}
   );
   gpc1_1 gpc3220 (
      {stage1_56[58]},
      {stage2_56[31]}
   );
   gpc1_1 gpc3221 (
      {stage1_56[59]},
      {stage2_56[32]}
   );
   gpc1_1 gpc3222 (
      {stage1_56[60]},
      {stage2_56[33]}
   );
   gpc1_1 gpc3223 (
      {stage1_56[61]},
      {stage2_56[34]}
   );
   gpc1_1 gpc3224 (
      {stage1_56[62]},
      {stage2_56[35]}
   );
   gpc1_1 gpc3225 (
      {stage1_56[63]},
      {stage2_56[36]}
   );
   gpc1_1 gpc3226 (
      {stage1_56[64]},
      {stage2_56[37]}
   );
   gpc1_1 gpc3227 (
      {stage1_56[65]},
      {stage2_56[38]}
   );
   gpc1_1 gpc3228 (
      {stage1_56[66]},
      {stage2_56[39]}
   );
   gpc1_1 gpc3229 (
      {stage1_56[67]},
      {stage2_56[40]}
   );
   gpc1_1 gpc3230 (
      {stage1_56[68]},
      {stage2_56[41]}
   );
   gpc1_1 gpc3231 (
      {stage1_56[69]},
      {stage2_56[42]}
   );
   gpc1_1 gpc3232 (
      {stage1_56[70]},
      {stage2_56[43]}
   );
   gpc1_1 gpc3233 (
      {stage1_56[71]},
      {stage2_56[44]}
   );
   gpc1_1 gpc3234 (
      {stage1_56[72]},
      {stage2_56[45]}
   );
   gpc1_1 gpc3235 (
      {stage1_56[73]},
      {stage2_56[46]}
   );
   gpc1_1 gpc3236 (
      {stage1_56[74]},
      {stage2_56[47]}
   );
   gpc1_1 gpc3237 (
      {stage1_56[75]},
      {stage2_56[48]}
   );
   gpc1_1 gpc3238 (
      {stage1_56[76]},
      {stage2_56[49]}
   );
   gpc1_1 gpc3239 (
      {stage1_56[77]},
      {stage2_56[50]}
   );
   gpc1_1 gpc3240 (
      {stage1_56[78]},
      {stage2_56[51]}
   );
   gpc1_1 gpc3241 (
      {stage1_56[79]},
      {stage2_56[52]}
   );
   gpc1_1 gpc3242 (
      {stage1_57[66]},
      {stage2_57[24]}
   );
   gpc1_1 gpc3243 (
      {stage1_57[67]},
      {stage2_57[25]}
   );
   gpc1_1 gpc3244 (
      {stage1_57[68]},
      {stage2_57[26]}
   );
   gpc1_1 gpc3245 (
      {stage1_57[69]},
      {stage2_57[27]}
   );
   gpc1_1 gpc3246 (
      {stage1_57[70]},
      {stage2_57[28]}
   );
   gpc1_1 gpc3247 (
      {stage1_57[71]},
      {stage2_57[29]}
   );
   gpc1_1 gpc3248 (
      {stage1_58[65]},
      {stage2_58[24]}
   );
   gpc1_1 gpc3249 (
      {stage1_58[66]},
      {stage2_58[25]}
   );
   gpc1_1 gpc3250 (
      {stage1_58[67]},
      {stage2_58[26]}
   );
   gpc1_1 gpc3251 (
      {stage1_58[68]},
      {stage2_58[27]}
   );
   gpc1_1 gpc3252 (
      {stage1_58[69]},
      {stage2_58[28]}
   );
   gpc1_1 gpc3253 (
      {stage1_58[70]},
      {stage2_58[29]}
   );
   gpc1_1 gpc3254 (
      {stage1_58[71]},
      {stage2_58[30]}
   );
   gpc1_1 gpc3255 (
      {stage1_58[72]},
      {stage2_58[31]}
   );
   gpc1_1 gpc3256 (
      {stage1_58[73]},
      {stage2_58[32]}
   );
   gpc1_1 gpc3257 (
      {stage1_59[25]},
      {stage2_59[26]}
   );
   gpc1_1 gpc3258 (
      {stage1_59[26]},
      {stage2_59[27]}
   );
   gpc1_1 gpc3259 (
      {stage1_59[27]},
      {stage2_59[28]}
   );
   gpc1_1 gpc3260 (
      {stage1_59[28]},
      {stage2_59[29]}
   );
   gpc1_1 gpc3261 (
      {stage1_59[29]},
      {stage2_59[30]}
   );
   gpc1_1 gpc3262 (
      {stage1_59[30]},
      {stage2_59[31]}
   );
   gpc1_1 gpc3263 (
      {stage1_59[31]},
      {stage2_59[32]}
   );
   gpc1_1 gpc3264 (
      {stage1_59[32]},
      {stage2_59[33]}
   );
   gpc1_1 gpc3265 (
      {stage1_59[33]},
      {stage2_59[34]}
   );
   gpc1_1 gpc3266 (
      {stage1_59[34]},
      {stage2_59[35]}
   );
   gpc1_1 gpc3267 (
      {stage1_59[35]},
      {stage2_59[36]}
   );
   gpc1_1 gpc3268 (
      {stage1_59[36]},
      {stage2_59[37]}
   );
   gpc1_1 gpc3269 (
      {stage1_59[37]},
      {stage2_59[38]}
   );
   gpc1_1 gpc3270 (
      {stage1_59[38]},
      {stage2_59[39]}
   );
   gpc1_1 gpc3271 (
      {stage1_59[39]},
      {stage2_59[40]}
   );
   gpc1_1 gpc3272 (
      {stage1_59[40]},
      {stage2_59[41]}
   );
   gpc1_1 gpc3273 (
      {stage1_59[41]},
      {stage2_59[42]}
   );
   gpc1_1 gpc3274 (
      {stage1_59[42]},
      {stage2_59[43]}
   );
   gpc1_1 gpc3275 (
      {stage1_59[43]},
      {stage2_59[44]}
   );
   gpc1_1 gpc3276 (
      {stage1_59[44]},
      {stage2_59[45]}
   );
   gpc1_1 gpc3277 (
      {stage1_59[45]},
      {stage2_59[46]}
   );
   gpc1_1 gpc3278 (
      {stage1_59[46]},
      {stage2_59[47]}
   );
   gpc1_1 gpc3279 (
      {stage1_59[47]},
      {stage2_59[48]}
   );
   gpc1_1 gpc3280 (
      {stage1_59[48]},
      {stage2_59[49]}
   );
   gpc1_1 gpc3281 (
      {stage1_59[49]},
      {stage2_59[50]}
   );
   gpc1_1 gpc3282 (
      {stage1_59[50]},
      {stage2_59[51]}
   );
   gpc1_1 gpc3283 (
      {stage1_59[51]},
      {stage2_59[52]}
   );
   gpc1_1 gpc3284 (
      {stage1_59[52]},
      {stage2_59[53]}
   );
   gpc1_1 gpc3285 (
      {stage1_59[53]},
      {stage2_59[54]}
   );
   gpc1_1 gpc3286 (
      {stage1_59[54]},
      {stage2_59[55]}
   );
   gpc1_1 gpc3287 (
      {stage1_59[55]},
      {stage2_59[56]}
   );
   gpc1_1 gpc3288 (
      {stage1_59[56]},
      {stage2_59[57]}
   );
   gpc1_1 gpc3289 (
      {stage1_59[57]},
      {stage2_59[58]}
   );
   gpc1_1 gpc3290 (
      {stage1_59[58]},
      {stage2_59[59]}
   );
   gpc1_1 gpc3291 (
      {stage1_59[59]},
      {stage2_59[60]}
   );
   gpc1_1 gpc3292 (
      {stage1_59[60]},
      {stage2_59[61]}
   );
   gpc1_1 gpc3293 (
      {stage1_59[61]},
      {stage2_59[62]}
   );
   gpc1_1 gpc3294 (
      {stage1_59[62]},
      {stage2_59[63]}
   );
   gpc1_1 gpc3295 (
      {stage1_59[63]},
      {stage2_59[64]}
   );
   gpc1_1 gpc3296 (
      {stage1_59[64]},
      {stage2_59[65]}
   );
   gpc1_1 gpc3297 (
      {stage1_59[65]},
      {stage2_59[66]}
   );
   gpc1_1 gpc3298 (
      {stage1_59[66]},
      {stage2_59[67]}
   );
   gpc1_1 gpc3299 (
      {stage1_59[67]},
      {stage2_59[68]}
   );
   gpc1_1 gpc3300 (
      {stage1_59[68]},
      {stage2_59[69]}
   );
   gpc1_1 gpc3301 (
      {stage1_59[69]},
      {stage2_59[70]}
   );
   gpc1_1 gpc3302 (
      {stage1_59[70]},
      {stage2_59[71]}
   );
   gpc1_1 gpc3303 (
      {stage1_59[71]},
      {stage2_59[72]}
   );
   gpc1_1 gpc3304 (
      {stage1_59[72]},
      {stage2_59[73]}
   );
   gpc1_1 gpc3305 (
      {stage1_59[73]},
      {stage2_59[74]}
   );
   gpc1_1 gpc3306 (
      {stage1_59[74]},
      {stage2_59[75]}
   );
   gpc1_1 gpc3307 (
      {stage1_59[75]},
      {stage2_59[76]}
   );
   gpc1_1 gpc3308 (
      {stage1_59[76]},
      {stage2_59[77]}
   );
   gpc1_1 gpc3309 (
      {stage1_59[77]},
      {stage2_59[78]}
   );
   gpc1_1 gpc3310 (
      {stage1_59[78]},
      {stage2_59[79]}
   );
   gpc1_1 gpc3311 (
      {stage1_59[79]},
      {stage2_59[80]}
   );
   gpc1_1 gpc3312 (
      {stage1_60[66]},
      {stage2_60[21]}
   );
   gpc1_1 gpc3313 (
      {stage1_61[42]},
      {stage2_61[18]}
   );
   gpc1_1 gpc3314 (
      {stage1_61[43]},
      {stage2_61[19]}
   );
   gpc1_1 gpc3315 (
      {stage1_61[44]},
      {stage2_61[20]}
   );
   gpc1_1 gpc3316 (
      {stage1_61[45]},
      {stage2_61[21]}
   );
   gpc1_1 gpc3317 (
      {stage1_61[46]},
      {stage2_61[22]}
   );
   gpc1_1 gpc3318 (
      {stage1_61[47]},
      {stage2_61[23]}
   );
   gpc1_1 gpc3319 (
      {stage1_61[48]},
      {stage2_61[24]}
   );
   gpc1_1 gpc3320 (
      {stage1_61[49]},
      {stage2_61[25]}
   );
   gpc1_1 gpc3321 (
      {stage1_61[50]},
      {stage2_61[26]}
   );
   gpc1_1 gpc3322 (
      {stage1_61[51]},
      {stage2_61[27]}
   );
   gpc1_1 gpc3323 (
      {stage1_61[52]},
      {stage2_61[28]}
   );
   gpc1_1 gpc3324 (
      {stage1_61[53]},
      {stage2_61[29]}
   );
   gpc1_1 gpc3325 (
      {stage1_61[54]},
      {stage2_61[30]}
   );
   gpc1_1 gpc3326 (
      {stage1_61[55]},
      {stage2_61[31]}
   );
   gpc1_1 gpc3327 (
      {stage1_61[56]},
      {stage2_61[32]}
   );
   gpc1_1 gpc3328 (
      {stage1_61[57]},
      {stage2_61[33]}
   );
   gpc1_1 gpc3329 (
      {stage1_61[58]},
      {stage2_61[34]}
   );
   gpc1_1 gpc3330 (
      {stage1_61[59]},
      {stage2_61[35]}
   );
   gpc1_1 gpc3331 (
      {stage1_61[60]},
      {stage2_61[36]}
   );
   gpc1_1 gpc3332 (
      {stage1_61[61]},
      {stage2_61[37]}
   );
   gpc1_1 gpc3333 (
      {stage1_61[62]},
      {stage2_61[38]}
   );
   gpc1_1 gpc3334 (
      {stage1_61[63]},
      {stage2_61[39]}
   );
   gpc1_1 gpc3335 (
      {stage1_61[64]},
      {stage2_61[40]}
   );
   gpc1_1 gpc3336 (
      {stage1_61[65]},
      {stage2_61[41]}
   );
   gpc1_1 gpc3337 (
      {stage1_61[66]},
      {stage2_61[42]}
   );
   gpc1_1 gpc3338 (
      {stage1_61[67]},
      {stage2_61[43]}
   );
   gpc1_1 gpc3339 (
      {stage1_61[68]},
      {stage2_61[44]}
   );
   gpc1_1 gpc3340 (
      {stage1_61[69]},
      {stage2_61[45]}
   );
   gpc1_1 gpc3341 (
      {stage1_61[70]},
      {stage2_61[46]}
   );
   gpc1_1 gpc3342 (
      {stage1_61[71]},
      {stage2_61[47]}
   );
   gpc1_1 gpc3343 (
      {stage1_61[72]},
      {stage2_61[48]}
   );
   gpc1_1 gpc3344 (
      {stage1_61[73]},
      {stage2_61[49]}
   );
   gpc1_1 gpc3345 (
      {stage1_61[74]},
      {stage2_61[50]}
   );
   gpc1_1 gpc3346 (
      {stage1_61[75]},
      {stage2_61[51]}
   );
   gpc1_1 gpc3347 (
      {stage1_61[76]},
      {stage2_61[52]}
   );
   gpc1_1 gpc3348 (
      {stage1_61[77]},
      {stage2_61[53]}
   );
   gpc1_1 gpc3349 (
      {stage1_61[78]},
      {stage2_61[54]}
   );
   gpc1_1 gpc3350 (
      {stage1_61[79]},
      {stage2_61[55]}
   );
   gpc1_1 gpc3351 (
      {stage1_61[80]},
      {stage2_61[56]}
   );
   gpc1_1 gpc3352 (
      {stage1_61[81]},
      {stage2_61[57]}
   );
   gpc1_1 gpc3353 (
      {stage1_61[82]},
      {stage2_61[58]}
   );
   gpc1_1 gpc3354 (
      {stage1_61[83]},
      {stage2_61[59]}
   );
   gpc1_1 gpc3355 (
      {stage1_61[84]},
      {stage2_61[60]}
   );
   gpc1_1 gpc3356 (
      {stage1_61[85]},
      {stage2_61[61]}
   );
   gpc1_1 gpc3357 (
      {stage1_61[86]},
      {stage2_61[62]}
   );
   gpc1_1 gpc3358 (
      {stage1_61[87]},
      {stage2_61[63]}
   );
   gpc1_1 gpc3359 (
      {stage1_61[88]},
      {stage2_61[64]}
   );
   gpc1_1 gpc3360 (
      {stage1_61[89]},
      {stage2_61[65]}
   );
   gpc1_1 gpc3361 (
      {stage1_61[90]},
      {stage2_61[66]}
   );
   gpc1_1 gpc3362 (
      {stage1_62[78]},
      {stage2_62[26]}
   );
   gpc1_1 gpc3363 (
      {stage1_62[79]},
      {stage2_62[27]}
   );
   gpc1_1 gpc3364 (
      {stage1_62[80]},
      {stage2_62[28]}
   );
   gpc1_1 gpc3365 (
      {stage1_62[81]},
      {stage2_62[29]}
   );
   gpc1_1 gpc3366 (
      {stage1_62[82]},
      {stage2_62[30]}
   );
   gpc1_1 gpc3367 (
      {stage1_62[83]},
      {stage2_62[31]}
   );
   gpc1_1 gpc3368 (
      {stage1_62[84]},
      {stage2_62[32]}
   );
   gpc1_1 gpc3369 (
      {stage1_62[85]},
      {stage2_62[33]}
   );
   gpc1_1 gpc3370 (
      {stage1_62[86]},
      {stage2_62[34]}
   );
   gpc1_1 gpc3371 (
      {stage1_63[48]},
      {stage2_63[23]}
   );
   gpc1_1 gpc3372 (
      {stage1_63[49]},
      {stage2_63[24]}
   );
   gpc1_1 gpc3373 (
      {stage1_63[50]},
      {stage2_63[25]}
   );
   gpc1_1 gpc3374 (
      {stage1_63[51]},
      {stage2_63[26]}
   );
   gpc1_1 gpc3375 (
      {stage1_63[52]},
      {stage2_63[27]}
   );
   gpc1_1 gpc3376 (
      {stage1_63[53]},
      {stage2_63[28]}
   );
   gpc1_1 gpc3377 (
      {stage1_63[54]},
      {stage2_63[29]}
   );
   gpc1_1 gpc3378 (
      {stage1_63[55]},
      {stage2_63[30]}
   );
   gpc1_1 gpc3379 (
      {stage1_63[56]},
      {stage2_63[31]}
   );
   gpc1_1 gpc3380 (
      {stage1_63[57]},
      {stage2_63[32]}
   );
   gpc1_1 gpc3381 (
      {stage1_63[58]},
      {stage2_63[33]}
   );
   gpc1_1 gpc3382 (
      {stage1_63[59]},
      {stage2_63[34]}
   );
   gpc1_1 gpc3383 (
      {stage1_63[60]},
      {stage2_63[35]}
   );
   gpc1_1 gpc3384 (
      {stage1_63[61]},
      {stage2_63[36]}
   );
   gpc1_1 gpc3385 (
      {stage1_63[62]},
      {stage2_63[37]}
   );
   gpc1_1 gpc3386 (
      {stage1_64[18]},
      {stage2_64[19]}
   );
   gpc1_1 gpc3387 (
      {stage1_64[19]},
      {stage2_64[20]}
   );
   gpc1_1 gpc3388 (
      {stage1_64[20]},
      {stage2_64[21]}
   );
   gpc1_1 gpc3389 (
      {stage1_64[21]},
      {stage2_64[22]}
   );
   gpc1_1 gpc3390 (
      {stage1_64[22]},
      {stage2_64[23]}
   );
   gpc1_1 gpc3391 (
      {stage1_64[23]},
      {stage2_64[24]}
   );
   gpc1_1 gpc3392 (
      {stage1_64[24]},
      {stage2_64[25]}
   );
   gpc1_1 gpc3393 (
      {stage1_64[25]},
      {stage2_64[26]}
   );
   gpc1_1 gpc3394 (
      {stage1_64[26]},
      {stage2_64[27]}
   );
   gpc1_1 gpc3395 (
      {stage1_64[27]},
      {stage2_64[28]}
   );
   gpc1_1 gpc3396 (
      {stage1_64[28]},
      {stage2_64[29]}
   );
   gpc1_1 gpc3397 (
      {stage1_64[29]},
      {stage2_64[30]}
   );
   gpc1_1 gpc3398 (
      {stage1_64[30]},
      {stage2_64[31]}
   );
   gpc1_1 gpc3399 (
      {stage1_64[31]},
      {stage2_64[32]}
   );
   gpc1_1 gpc3400 (
      {stage1_64[32]},
      {stage2_64[33]}
   );
   gpc1_1 gpc3401 (
      {stage1_64[33]},
      {stage2_64[34]}
   );
   gpc1_1 gpc3402 (
      {stage1_64[34]},
      {stage2_64[35]}
   );
   gpc1_1 gpc3403 (
      {stage1_64[35]},
      {stage2_64[36]}
   );
   gpc1_1 gpc3404 (
      {stage1_64[36]},
      {stage2_64[37]}
   );
   gpc1_1 gpc3405 (
      {stage1_64[37]},
      {stage2_64[38]}
   );
   gpc1_1 gpc3406 (
      {stage1_64[38]},
      {stage2_64[39]}
   );
   gpc1_1 gpc3407 (
      {stage1_64[39]},
      {stage2_64[40]}
   );
   gpc1_1 gpc3408 (
      {stage1_64[40]},
      {stage2_64[41]}
   );
   gpc1_1 gpc3409 (
      {stage1_64[41]},
      {stage2_64[42]}
   );
   gpc1_1 gpc3410 (
      {stage1_64[42]},
      {stage2_64[43]}
   );
   gpc1_1 gpc3411 (
      {stage1_64[43]},
      {stage2_64[44]}
   );
   gpc1_1 gpc3412 (
      {stage1_64[44]},
      {stage2_64[45]}
   );
   gpc1163_5 gpc3413 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3414 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc3415 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc3416 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[2],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc3417 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[1]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[3],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc3418 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[2]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[4],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc3419 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[3]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[5],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc3420 (
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[6],stage3_4[7],stage3_3[7]}
   );
   gpc615_5 gpc3421 (
      {stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[7],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc3422 (
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[8],stage3_4[9],stage3_3[9]}
   );
   gpc606_5 gpc3423 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[9],stage3_4[10]}
   );
   gpc606_5 gpc3424 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[10]}
   );
   gpc606_5 gpc3425 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[11]}
   );
   gpc606_5 gpc3426 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[3],stage3_7[6],stage3_6[12]}
   );
   gpc606_5 gpc3427 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[4],stage3_7[7],stage3_6[13]}
   );
   gpc606_5 gpc3428 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[5],stage3_7[8],stage3_6[14]}
   );
   gpc207_4 gpc3429 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[3],stage3_9[5],stage3_8[6],stage3_7[9]}
   );
   gpc207_4 gpc3430 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25]},
      {stage2_9[2], stage2_9[3]},
      {stage3_10[4],stage3_9[6],stage3_8[7],stage3_7[10]}
   );
   gpc606_5 gpc3431 (
      {stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9]},
      {stage3_11[0],stage3_10[5],stage3_9[7],stage3_8[8],stage3_7[11]}
   );
   gpc615_5 gpc3432 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[18]},
      {stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15]},
      {stage3_11[1],stage3_10[6],stage3_9[8],stage3_8[9],stage3_7[12]}
   );
   gpc606_5 gpc3433 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[7],stage3_9[9],stage3_8[10]}
   );
   gpc606_5 gpc3434 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[8],stage3_9[10],stage3_8[11]}
   );
   gpc606_5 gpc3435 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[4],stage3_10[9],stage3_9[11],stage3_8[12]}
   );
   gpc606_5 gpc3436 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[5],stage3_10[10],stage3_9[12],stage3_8[13]}
   );
   gpc606_5 gpc3437 (
      {stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[6],stage3_10[11],stage3_9[13],stage3_8[14]}
   );
   gpc606_5 gpc3438 (
      {stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[7],stage3_10[12],stage3_9[14],stage3_8[15]}
   );
   gpc606_5 gpc3439 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], 1'b0},
      {stage3_12[6],stage3_11[8],stage3_10[13],stage3_9[15],stage3_8[16]}
   );
   gpc606_5 gpc3440 (
      {stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[9],stage3_10[14],stage3_9[16]}
   );
   gpc606_5 gpc3441 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[8],stage3_11[10]}
   );
   gpc606_5 gpc3442 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[2],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc3443 (
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[3],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc3444 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[4],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc3445 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[5],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc3446 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[5],stage3_13[6],stage3_12[13]}
   );
   gpc606_5 gpc3447 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[6],stage3_14[6],stage3_13[7],stage3_12[14]}
   );
   gpc606_5 gpc3448 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[7],stage3_14[7],stage3_13[8],stage3_12[15]}
   );
   gpc606_5 gpc3449 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[8],stage3_14[8],stage3_13[9],stage3_12[16]}
   );
   gpc606_5 gpc3450 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[9],stage3_14[9],stage3_13[10]}
   );
   gpc615_5 gpc3451 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[10],stage3_14[10]}
   );
   gpc615_5 gpc3452 (
      {stage2_14[29], stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33]},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[11],stage3_14[11]}
   );
   gpc615_5 gpc3453 (
      {stage2_14[34], stage2_14[35], stage2_14[36], stage2_14[37], stage2_14[38]},
      {stage2_15[8]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[12],stage3_14[12]}
   );
   gpc615_5 gpc3454 (
      {stage2_14[39], stage2_14[40], stage2_14[41], stage2_14[42], stage2_14[43]},
      {stage2_15[9]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[13],stage3_14[13]}
   );
   gpc615_5 gpc3455 (
      {stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47], stage2_14[48]},
      {stage2_15[10]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[5],stage3_16[9],stage3_15[14],stage3_14[14]}
   );
   gpc615_5 gpc3456 (
      {stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage2_15[11]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[6],stage3_16[10],stage3_15[15],stage3_14[15]}
   );
   gpc615_5 gpc3457 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[7],stage3_16[11],stage3_15[16]}
   );
   gpc606_5 gpc3458 (
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[7],stage3_17[8]}
   );
   gpc606_5 gpc3459 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[2],stage3_18[8],stage3_17[9]}
   );
   gpc606_5 gpc3460 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[2],stage3_19[3],stage3_18[9],stage3_17[10]}
   );
   gpc606_5 gpc3461 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[3],stage3_19[4],stage3_18[10],stage3_17[11]}
   );
   gpc606_5 gpc3462 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[4],stage3_19[5],stage3_18[11],stage3_17[12]}
   );
   gpc615_5 gpc3463 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[30]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[5],stage3_20[5],stage3_19[6],stage3_18[12]}
   );
   gpc615_5 gpc3464 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[31]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[6],stage3_20[6],stage3_19[7],stage3_18[13]}
   );
   gpc615_5 gpc3465 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[32]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[7],stage3_20[7],stage3_19[8],stage3_18[14]}
   );
   gpc615_5 gpc3466 (
      {stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[33]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[8],stage3_20[8],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc3467 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[34]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[9],stage3_20[9],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc3468 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[35]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[10],stage3_20[10],stage3_19[11],stage3_18[17]}
   );
   gpc615_5 gpc3469 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[36]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[11],stage3_20[11],stage3_19[12],stage3_18[18]}
   );
   gpc615_5 gpc3470 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[37]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[12],stage3_20[12],stage3_19[13],stage3_18[19]}
   );
   gpc615_5 gpc3471 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[8],stage3_21[13]}
   );
   gpc615_5 gpc3472 (
      {stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[9],stage3_21[14]}
   );
   gpc615_5 gpc3473 (
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[10],stage3_21[15]}
   );
   gpc615_5 gpc3474 (
      {stage2_21[15], stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19]},
      {stage2_22[3]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[11],stage3_21[16]}
   );
   gpc615_5 gpc3475 (
      {stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[4]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[12],stage3_21[17]}
   );
   gpc615_5 gpc3476 (
      {stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage2_22[5]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[5],stage3_24[5],stage3_23[5],stage3_22[13],stage3_21[18]}
   );
   gpc615_5 gpc3477 (
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34]},
      {stage2_22[6]},
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage3_25[6],stage3_24[6],stage3_23[6],stage3_22[14],stage3_21[19]}
   );
   gpc615_5 gpc3478 (
      {stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_23[42]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[7],stage3_24[7],stage3_23[7],stage3_22[15]}
   );
   gpc615_5 gpc3479 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16]},
      {stage2_23[43]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[8],stage3_24[8],stage3_23[8],stage3_22[16]}
   );
   gpc615_5 gpc3480 (
      {stage2_22[17], stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[44]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[9],stage3_24[9],stage3_23[9],stage3_22[17]}
   );
   gpc615_5 gpc3481 (
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[3],stage3_25[10],stage3_24[10]}
   );
   gpc615_5 gpc3482 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_25[1]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[1],stage3_26[4],stage3_25[11],stage3_24[11]}
   );
   gpc615_5 gpc3483 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32]},
      {stage2_25[2]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[2],stage3_26[5],stage3_25[12],stage3_24[12]}
   );
   gpc606_5 gpc3484 (
      {stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[3],stage3_27[3],stage3_26[6],stage3_25[13]}
   );
   gpc606_5 gpc3485 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], stage2_25[13], stage2_25[14]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[4],stage3_27[4],stage3_26[7],stage3_25[14]}
   );
   gpc606_5 gpc3486 (
      {stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18], stage2_25[19], stage2_25[20]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[5],stage3_27[5],stage3_26[8],stage3_25[15]}
   );
   gpc606_5 gpc3487 (
      {stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24], stage2_25[25], stage2_25[26]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[6],stage3_27[6],stage3_26[9],stage3_25[16]}
   );
   gpc606_5 gpc3488 (
      {stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30], stage2_25[31], stage2_25[32]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[7],stage3_27[7],stage3_26[10],stage3_25[17]}
   );
   gpc207_4 gpc3489 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24]},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[5],stage3_28[8],stage3_27[8],stage3_26[11]}
   );
   gpc207_4 gpc3490 (
      {stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31]},
      {stage2_28[2], stage2_28[3]},
      {stage3_29[6],stage3_28[9],stage3_27[9],stage3_26[12]}
   );
   gpc207_4 gpc3491 (
      {stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[4], stage2_28[5]},
      {stage3_29[7],stage3_28[10],stage3_27[10],stage3_26[13]}
   );
   gpc207_4 gpc3492 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45]},
      {stage2_28[6], stage2_28[7]},
      {stage3_29[8],stage3_28[11],stage3_27[11],stage3_26[14]}
   );
   gpc207_4 gpc3493 (
      {stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_28[8], stage2_28[9]},
      {stage3_29[9],stage3_28[12],stage3_27[12],stage3_26[15]}
   );
   gpc606_5 gpc3494 (
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[10],stage3_28[13],stage3_27[13]}
   );
   gpc606_5 gpc3495 (
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[1],stage3_29[11],stage3_28[14],stage3_27[14]}
   );
   gpc615_5 gpc3496 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[10]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[2],stage3_29[12],stage3_28[15],stage3_27[15]}
   );
   gpc606_5 gpc3497 (
      {stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[3],stage3_29[13],stage3_28[16]}
   );
   gpc606_5 gpc3498 (
      {stage2_28[17], stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[4],stage3_29[14],stage3_28[17]}
   );
   gpc606_5 gpc3499 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[5],stage3_29[15],stage3_28[18]}
   );
   gpc606_5 gpc3500 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[6],stage3_29[16],stage3_28[19]}
   );
   gpc606_5 gpc3501 (
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[4],stage3_31[7],stage3_30[7],stage3_29[17]}
   );
   gpc606_5 gpc3502 (
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[5],stage3_31[8],stage3_30[8],stage3_29[18]}
   );
   gpc606_5 gpc3503 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[6],stage3_31[9],stage3_30[9],stage3_29[19]}
   );
   gpc606_5 gpc3504 (
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[7],stage3_31[10],stage3_30[10],stage3_29[20]}
   );
   gpc606_5 gpc3505 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[8],stage3_31[11],stage3_30[11],stage3_29[21]}
   );
   gpc615_5 gpc3506 (
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28]},
      {stage2_31[30]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[5],stage3_32[9],stage3_31[12],stage3_30[12]}
   );
   gpc615_5 gpc3507 (
      {stage2_30[29], stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33]},
      {stage2_31[31]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[6],stage3_32[10],stage3_31[13],stage3_30[13]}
   );
   gpc615_5 gpc3508 (
      {stage2_30[34], stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38]},
      {stage2_31[32]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[7],stage3_32[11],stage3_31[14],stage3_30[14]}
   );
   gpc606_5 gpc3509 (
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[0],stage3_34[3],stage3_33[8],stage3_32[12]}
   );
   gpc606_5 gpc3510 (
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[1],stage3_34[4],stage3_33[9],stage3_32[13]}
   );
   gpc606_5 gpc3511 (
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[2],stage3_34[5],stage3_33[10],stage3_32[14]}
   );
   gpc7_3 gpc3512 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[3],stage3_34[6],stage3_33[11]}
   );
   gpc7_3 gpc3513 (
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12], stage2_33[13]},
      {stage3_35[4],stage3_34[7],stage3_33[12]}
   );
   gpc7_3 gpc3514 (
      {stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18], stage2_33[19], stage2_33[20]},
      {stage3_35[5],stage3_34[8],stage3_33[13]}
   );
   gpc7_3 gpc3515 (
      {stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27]},
      {stage3_35[6],stage3_34[9],stage3_33[14]}
   );
   gpc615_5 gpc3516 (
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22]},
      {stage2_35[0]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[3],stage3_35[7],stage3_34[10]}
   );
   gpc606_5 gpc3517 (
      {stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5], stage2_35[6]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[1],stage3_37[1],stage3_36[4],stage3_35[8]}
   );
   gpc606_5 gpc3518 (
      {stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[2],stage3_37[2],stage3_36[5],stage3_35[9]}
   );
   gpc615_5 gpc3519 (
      {stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage2_36[6]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[3],stage3_37[3],stage3_36[6],stage3_35[10]}
   );
   gpc615_5 gpc3520 (
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22]},
      {stage2_36[7]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[4],stage3_37[4],stage3_36[7],stage3_35[11]}
   );
   gpc615_5 gpc3521 (
      {stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_36[8]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[5],stage3_37[5],stage3_36[8],stage3_35[12]}
   );
   gpc615_5 gpc3522 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[9]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[6],stage3_37[6],stage3_36[9],stage3_35[13]}
   );
   gpc606_5 gpc3523 (
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[6],stage3_38[7],stage3_37[7],stage3_36[10]}
   );
   gpc606_5 gpc3524 (
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage3_40[1],stage3_39[7],stage3_38[8],stage3_37[8],stage3_36[11]}
   );
   gpc606_5 gpc3525 (
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage3_40[2],stage3_39[8],stage3_38[9],stage3_37[9],stage3_36[12]}
   );
   gpc606_5 gpc3526 (
      {stage2_36[28], stage2_36[29], stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33]},
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage3_40[3],stage3_39[9],stage3_38[10],stage3_37[10],stage3_36[13]}
   );
   gpc606_5 gpc3527 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[4],stage3_39[10],stage3_38[11],stage3_37[11]}
   );
   gpc615_5 gpc3528 (
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28]},
      {stage2_39[6]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[1],stage3_40[5],stage3_39[11],stage3_38[12]}
   );
   gpc615_5 gpc3529 (
      {stage2_38[29], stage2_38[30], stage2_38[31], stage2_38[32], 1'b0},
      {stage2_39[7]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[2],stage3_40[6],stage3_39[12],stage3_38[13]}
   );
   gpc606_5 gpc3530 (
      {stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11], stage2_39[12], stage2_39[13]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[2],stage3_41[3],stage3_40[7],stage3_39[13]}
   );
   gpc606_5 gpc3531 (
      {stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[3],stage3_41[4],stage3_40[8],stage3_39[14]}
   );
   gpc606_5 gpc3532 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24], stage2_39[25]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[4],stage3_41[5],stage3_40[9],stage3_39[15]}
   );
   gpc606_5 gpc3533 (
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[3],stage3_42[5],stage3_41[6],stage3_40[10]}
   );
   gpc606_5 gpc3534 (
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[4],stage3_42[6],stage3_41[7],stage3_40[11]}
   );
   gpc606_5 gpc3535 (
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[5],stage3_42[7],stage3_41[8],stage3_40[12]}
   );
   gpc606_5 gpc3536 (
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[3],stage3_43[6],stage3_42[8],stage3_41[9]}
   );
   gpc606_5 gpc3537 (
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11]},
      {stage3_45[1],stage3_44[4],stage3_43[7],stage3_42[9],stage3_41[10]}
   );
   gpc615_5 gpc3538 (
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34]},
      {stage2_42[18]},
      {stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17]},
      {stage3_45[2],stage3_44[5],stage3_43[8],stage3_42[10],stage3_41[11]}
   );
   gpc615_5 gpc3539 (
      {stage2_41[35], stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39]},
      {stage2_42[19]},
      {stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage3_45[3],stage3_44[6],stage3_43[9],stage3_42[11],stage3_41[12]}
   );
   gpc615_5 gpc3540 (
      {stage2_41[40], stage2_41[41], stage2_41[42], stage2_41[43], stage2_41[44]},
      {stage2_42[20]},
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28], stage2_43[29]},
      {stage3_45[4],stage3_44[7],stage3_43[10],stage3_42[12],stage3_41[13]}
   );
   gpc615_5 gpc3541 (
      {stage2_42[21], stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25]},
      {stage2_43[30]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[5],stage3_44[8],stage3_43[11],stage3_42[13]}
   );
   gpc615_5 gpc3542 (
      {stage2_42[26], stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30]},
      {stage2_43[31]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[6],stage3_44[9],stage3_43[12],stage3_42[14]}
   );
   gpc615_5 gpc3543 (
      {stage2_42[31], stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35]},
      {stage2_43[32]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[7],stage3_44[10],stage3_43[13],stage3_42[15]}
   );
   gpc615_5 gpc3544 (
      {stage2_42[36], stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40]},
      {stage2_43[33]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[8],stage3_44[11],stage3_43[14],stage3_42[16]}
   );
   gpc615_5 gpc3545 (
      {stage2_42[41], stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45]},
      {stage2_43[34]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[9],stage3_44[12],stage3_43[15],stage3_42[17]}
   );
   gpc615_5 gpc3546 (
      {stage2_42[46], stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50]},
      {stage2_43[35]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[10],stage3_44[13],stage3_43[16],stage3_42[18]}
   );
   gpc615_5 gpc3547 (
      {stage2_42[51], stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55]},
      {stage2_43[36]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[11],stage3_44[14],stage3_43[17],stage3_42[19]}
   );
   gpc615_5 gpc3548 (
      {stage2_43[37], stage2_43[38], stage2_43[39], stage2_43[40], stage2_43[41]},
      {stage2_44[42]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[7],stage3_45[12],stage3_44[15],stage3_43[18]}
   );
   gpc615_5 gpc3549 (
      {stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45], stage2_43[46]},
      {stage2_44[43]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[8],stage3_45[13],stage3_44[16],stage3_43[19]}
   );
   gpc615_5 gpc3550 (
      {stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_44[44]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[9],stage3_45[14],stage3_44[17],stage3_43[20]}
   );
   gpc615_5 gpc3551 (
      {stage2_44[45], stage2_44[46], stage2_44[47], stage2_44[48], stage2_44[49]},
      {stage2_45[18]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[3],stage3_46[10],stage3_45[15],stage3_44[18]}
   );
   gpc615_5 gpc3552 (
      {stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53], stage2_44[54]},
      {stage2_45[19]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[4],stage3_46[11],stage3_45[16],stage3_44[19]}
   );
   gpc606_5 gpc3553 (
      {stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23], stage2_45[24], stage2_45[25]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[5],stage3_46[12],stage3_45[17]}
   );
   gpc606_5 gpc3554 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[1],stage3_48[3],stage3_47[6],stage3_46[13]}
   );
   gpc1325_5 gpc3555 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[6], stage2_47[7]},
      {stage2_48[6], stage2_48[7], stage2_48[8]},
      {stage2_49[0]},
      {stage3_50[1],stage3_49[2],stage3_48[4],stage3_47[7],stage3_46[14]}
   );
   gpc1325_5 gpc3556 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[8], stage2_47[9]},
      {stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage2_49[1]},
      {stage3_50[2],stage3_49[3],stage3_48[5],stage3_47[8],stage3_46[15]}
   );
   gpc1325_5 gpc3557 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[10], stage2_47[11]},
      {stage2_48[12], stage2_48[13], stage2_48[14]},
      {stage2_49[2]},
      {stage3_50[3],stage3_49[4],stage3_48[6],stage3_47[9],stage3_46[16]}
   );
   gpc615_5 gpc3558 (
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16]},
      {stage2_48[15]},
      {stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7], stage2_49[8]},
      {stage3_51[0],stage3_50[4],stage3_49[5],stage3_48[7],stage3_47[10]}
   );
   gpc615_5 gpc3559 (
      {stage2_47[17], stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21]},
      {stage2_48[16]},
      {stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13], stage2_49[14]},
      {stage3_51[1],stage3_50[5],stage3_49[6],stage3_48[8],stage3_47[11]}
   );
   gpc615_5 gpc3560 (
      {stage2_47[22], stage2_47[23], stage2_47[24], stage2_47[25], stage2_47[26]},
      {stage2_48[17]},
      {stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19], stage2_49[20]},
      {stage3_51[2],stage3_50[6],stage3_49[7],stage3_48[9],stage3_47[12]}
   );
   gpc615_5 gpc3561 (
      {stage2_47[27], stage2_47[28], stage2_47[29], stage2_47[30], stage2_47[31]},
      {stage2_48[18]},
      {stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25], stage2_49[26]},
      {stage3_51[3],stage3_50[7],stage3_49[8],stage3_48[10],stage3_47[13]}
   );
   gpc615_5 gpc3562 (
      {stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35], stage2_47[36]},
      {stage2_48[19]},
      {stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31], stage2_49[32]},
      {stage3_51[4],stage3_50[8],stage3_49[9],stage3_48[11],stage3_47[14]}
   );
   gpc2116_5 gpc3563 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[0],stage3_52[0],stage3_51[5],stage3_50[9]}
   );
   gpc2116_5 gpc3564 (
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage2_51[1]},
      {stage2_52[1]},
      {stage2_53[2], stage2_53[3]},
      {stage3_54[1],stage3_53[1],stage3_52[1],stage3_51[6],stage3_50[10]}
   );
   gpc615_5 gpc3565 (
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16]},
      {stage2_51[2]},
      {stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5], stage2_52[6], stage2_52[7]},
      {stage3_54[2],stage3_53[2],stage3_52[2],stage3_51[7],stage3_50[11]}
   );
   gpc615_5 gpc3566 (
      {stage2_50[17], stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21]},
      {stage2_51[3]},
      {stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12], stage2_52[13]},
      {stage3_54[3],stage3_53[3],stage3_52[3],stage3_51[8],stage3_50[12]}
   );
   gpc615_5 gpc3567 (
      {stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7], stage2_51[8]},
      {stage2_52[14]},
      {stage2_53[4], stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9]},
      {stage3_55[0],stage3_54[4],stage3_53[4],stage3_52[4],stage3_51[9]}
   );
   gpc615_5 gpc3568 (
      {stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12], stage2_51[13]},
      {stage2_52[15]},
      {stage2_53[10], stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15]},
      {stage3_55[1],stage3_54[5],stage3_53[5],stage3_52[5],stage3_51[10]}
   );
   gpc615_5 gpc3569 (
      {stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17], stage2_51[18]},
      {stage2_52[16]},
      {stage2_53[16], stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21]},
      {stage3_55[2],stage3_54[6],stage3_53[6],stage3_52[6],stage3_51[11]}
   );
   gpc615_5 gpc3570 (
      {stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage2_52[17]},
      {stage2_53[22], stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27]},
      {stage3_55[3],stage3_54[7],stage3_53[7],stage3_52[7],stage3_51[12]}
   );
   gpc606_5 gpc3571 (
      {stage2_53[28], stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[4],stage3_54[8],stage3_53[8]}
   );
   gpc606_5 gpc3572 (
      {stage2_53[34], stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[5],stage3_54[9],stage3_53[9]}
   );
   gpc606_5 gpc3573 (
      {stage2_53[40], stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[6],stage3_54[10],stage3_53[10]}
   );
   gpc606_5 gpc3574 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[3],stage3_56[3],stage3_55[7],stage3_54[11]}
   );
   gpc606_5 gpc3575 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[4],stage3_56[4],stage3_55[8],stage3_54[12]}
   );
   gpc606_5 gpc3576 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[5],stage3_56[5],stage3_55[9],stage3_54[13]}
   );
   gpc615_5 gpc3577 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22]},
      {stage2_55[18]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[6],stage3_56[6],stage3_55[10],stage3_54[14]}
   );
   gpc615_5 gpc3578 (
      {stage2_54[23], stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27]},
      {stage2_55[19]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[7],stage3_56[7],stage3_55[11],stage3_54[15]}
   );
   gpc615_5 gpc3579 (
      {stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23], stage2_55[24]},
      {stage2_56[30]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[5],stage3_57[8],stage3_56[8],stage3_55[12]}
   );
   gpc615_5 gpc3580 (
      {stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage2_56[31]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[6],stage3_57[9],stage3_56[9],stage3_55[13]}
   );
   gpc615_5 gpc3581 (
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34]},
      {stage2_56[32]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[7],stage3_57[10],stage3_56[10],stage3_55[14]}
   );
   gpc606_5 gpc3582 (
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[0],stage3_59[3],stage3_58[8],stage3_57[11]}
   );
   gpc606_5 gpc3583 (
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[1],stage3_59[4],stage3_58[9],stage3_57[12]}
   );
   gpc1163_5 gpc3584 (
      {stage2_58[0], stage2_58[1], stage2_58[2]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage2_60[0]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[2],stage3_60[2],stage3_59[5],stage3_58[10]}
   );
   gpc615_5 gpc3585 (
      {stage2_58[3], stage2_58[4], stage2_58[5], stage2_58[6], stage2_58[7]},
      {stage2_59[18]},
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage3_62[1],stage3_61[3],stage3_60[3],stage3_59[6],stage3_58[11]}
   );
   gpc615_5 gpc3586 (
      {stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11], stage2_58[12]},
      {stage2_59[19]},
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage3_62[2],stage3_61[4],stage3_60[4],stage3_59[7],stage3_58[12]}
   );
   gpc135_4 gpc3587 (
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24]},
      {stage2_60[13], stage2_60[14], stage2_60[15]},
      {stage2_61[1]},
      {stage3_62[3],stage3_61[5],stage3_60[5],stage3_59[8]}
   );
   gpc606_5 gpc3588 (
      {stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30]},
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6], stage2_61[7]},
      {stage3_63[0],stage3_62[4],stage3_61[6],stage3_60[6],stage3_59[9]}
   );
   gpc606_5 gpc3589 (
      {stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36]},
      {stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12], stage2_61[13]},
      {stage3_63[1],stage3_62[5],stage3_61[7],stage3_60[7],stage3_59[10]}
   );
   gpc606_5 gpc3590 (
      {stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42]},
      {stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17], stage2_61[18], stage2_61[19]},
      {stage3_63[2],stage3_62[6],stage3_61[8],stage3_60[8],stage3_59[11]}
   );
   gpc606_5 gpc3591 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23], stage2_61[24], stage2_61[25]},
      {stage3_63[3],stage3_62[7],stage3_61[9],stage3_60[9],stage3_59[12]}
   );
   gpc606_5 gpc3592 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29], stage2_61[30], stage2_61[31]},
      {stage3_63[4],stage3_62[8],stage3_61[10],stage3_60[10],stage3_59[13]}
   );
   gpc615_5 gpc3593 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[16]},
      {stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35], stage2_61[36], stage2_61[37]},
      {stage3_63[5],stage3_62[9],stage3_61[11],stage3_60[11],stage3_59[14]}
   );
   gpc615_5 gpc3594 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[17]},
      {stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41], stage2_61[42], stage2_61[43]},
      {stage3_63[6],stage3_62[10],stage3_61[12],stage3_60[12],stage3_59[15]}
   );
   gpc615_5 gpc3595 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[18]},
      {stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47], stage2_61[48], stage2_61[49]},
      {stage3_63[7],stage3_62[11],stage3_61[13],stage3_60[13],stage3_59[16]}
   );
   gpc606_5 gpc3596 (
      {stage2_60[19], stage2_60[20], stage2_60[21], 1'b0, 1'b0, 1'b0},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[8],stage3_62[12],stage3_61[14],stage3_60[14]}
   );
   gpc1163_5 gpc3597 (
      {stage2_61[50], stage2_61[51], stage2_61[52]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_63[0]},
      {stage2_64[0]},
      {stage3_65[0],stage3_64[1],stage3_63[9],stage3_62[13],stage3_61[15]}
   );
   gpc606_5 gpc3598 (
      {stage2_61[53], stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58]},
      {stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage3_65[1],stage3_64[2],stage3_63[10],stage3_62[14],stage3_61[16]}
   );
   gpc1163_5 gpc3599 (
      {stage2_62[12], stage2_62[13], stage2_62[14]},
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12]},
      {stage2_64[1]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[2],stage3_64[3],stage3_63[11],stage3_62[15]}
   );
   gpc1163_5 gpc3600 (
      {stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18]},
      {stage2_64[2]},
      {stage2_65[1]},
      {stage3_66[1],stage3_65[3],stage3_64[4],stage3_63[12],stage3_62[16]}
   );
   gpc1163_5 gpc3601 (
      {stage2_62[18], stage2_62[19], stage2_62[20]},
      {stage2_63[19], stage2_63[20], stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24]},
      {stage2_64[3]},
      {stage2_65[2]},
      {stage3_66[2],stage3_65[4],stage3_64[5],stage3_63[13],stage3_62[17]}
   );
   gpc1163_5 gpc3602 (
      {stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage2_63[25], stage2_63[26], stage2_63[27], stage2_63[28], stage2_63[29], stage2_63[30]},
      {stage2_64[4]},
      {stage2_65[3]},
      {stage3_66[3],stage3_65[5],stage3_64[6],stage3_63[14],stage3_62[18]}
   );
   gpc606_5 gpc3603 (
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage2_64[5], stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10]},
      {stage3_66[4],stage3_65[6],stage3_64[7],stage3_63[15],stage3_62[19]}
   );
   gpc615_5 gpc3604 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[31]},
      {stage2_64[11], stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16]},
      {stage3_66[5],stage3_65[7],stage3_64[8],stage3_63[16],stage3_62[20]}
   );
   gpc606_5 gpc3605 (
      {stage2_63[32], stage2_63[33], stage2_63[34], stage2_63[35], stage2_63[36], stage2_63[37]},
      {stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9]},
      {stage3_67[0],stage3_66[6],stage3_65[8],stage3_64[9],stage3_63[17]}
   );
   gpc606_5 gpc3606 (
      {stage2_64[17], stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[1],stage3_66[7],stage3_65[9],stage3_64[10]}
   );
   gpc606_5 gpc3607 (
      {stage2_64[23], stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], 1'b0, 1'b0},
      {stage3_68[1],stage3_67[2],stage3_66[8],stage3_65[10],stage3_64[11]}
   );
   gpc1_1 gpc3608 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc3609 (
      {stage2_0[4]},
      {stage3_0[2]}
   );
   gpc1_1 gpc3610 (
      {stage2_0[5]},
      {stage3_0[3]}
   );
   gpc1_1 gpc3611 (
      {stage2_0[6]},
      {stage3_0[4]}
   );
   gpc1_1 gpc3612 (
      {stage2_0[7]},
      {stage3_0[5]}
   );
   gpc1_1 gpc3613 (
      {stage2_0[8]},
      {stage3_0[6]}
   );
   gpc1_1 gpc3614 (
      {stage2_0[9]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3615 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc3616 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc3617 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc3618 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc3619 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc3620 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc3621 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc3622 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc3623 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc3624 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc3625 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc3626 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc3627 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc3628 (
      {stage2_2[34]},
      {stage3_2[7]}
   );
   gpc1_1 gpc3629 (
      {stage2_2[35]},
      {stage3_2[8]}
   );
   gpc1_1 gpc3630 (
      {stage2_2[36]},
      {stage3_2[9]}
   );
   gpc1_1 gpc3631 (
      {stage2_2[37]},
      {stage3_2[10]}
   );
   gpc1_1 gpc3632 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc3633 (
      {stage2_3[20]},
      {stage3_3[11]}
   );
   gpc1_1 gpc3634 (
      {stage2_3[21]},
      {stage3_3[12]}
   );
   gpc1_1 gpc3635 (
      {stage2_3[22]},
      {stage3_3[13]}
   );
   gpc1_1 gpc3636 (
      {stage2_4[45]},
      {stage3_4[11]}
   );
   gpc1_1 gpc3637 (
      {stage2_4[46]},
      {stage3_4[12]}
   );
   gpc1_1 gpc3638 (
      {stage2_4[47]},
      {stage3_4[13]}
   );
   gpc1_1 gpc3639 (
      {stage2_5[30]},
      {stage3_5[12]}
   );
   gpc1_1 gpc3640 (
      {stage2_5[31]},
      {stage3_5[13]}
   );
   gpc1_1 gpc3641 (
      {stage2_5[32]},
      {stage3_5[14]}
   );
   gpc1_1 gpc3642 (
      {stage2_5[33]},
      {stage3_5[15]}
   );
   gpc1_1 gpc3643 (
      {stage2_5[34]},
      {stage3_5[16]}
   );
   gpc1_1 gpc3644 (
      {stage2_5[35]},
      {stage3_5[17]}
   );
   gpc1_1 gpc3645 (
      {stage2_6[24]},
      {stage3_6[15]}
   );
   gpc1_1 gpc3646 (
      {stage2_6[25]},
      {stage3_6[16]}
   );
   gpc1_1 gpc3647 (
      {stage2_6[26]},
      {stage3_6[17]}
   );
   gpc1_1 gpc3648 (
      {stage2_6[27]},
      {stage3_6[18]}
   );
   gpc1_1 gpc3649 (
      {stage2_6[28]},
      {stage3_6[19]}
   );
   gpc1_1 gpc3650 (
      {stage2_7[37]},
      {stage3_7[13]}
   );
   gpc1_1 gpc3651 (
      {stage2_7[38]},
      {stage3_7[14]}
   );
   gpc1_1 gpc3652 (
      {stage2_7[39]},
      {stage3_7[15]}
   );
   gpc1_1 gpc3653 (
      {stage2_7[40]},
      {stage3_7[16]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[22]},
      {stage3_9[17]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[23]},
      {stage3_9[18]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[24]},
      {stage3_9[19]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[25]},
      {stage3_9[20]}
   );
   gpc1_1 gpc3658 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc3659 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc3660 (
      {stage2_11[38]},
      {stage3_11[17]}
   );
   gpc1_1 gpc3661 (
      {stage2_12[24]},
      {stage3_12[17]}
   );
   gpc1_1 gpc3662 (
      {stage2_12[25]},
      {stage3_12[18]}
   );
   gpc1_1 gpc3663 (
      {stage2_12[26]},
      {stage3_12[19]}
   );
   gpc1_1 gpc3664 (
      {stage2_12[27]},
      {stage3_12[20]}
   );
   gpc1_1 gpc3665 (
      {stage2_12[28]},
      {stage3_12[21]}
   );
   gpc1_1 gpc3666 (
      {stage2_12[29]},
      {stage3_12[22]}
   );
   gpc1_1 gpc3667 (
      {stage2_12[30]},
      {stage3_12[23]}
   );
   gpc1_1 gpc3668 (
      {stage2_13[36]},
      {stage3_13[11]}
   );
   gpc1_1 gpc3669 (
      {stage2_13[37]},
      {stage3_13[12]}
   );
   gpc1_1 gpc3670 (
      {stage2_13[38]},
      {stage3_13[13]}
   );
   gpc1_1 gpc3671 (
      {stage2_13[39]},
      {stage3_13[14]}
   );
   gpc1_1 gpc3672 (
      {stage2_13[40]},
      {stage3_13[15]}
   );
   gpc1_1 gpc3673 (
      {stage2_13[41]},
      {stage3_13[16]}
   );
   gpc1_1 gpc3674 (
      {stage2_13[42]},
      {stage3_13[17]}
   );
   gpc1_1 gpc3675 (
      {stage2_13[43]},
      {stage3_13[18]}
   );
   gpc1_1 gpc3676 (
      {stage2_13[44]},
      {stage3_13[19]}
   );
   gpc1_1 gpc3677 (
      {stage2_14[54]},
      {stage3_14[16]}
   );
   gpc1_1 gpc3678 (
      {stage2_14[55]},
      {stage3_14[17]}
   );
   gpc1_1 gpc3679 (
      {stage2_14[56]},
      {stage3_14[18]}
   );
   gpc1_1 gpc3680 (
      {stage2_14[57]},
      {stage3_14[19]}
   );
   gpc1_1 gpc3681 (
      {stage2_14[58]},
      {stage3_14[20]}
   );
   gpc1_1 gpc3682 (
      {stage2_14[59]},
      {stage3_14[21]}
   );
   gpc1_1 gpc3683 (
      {stage2_14[60]},
      {stage3_14[22]}
   );
   gpc1_1 gpc3684 (
      {stage2_14[61]},
      {stage3_14[23]}
   );
   gpc1_1 gpc3685 (
      {stage2_14[62]},
      {stage3_14[24]}
   );
   gpc1_1 gpc3686 (
      {stage2_14[63]},
      {stage3_14[25]}
   );
   gpc1_1 gpc3687 (
      {stage2_14[64]},
      {stage3_14[26]}
   );
   gpc1_1 gpc3688 (
      {stage2_14[65]},
      {stage3_14[27]}
   );
   gpc1_1 gpc3689 (
      {stage2_14[66]},
      {stage3_14[28]}
   );
   gpc1_1 gpc3690 (
      {stage2_14[67]},
      {stage3_14[29]}
   );
   gpc1_1 gpc3691 (
      {stage2_14[68]},
      {stage3_14[30]}
   );
   gpc1_1 gpc3692 (
      {stage2_14[69]},
      {stage3_14[31]}
   );
   gpc1_1 gpc3693 (
      {stage2_14[70]},
      {stage3_14[32]}
   );
   gpc1_1 gpc3694 (
      {stage2_14[71]},
      {stage3_14[33]}
   );
   gpc1_1 gpc3695 (
      {stage2_14[72]},
      {stage3_14[34]}
   );
   gpc1_1 gpc3696 (
      {stage2_14[73]},
      {stage3_14[35]}
   );
   gpc1_1 gpc3697 (
      {stage2_15[17]},
      {stage3_15[17]}
   );
   gpc1_1 gpc3698 (
      {stage2_15[18]},
      {stage3_15[18]}
   );
   gpc1_1 gpc3699 (
      {stage2_15[19]},
      {stage3_15[19]}
   );
   gpc1_1 gpc3700 (
      {stage2_15[20]},
      {stage3_15[20]}
   );
   gpc1_1 gpc3701 (
      {stage2_15[21]},
      {stage3_15[21]}
   );
   gpc1_1 gpc3702 (
      {stage2_15[22]},
      {stage3_15[22]}
   );
   gpc1_1 gpc3703 (
      {stage2_15[23]},
      {stage3_15[23]}
   );
   gpc1_1 gpc3704 (
      {stage2_15[24]},
      {stage3_15[24]}
   );
   gpc1_1 gpc3705 (
      {stage2_15[25]},
      {stage3_15[25]}
   );
   gpc1_1 gpc3706 (
      {stage2_15[26]},
      {stage3_15[26]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[27]},
      {stage3_15[27]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[28]},
      {stage3_15[28]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[29]},
      {stage3_15[29]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[30]},
      {stage3_15[30]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[31]},
      {stage3_15[31]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[32]},
      {stage3_15[32]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[33]},
      {stage3_15[33]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[34]},
      {stage3_15[34]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[35]},
      {stage3_15[35]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[36]},
      {stage3_15[36]}
   );
   gpc1_1 gpc3717 (
      {stage2_16[37]},
      {stage3_16[12]}
   );
   gpc1_1 gpc3718 (
      {stage2_16[38]},
      {stage3_16[13]}
   );
   gpc1_1 gpc3719 (
      {stage2_16[39]},
      {stage3_16[14]}
   );
   gpc1_1 gpc3720 (
      {stage2_16[40]},
      {stage3_16[15]}
   );
   gpc1_1 gpc3721 (
      {stage2_16[41]},
      {stage3_16[16]}
   );
   gpc1_1 gpc3722 (
      {stage2_16[42]},
      {stage3_16[17]}
   );
   gpc1_1 gpc3723 (
      {stage2_16[43]},
      {stage3_16[18]}
   );
   gpc1_1 gpc3724 (
      {stage2_16[44]},
      {stage3_16[19]}
   );
   gpc1_1 gpc3725 (
      {stage2_16[45]},
      {stage3_16[20]}
   );
   gpc1_1 gpc3726 (
      {stage2_16[46]},
      {stage3_16[21]}
   );
   gpc1_1 gpc3727 (
      {stage2_17[36]},
      {stage3_17[13]}
   );
   gpc1_1 gpc3728 (
      {stage2_17[37]},
      {stage3_17[14]}
   );
   gpc1_1 gpc3729 (
      {stage2_17[38]},
      {stage3_17[15]}
   );
   gpc1_1 gpc3730 (
      {stage2_17[39]},
      {stage3_17[16]}
   );
   gpc1_1 gpc3731 (
      {stage2_18[40]},
      {stage3_18[20]}
   );
   gpc1_1 gpc3732 (
      {stage2_18[41]},
      {stage3_18[21]}
   );
   gpc1_1 gpc3733 (
      {stage2_18[42]},
      {stage3_18[22]}
   );
   gpc1_1 gpc3734 (
      {stage2_19[38]},
      {stage3_19[14]}
   );
   gpc1_1 gpc3735 (
      {stage2_19[39]},
      {stage3_19[15]}
   );
   gpc1_1 gpc3736 (
      {stage2_19[40]},
      {stage3_19[16]}
   );
   gpc1_1 gpc3737 (
      {stage2_19[41]},
      {stage3_19[17]}
   );
   gpc1_1 gpc3738 (
      {stage2_19[42]},
      {stage3_19[18]}
   );
   gpc1_1 gpc3739 (
      {stage2_19[43]},
      {stage3_19[19]}
   );
   gpc1_1 gpc3740 (
      {stage2_19[44]},
      {stage3_19[20]}
   );
   gpc1_1 gpc3741 (
      {stage2_19[45]},
      {stage3_19[21]}
   );
   gpc1_1 gpc3742 (
      {stage2_19[46]},
      {stage3_19[22]}
   );
   gpc1_1 gpc3743 (
      {stage2_19[47]},
      {stage3_19[23]}
   );
   gpc1_1 gpc3744 (
      {stage2_19[48]},
      {stage3_19[24]}
   );
   gpc1_1 gpc3745 (
      {stage2_19[49]},
      {stage3_19[25]}
   );
   gpc1_1 gpc3746 (
      {stage2_19[50]},
      {stage3_19[26]}
   );
   gpc1_1 gpc3747 (
      {stage2_20[48]},
      {stage3_20[13]}
   );
   gpc1_1 gpc3748 (
      {stage2_20[49]},
      {stage3_20[14]}
   );
   gpc1_1 gpc3749 (
      {stage2_20[50]},
      {stage3_20[15]}
   );
   gpc1_1 gpc3750 (
      {stage2_20[51]},
      {stage3_20[16]}
   );
   gpc1_1 gpc3751 (
      {stage2_20[52]},
      {stage3_20[17]}
   );
   gpc1_1 gpc3752 (
      {stage2_20[53]},
      {stage3_20[18]}
   );
   gpc1_1 gpc3753 (
      {stage2_20[54]},
      {stage3_20[19]}
   );
   gpc1_1 gpc3754 (
      {stage2_20[55]},
      {stage3_20[20]}
   );
   gpc1_1 gpc3755 (
      {stage2_20[56]},
      {stage3_20[21]}
   );
   gpc1_1 gpc3756 (
      {stage2_20[57]},
      {stage3_20[22]}
   );
   gpc1_1 gpc3757 (
      {stage2_21[35]},
      {stage3_21[20]}
   );
   gpc1_1 gpc3758 (
      {stage2_21[36]},
      {stage3_21[21]}
   );
   gpc1_1 gpc3759 (
      {stage2_21[37]},
      {stage3_21[22]}
   );
   gpc1_1 gpc3760 (
      {stage2_21[38]},
      {stage3_21[23]}
   );
   gpc1_1 gpc3761 (
      {stage2_21[39]},
      {stage3_21[24]}
   );
   gpc1_1 gpc3762 (
      {stage2_22[22]},
      {stage3_22[18]}
   );
   gpc1_1 gpc3763 (
      {stage2_22[23]},
      {stage3_22[19]}
   );
   gpc1_1 gpc3764 (
      {stage2_22[24]},
      {stage3_22[20]}
   );
   gpc1_1 gpc3765 (
      {stage2_22[25]},
      {stage3_22[21]}
   );
   gpc1_1 gpc3766 (
      {stage2_22[26]},
      {stage3_22[22]}
   );
   gpc1_1 gpc3767 (
      {stage2_22[27]},
      {stage3_22[23]}
   );
   gpc1_1 gpc3768 (
      {stage2_22[28]},
      {stage3_22[24]}
   );
   gpc1_1 gpc3769 (
      {stage2_22[29]},
      {stage3_22[25]}
   );
   gpc1_1 gpc3770 (
      {stage2_22[30]},
      {stage3_22[26]}
   );
   gpc1_1 gpc3771 (
      {stage2_23[45]},
      {stage3_23[10]}
   );
   gpc1_1 gpc3772 (
      {stage2_23[46]},
      {stage3_23[11]}
   );
   gpc1_1 gpc3773 (
      {stage2_24[33]},
      {stage3_24[13]}
   );
   gpc1_1 gpc3774 (
      {stage2_24[34]},
      {stage3_24[14]}
   );
   gpc1_1 gpc3775 (
      {stage2_24[35]},
      {stage3_24[15]}
   );
   gpc1_1 gpc3776 (
      {stage2_24[36]},
      {stage3_24[16]}
   );
   gpc1_1 gpc3777 (
      {stage2_24[37]},
      {stage3_24[17]}
   );
   gpc1_1 gpc3778 (
      {stage2_24[38]},
      {stage3_24[18]}
   );
   gpc1_1 gpc3779 (
      {stage2_24[39]},
      {stage3_24[19]}
   );
   gpc1_1 gpc3780 (
      {stage2_24[40]},
      {stage3_24[20]}
   );
   gpc1_1 gpc3781 (
      {stage2_24[41]},
      {stage3_24[21]}
   );
   gpc1_1 gpc3782 (
      {stage2_24[42]},
      {stage3_24[22]}
   );
   gpc1_1 gpc3783 (
      {stage2_24[43]},
      {stage3_24[23]}
   );
   gpc1_1 gpc3784 (
      {stage2_24[44]},
      {stage3_24[24]}
   );
   gpc1_1 gpc3785 (
      {stage2_24[45]},
      {stage3_24[25]}
   );
   gpc1_1 gpc3786 (
      {stage2_25[33]},
      {stage3_25[18]}
   );
   gpc1_1 gpc3787 (
      {stage2_25[34]},
      {stage3_25[19]}
   );
   gpc1_1 gpc3788 (
      {stage2_25[35]},
      {stage3_25[20]}
   );
   gpc1_1 gpc3789 (
      {stage2_25[36]},
      {stage3_25[21]}
   );
   gpc1_1 gpc3790 (
      {stage2_27[47]},
      {stage3_27[16]}
   );
   gpc1_1 gpc3791 (
      {stage2_27[48]},
      {stage3_27[17]}
   );
   gpc1_1 gpc3792 (
      {stage2_27[49]},
      {stage3_27[18]}
   );
   gpc1_1 gpc3793 (
      {stage2_29[48]},
      {stage3_29[22]}
   );
   gpc1_1 gpc3794 (
      {stage2_29[49]},
      {stage3_29[23]}
   );
   gpc1_1 gpc3795 (
      {stage2_30[39]},
      {stage3_30[15]}
   );
   gpc1_1 gpc3796 (
      {stage2_30[40]},
      {stage3_30[16]}
   );
   gpc1_1 gpc3797 (
      {stage2_30[41]},
      {stage3_30[17]}
   );
   gpc1_1 gpc3798 (
      {stage2_30[42]},
      {stage3_30[18]}
   );
   gpc1_1 gpc3799 (
      {stage2_30[43]},
      {stage3_30[19]}
   );
   gpc1_1 gpc3800 (
      {stage2_30[44]},
      {stage3_30[20]}
   );
   gpc1_1 gpc3801 (
      {stage2_30[45]},
      {stage3_30[21]}
   );
   gpc1_1 gpc3802 (
      {stage2_30[46]},
      {stage3_30[22]}
   );
   gpc1_1 gpc3803 (
      {stage2_30[47]},
      {stage3_30[23]}
   );
   gpc1_1 gpc3804 (
      {stage2_30[48]},
      {stage3_30[24]}
   );
   gpc1_1 gpc3805 (
      {stage2_30[49]},
      {stage3_30[25]}
   );
   gpc1_1 gpc3806 (
      {stage2_31[33]},
      {stage3_31[15]}
   );
   gpc1_1 gpc3807 (
      {stage2_31[34]},
      {stage3_31[16]}
   );
   gpc1_1 gpc3808 (
      {stage2_31[35]},
      {stage3_31[17]}
   );
   gpc1_1 gpc3809 (
      {stage2_31[36]},
      {stage3_31[18]}
   );
   gpc1_1 gpc3810 (
      {stage2_31[37]},
      {stage3_31[19]}
   );
   gpc1_1 gpc3811 (
      {stage2_31[38]},
      {stage3_31[20]}
   );
   gpc1_1 gpc3812 (
      {stage2_32[36]},
      {stage3_32[15]}
   );
   gpc1_1 gpc3813 (
      {stage2_32[37]},
      {stage3_32[16]}
   );
   gpc1_1 gpc3814 (
      {stage2_32[38]},
      {stage3_32[17]}
   );
   gpc1_1 gpc3815 (
      {stage2_32[39]},
      {stage3_32[18]}
   );
   gpc1_1 gpc3816 (
      {stage2_32[40]},
      {stage3_32[19]}
   );
   gpc1_1 gpc3817 (
      {stage2_32[41]},
      {stage3_32[20]}
   );
   gpc1_1 gpc3818 (
      {stage2_32[42]},
      {stage3_32[21]}
   );
   gpc1_1 gpc3819 (
      {stage2_32[43]},
      {stage3_32[22]}
   );
   gpc1_1 gpc3820 (
      {stage2_32[44]},
      {stage3_32[23]}
   );
   gpc1_1 gpc3821 (
      {stage2_32[45]},
      {stage3_32[24]}
   );
   gpc1_1 gpc3822 (
      {stage2_32[46]},
      {stage3_32[25]}
   );
   gpc1_1 gpc3823 (
      {stage2_32[47]},
      {stage3_32[26]}
   );
   gpc1_1 gpc3824 (
      {stage2_32[48]},
      {stage3_32[27]}
   );
   gpc1_1 gpc3825 (
      {stage2_32[49]},
      {stage3_32[28]}
   );
   gpc1_1 gpc3826 (
      {stage2_32[50]},
      {stage3_32[29]}
   );
   gpc1_1 gpc3827 (
      {stage2_32[51]},
      {stage3_32[30]}
   );
   gpc1_1 gpc3828 (
      {stage2_32[52]},
      {stage3_32[31]}
   );
   gpc1_1 gpc3829 (
      {stage2_32[53]},
      {stage3_32[32]}
   );
   gpc1_1 gpc3830 (
      {stage2_32[54]},
      {stage3_32[33]}
   );
   gpc1_1 gpc3831 (
      {stage2_32[55]},
      {stage3_32[34]}
   );
   gpc1_1 gpc3832 (
      {stage2_34[23]},
      {stage3_34[11]}
   );
   gpc1_1 gpc3833 (
      {stage2_34[24]},
      {stage3_34[12]}
   );
   gpc1_1 gpc3834 (
      {stage2_34[25]},
      {stage3_34[13]}
   );
   gpc1_1 gpc3835 (
      {stage2_34[26]},
      {stage3_34[14]}
   );
   gpc1_1 gpc3836 (
      {stage2_34[27]},
      {stage3_34[15]}
   );
   gpc1_1 gpc3837 (
      {stage2_34[28]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3838 (
      {stage2_34[29]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3839 (
      {stage2_34[30]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3840 (
      {stage2_34[31]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3841 (
      {stage2_34[32]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3842 (
      {stage2_34[33]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3843 (
      {stage2_34[34]},
      {stage3_34[22]}
   );
   gpc1_1 gpc3844 (
      {stage2_35[33]},
      {stage3_35[14]}
   );
   gpc1_1 gpc3845 (
      {stage2_35[34]},
      {stage3_35[15]}
   );
   gpc1_1 gpc3846 (
      {stage2_35[35]},
      {stage3_35[16]}
   );
   gpc1_1 gpc3847 (
      {stage2_35[36]},
      {stage3_35[17]}
   );
   gpc1_1 gpc3848 (
      {stage2_35[37]},
      {stage3_35[18]}
   );
   gpc1_1 gpc3849 (
      {stage2_35[38]},
      {stage3_35[19]}
   );
   gpc1_1 gpc3850 (
      {stage2_35[39]},
      {stage3_35[20]}
   );
   gpc1_1 gpc3851 (
      {stage2_35[40]},
      {stage3_35[21]}
   );
   gpc1_1 gpc3852 (
      {stage2_35[41]},
      {stage3_35[22]}
   );
   gpc1_1 gpc3853 (
      {stage2_35[42]},
      {stage3_35[23]}
   );
   gpc1_1 gpc3854 (
      {stage2_35[43]},
      {stage3_35[24]}
   );
   gpc1_1 gpc3855 (
      {stage2_35[44]},
      {stage3_35[25]}
   );
   gpc1_1 gpc3856 (
      {stage2_36[34]},
      {stage3_36[14]}
   );
   gpc1_1 gpc3857 (
      {stage2_36[35]},
      {stage3_36[15]}
   );
   gpc1_1 gpc3858 (
      {stage2_36[36]},
      {stage3_36[16]}
   );
   gpc1_1 gpc3859 (
      {stage2_39[26]},
      {stage3_39[16]}
   );
   gpc1_1 gpc3860 (
      {stage2_39[27]},
      {stage3_39[17]}
   );
   gpc1_1 gpc3861 (
      {stage2_39[28]},
      {stage3_39[18]}
   );
   gpc1_1 gpc3862 (
      {stage2_39[29]},
      {stage3_39[19]}
   );
   gpc1_1 gpc3863 (
      {stage2_39[30]},
      {stage3_39[20]}
   );
   gpc1_1 gpc3864 (
      {stage2_39[31]},
      {stage3_39[21]}
   );
   gpc1_1 gpc3865 (
      {stage2_39[32]},
      {stage3_39[22]}
   );
   gpc1_1 gpc3866 (
      {stage2_39[33]},
      {stage3_39[23]}
   );
   gpc1_1 gpc3867 (
      {stage2_40[30]},
      {stage3_40[13]}
   );
   gpc1_1 gpc3868 (
      {stage2_40[31]},
      {stage3_40[14]}
   );
   gpc1_1 gpc3869 (
      {stage2_40[32]},
      {stage3_40[15]}
   );
   gpc1_1 gpc3870 (
      {stage2_40[33]},
      {stage3_40[16]}
   );
   gpc1_1 gpc3871 (
      {stage2_40[34]},
      {stage3_40[17]}
   );
   gpc1_1 gpc3872 (
      {stage2_40[35]},
      {stage3_40[18]}
   );
   gpc1_1 gpc3873 (
      {stage2_40[36]},
      {stage3_40[19]}
   );
   gpc1_1 gpc3874 (
      {stage2_40[37]},
      {stage3_40[20]}
   );
   gpc1_1 gpc3875 (
      {stage2_40[38]},
      {stage3_40[21]}
   );
   gpc1_1 gpc3876 (
      {stage2_40[39]},
      {stage3_40[22]}
   );
   gpc1_1 gpc3877 (
      {stage2_40[40]},
      {stage3_40[23]}
   );
   gpc1_1 gpc3878 (
      {stage2_41[45]},
      {stage3_41[14]}
   );
   gpc1_1 gpc3879 (
      {stage2_41[46]},
      {stage3_41[15]}
   );
   gpc1_1 gpc3880 (
      {stage2_41[47]},
      {stage3_41[16]}
   );
   gpc1_1 gpc3881 (
      {stage2_41[48]},
      {stage3_41[17]}
   );
   gpc1_1 gpc3882 (
      {stage2_41[49]},
      {stage3_41[18]}
   );
   gpc1_1 gpc3883 (
      {stage2_41[50]},
      {stage3_41[19]}
   );
   gpc1_1 gpc3884 (
      {stage2_41[51]},
      {stage3_41[20]}
   );
   gpc1_1 gpc3885 (
      {stage2_41[52]},
      {stage3_41[21]}
   );
   gpc1_1 gpc3886 (
      {stage2_41[53]},
      {stage3_41[22]}
   );
   gpc1_1 gpc3887 (
      {stage2_41[54]},
      {stage3_41[23]}
   );
   gpc1_1 gpc3888 (
      {stage2_41[55]},
      {stage3_41[24]}
   );
   gpc1_1 gpc3889 (
      {stage2_42[56]},
      {stage3_42[20]}
   );
   gpc1_1 gpc3890 (
      {stage2_42[57]},
      {stage3_42[21]}
   );
   gpc1_1 gpc3891 (
      {stage2_42[58]},
      {stage3_42[22]}
   );
   gpc1_1 gpc3892 (
      {stage2_42[59]},
      {stage3_42[23]}
   );
   gpc1_1 gpc3893 (
      {stage2_42[60]},
      {stage3_42[24]}
   );
   gpc1_1 gpc3894 (
      {stage2_42[61]},
      {stage3_42[25]}
   );
   gpc1_1 gpc3895 (
      {stage2_44[55]},
      {stage3_44[20]}
   );
   gpc1_1 gpc3896 (
      {stage2_44[56]},
      {stage3_44[21]}
   );
   gpc1_1 gpc3897 (
      {stage2_44[57]},
      {stage3_44[22]}
   );
   gpc1_1 gpc3898 (
      {stage2_44[58]},
      {stage3_44[23]}
   );
   gpc1_1 gpc3899 (
      {stage2_44[59]},
      {stage3_44[24]}
   );
   gpc1_1 gpc3900 (
      {stage2_44[60]},
      {stage3_44[25]}
   );
   gpc1_1 gpc3901 (
      {stage2_44[61]},
      {stage3_44[26]}
   );
   gpc1_1 gpc3902 (
      {stage2_44[62]},
      {stage3_44[27]}
   );
   gpc1_1 gpc3903 (
      {stage2_44[63]},
      {stage3_44[28]}
   );
   gpc1_1 gpc3904 (
      {stage2_44[64]},
      {stage3_44[29]}
   );
   gpc1_1 gpc3905 (
      {stage2_44[65]},
      {stage3_44[30]}
   );
   gpc1_1 gpc3906 (
      {stage2_47[37]},
      {stage3_47[15]}
   );
   gpc1_1 gpc3907 (
      {stage2_47[38]},
      {stage3_47[16]}
   );
   gpc1_1 gpc3908 (
      {stage2_47[39]},
      {stage3_47[17]}
   );
   gpc1_1 gpc3909 (
      {stage2_47[40]},
      {stage3_47[18]}
   );
   gpc1_1 gpc3910 (
      {stage2_47[41]},
      {stage3_47[19]}
   );
   gpc1_1 gpc3911 (
      {stage2_47[42]},
      {stage3_47[20]}
   );
   gpc1_1 gpc3912 (
      {stage2_47[43]},
      {stage3_47[21]}
   );
   gpc1_1 gpc3913 (
      {stage2_47[44]},
      {stage3_47[22]}
   );
   gpc1_1 gpc3914 (
      {stage2_47[45]},
      {stage3_47[23]}
   );
   gpc1_1 gpc3915 (
      {stage2_48[20]},
      {stage3_48[12]}
   );
   gpc1_1 gpc3916 (
      {stage2_48[21]},
      {stage3_48[13]}
   );
   gpc1_1 gpc3917 (
      {stage2_48[22]},
      {stage3_48[14]}
   );
   gpc1_1 gpc3918 (
      {stage2_48[23]},
      {stage3_48[15]}
   );
   gpc1_1 gpc3919 (
      {stage2_49[33]},
      {stage3_49[10]}
   );
   gpc1_1 gpc3920 (
      {stage2_49[34]},
      {stage3_49[11]}
   );
   gpc1_1 gpc3921 (
      {stage2_49[35]},
      {stage3_49[12]}
   );
   gpc1_1 gpc3922 (
      {stage2_49[36]},
      {stage3_49[13]}
   );
   gpc1_1 gpc3923 (
      {stage2_50[22]},
      {stage3_50[13]}
   );
   gpc1_1 gpc3924 (
      {stage2_50[23]},
      {stage3_50[14]}
   );
   gpc1_1 gpc3925 (
      {stage2_50[24]},
      {stage3_50[15]}
   );
   gpc1_1 gpc3926 (
      {stage2_50[25]},
      {stage3_50[16]}
   );
   gpc1_1 gpc3927 (
      {stage2_50[26]},
      {stage3_50[17]}
   );
   gpc1_1 gpc3928 (
      {stage2_50[27]},
      {stage3_50[18]}
   );
   gpc1_1 gpc3929 (
      {stage2_50[28]},
      {stage3_50[19]}
   );
   gpc1_1 gpc3930 (
      {stage2_50[29]},
      {stage3_50[20]}
   );
   gpc1_1 gpc3931 (
      {stage2_50[30]},
      {stage3_50[21]}
   );
   gpc1_1 gpc3932 (
      {stage2_50[31]},
      {stage3_50[22]}
   );
   gpc1_1 gpc3933 (
      {stage2_50[32]},
      {stage3_50[23]}
   );
   gpc1_1 gpc3934 (
      {stage2_50[33]},
      {stage3_50[24]}
   );
   gpc1_1 gpc3935 (
      {stage2_50[34]},
      {stage3_50[25]}
   );
   gpc1_1 gpc3936 (
      {stage2_50[35]},
      {stage3_50[26]}
   );
   gpc1_1 gpc3937 (
      {stage2_50[36]},
      {stage3_50[27]}
   );
   gpc1_1 gpc3938 (
      {stage2_50[37]},
      {stage3_50[28]}
   );
   gpc1_1 gpc3939 (
      {stage2_50[38]},
      {stage3_50[29]}
   );
   gpc1_1 gpc3940 (
      {stage2_50[39]},
      {stage3_50[30]}
   );
   gpc1_1 gpc3941 (
      {stage2_50[40]},
      {stage3_50[31]}
   );
   gpc1_1 gpc3942 (
      {stage2_51[24]},
      {stage3_51[13]}
   );
   gpc1_1 gpc3943 (
      {stage2_52[18]},
      {stage3_52[8]}
   );
   gpc1_1 gpc3944 (
      {stage2_52[19]},
      {stage3_52[9]}
   );
   gpc1_1 gpc3945 (
      {stage2_52[20]},
      {stage3_52[10]}
   );
   gpc1_1 gpc3946 (
      {stage2_52[21]},
      {stage3_52[11]}
   );
   gpc1_1 gpc3947 (
      {stage2_52[22]},
      {stage3_52[12]}
   );
   gpc1_1 gpc3948 (
      {stage2_52[23]},
      {stage3_52[13]}
   );
   gpc1_1 gpc3949 (
      {stage2_52[24]},
      {stage3_52[14]}
   );
   gpc1_1 gpc3950 (
      {stage2_52[25]},
      {stage3_52[15]}
   );
   gpc1_1 gpc3951 (
      {stage2_52[26]},
      {stage3_52[16]}
   );
   gpc1_1 gpc3952 (
      {stage2_52[27]},
      {stage3_52[17]}
   );
   gpc1_1 gpc3953 (
      {stage2_52[28]},
      {stage3_52[18]}
   );
   gpc1_1 gpc3954 (
      {stage2_52[29]},
      {stage3_52[19]}
   );
   gpc1_1 gpc3955 (
      {stage2_52[30]},
      {stage3_52[20]}
   );
   gpc1_1 gpc3956 (
      {stage2_52[31]},
      {stage3_52[21]}
   );
   gpc1_1 gpc3957 (
      {stage2_52[32]},
      {stage3_52[22]}
   );
   gpc1_1 gpc3958 (
      {stage2_52[33]},
      {stage3_52[23]}
   );
   gpc1_1 gpc3959 (
      {stage2_53[46]},
      {stage3_53[11]}
   );
   gpc1_1 gpc3960 (
      {stage2_53[47]},
      {stage3_53[12]}
   );
   gpc1_1 gpc3961 (
      {stage2_53[48]},
      {stage3_53[13]}
   );
   gpc1_1 gpc3962 (
      {stage2_53[49]},
      {stage3_53[14]}
   );
   gpc1_1 gpc3963 (
      {stage2_53[50]},
      {stage3_53[15]}
   );
   gpc1_1 gpc3964 (
      {stage2_55[35]},
      {stage3_55[15]}
   );
   gpc1_1 gpc3965 (
      {stage2_55[36]},
      {stage3_55[16]}
   );
   gpc1_1 gpc3966 (
      {stage2_55[37]},
      {stage3_55[17]}
   );
   gpc1_1 gpc3967 (
      {stage2_56[33]},
      {stage3_56[11]}
   );
   gpc1_1 gpc3968 (
      {stage2_56[34]},
      {stage3_56[12]}
   );
   gpc1_1 gpc3969 (
      {stage2_56[35]},
      {stage3_56[13]}
   );
   gpc1_1 gpc3970 (
      {stage2_56[36]},
      {stage3_56[14]}
   );
   gpc1_1 gpc3971 (
      {stage2_56[37]},
      {stage3_56[15]}
   );
   gpc1_1 gpc3972 (
      {stage2_56[38]},
      {stage3_56[16]}
   );
   gpc1_1 gpc3973 (
      {stage2_56[39]},
      {stage3_56[17]}
   );
   gpc1_1 gpc3974 (
      {stage2_56[40]},
      {stage3_56[18]}
   );
   gpc1_1 gpc3975 (
      {stage2_56[41]},
      {stage3_56[19]}
   );
   gpc1_1 gpc3976 (
      {stage2_56[42]},
      {stage3_56[20]}
   );
   gpc1_1 gpc3977 (
      {stage2_56[43]},
      {stage3_56[21]}
   );
   gpc1_1 gpc3978 (
      {stage2_56[44]},
      {stage3_56[22]}
   );
   gpc1_1 gpc3979 (
      {stage2_56[45]},
      {stage3_56[23]}
   );
   gpc1_1 gpc3980 (
      {stage2_56[46]},
      {stage3_56[24]}
   );
   gpc1_1 gpc3981 (
      {stage2_56[47]},
      {stage3_56[25]}
   );
   gpc1_1 gpc3982 (
      {stage2_56[48]},
      {stage3_56[26]}
   );
   gpc1_1 gpc3983 (
      {stage2_56[49]},
      {stage3_56[27]}
   );
   gpc1_1 gpc3984 (
      {stage2_56[50]},
      {stage3_56[28]}
   );
   gpc1_1 gpc3985 (
      {stage2_56[51]},
      {stage3_56[29]}
   );
   gpc1_1 gpc3986 (
      {stage2_56[52]},
      {stage3_56[30]}
   );
   gpc1_1 gpc3987 (
      {stage2_58[13]},
      {stage3_58[13]}
   );
   gpc1_1 gpc3988 (
      {stage2_58[14]},
      {stage3_58[14]}
   );
   gpc1_1 gpc3989 (
      {stage2_58[15]},
      {stage3_58[15]}
   );
   gpc1_1 gpc3990 (
      {stage2_58[16]},
      {stage3_58[16]}
   );
   gpc1_1 gpc3991 (
      {stage2_58[17]},
      {stage3_58[17]}
   );
   gpc1_1 gpc3992 (
      {stage2_58[18]},
      {stage3_58[18]}
   );
   gpc1_1 gpc3993 (
      {stage2_58[19]},
      {stage3_58[19]}
   );
   gpc1_1 gpc3994 (
      {stage2_58[20]},
      {stage3_58[20]}
   );
   gpc1_1 gpc3995 (
      {stage2_58[21]},
      {stage3_58[21]}
   );
   gpc1_1 gpc3996 (
      {stage2_58[22]},
      {stage3_58[22]}
   );
   gpc1_1 gpc3997 (
      {stage2_58[23]},
      {stage3_58[23]}
   );
   gpc1_1 gpc3998 (
      {stage2_58[24]},
      {stage3_58[24]}
   );
   gpc1_1 gpc3999 (
      {stage2_58[25]},
      {stage3_58[25]}
   );
   gpc1_1 gpc4000 (
      {stage2_58[26]},
      {stage3_58[26]}
   );
   gpc1_1 gpc4001 (
      {stage2_58[27]},
      {stage3_58[27]}
   );
   gpc1_1 gpc4002 (
      {stage2_58[28]},
      {stage3_58[28]}
   );
   gpc1_1 gpc4003 (
      {stage2_58[29]},
      {stage3_58[29]}
   );
   gpc1_1 gpc4004 (
      {stage2_58[30]},
      {stage3_58[30]}
   );
   gpc1_1 gpc4005 (
      {stage2_58[31]},
      {stage3_58[31]}
   );
   gpc1_1 gpc4006 (
      {stage2_58[32]},
      {stage3_58[32]}
   );
   gpc1_1 gpc4007 (
      {stage2_59[70]},
      {stage3_59[17]}
   );
   gpc1_1 gpc4008 (
      {stage2_59[71]},
      {stage3_59[18]}
   );
   gpc1_1 gpc4009 (
      {stage2_59[72]},
      {stage3_59[19]}
   );
   gpc1_1 gpc4010 (
      {stage2_59[73]},
      {stage3_59[20]}
   );
   gpc1_1 gpc4011 (
      {stage2_59[74]},
      {stage3_59[21]}
   );
   gpc1_1 gpc4012 (
      {stage2_59[75]},
      {stage3_59[22]}
   );
   gpc1_1 gpc4013 (
      {stage2_59[76]},
      {stage3_59[23]}
   );
   gpc1_1 gpc4014 (
      {stage2_59[77]},
      {stage3_59[24]}
   );
   gpc1_1 gpc4015 (
      {stage2_59[78]},
      {stage3_59[25]}
   );
   gpc1_1 gpc4016 (
      {stage2_59[79]},
      {stage3_59[26]}
   );
   gpc1_1 gpc4017 (
      {stage2_59[80]},
      {stage3_59[27]}
   );
   gpc1_1 gpc4018 (
      {stage2_61[59]},
      {stage3_61[17]}
   );
   gpc1_1 gpc4019 (
      {stage2_61[60]},
      {stage3_61[18]}
   );
   gpc1_1 gpc4020 (
      {stage2_61[61]},
      {stage3_61[19]}
   );
   gpc1_1 gpc4021 (
      {stage2_61[62]},
      {stage3_61[20]}
   );
   gpc1_1 gpc4022 (
      {stage2_61[63]},
      {stage3_61[21]}
   );
   gpc1_1 gpc4023 (
      {stage2_61[64]},
      {stage3_61[22]}
   );
   gpc1_1 gpc4024 (
      {stage2_61[65]},
      {stage3_61[23]}
   );
   gpc1_1 gpc4025 (
      {stage2_61[66]},
      {stage3_61[24]}
   );
   gpc1_1 gpc4026 (
      {stage2_64[29]},
      {stage3_64[12]}
   );
   gpc1_1 gpc4027 (
      {stage2_64[30]},
      {stage3_64[13]}
   );
   gpc1_1 gpc4028 (
      {stage2_64[31]},
      {stage3_64[14]}
   );
   gpc1_1 gpc4029 (
      {stage2_64[32]},
      {stage3_64[15]}
   );
   gpc1_1 gpc4030 (
      {stage2_64[33]},
      {stage3_64[16]}
   );
   gpc1_1 gpc4031 (
      {stage2_64[34]},
      {stage3_64[17]}
   );
   gpc1_1 gpc4032 (
      {stage2_64[35]},
      {stage3_64[18]}
   );
   gpc1_1 gpc4033 (
      {stage2_64[36]},
      {stage3_64[19]}
   );
   gpc1_1 gpc4034 (
      {stage2_64[37]},
      {stage3_64[20]}
   );
   gpc1_1 gpc4035 (
      {stage2_64[38]},
      {stage3_64[21]}
   );
   gpc1_1 gpc4036 (
      {stage2_64[39]},
      {stage3_64[22]}
   );
   gpc1_1 gpc4037 (
      {stage2_64[40]},
      {stage3_64[23]}
   );
   gpc1_1 gpc4038 (
      {stage2_64[41]},
      {stage3_64[24]}
   );
   gpc1_1 gpc4039 (
      {stage2_64[42]},
      {stage3_64[25]}
   );
   gpc1_1 gpc4040 (
      {stage2_64[43]},
      {stage3_64[26]}
   );
   gpc1_1 gpc4041 (
      {stage2_64[44]},
      {stage3_64[27]}
   );
   gpc1_1 gpc4042 (
      {stage2_64[45]},
      {stage3_64[28]}
   );
   gpc1_1 gpc4043 (
      {stage2_65[10]},
      {stage3_65[11]}
   );
   gpc1_1 gpc4044 (
      {stage2_65[11]},
      {stage3_65[12]}
   );
   gpc1_1 gpc4045 (
      {stage2_65[12]},
      {stage3_65[13]}
   );
   gpc1_1 gpc4046 (
      {stage2_67[0]},
      {stage3_67[3]}
   );
   gpc1_1 gpc4047 (
      {stage2_67[1]},
      {stage3_67[4]}
   );
   gpc1163_5 gpc4048 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1163_5 gpc4049 (
      {stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_2[1]},
      {stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc4050 (
      {stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6]},
      {stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4051 (
      {stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc4052 (
      {stage3_3[9], stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], 1'b0},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc4053 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[12]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[5]}
   );
   gpc615_5 gpc4054 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4]}
   );
   gpc207_4 gpc4055 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4]}
   );
   gpc207_4 gpc4056 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_9[2], stage3_9[3]},
      {stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc4057 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[3],stage4_8[4]}
   );
   gpc2135_5 gpc4058 (
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[6], stage3_10[7], stage3_10[8]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc4059 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6]},
      {stage4_13[1],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[5]}
   );
   gpc606_5 gpc4060 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12]},
      {stage4_13[2],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[6]}
   );
   gpc2135_5 gpc4061 (
      {stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage3_11[13], stage3_11[14], stage3_11[15]},
      {stage3_12[2]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[3],stage4_12[4],stage4_11[4],stage4_10[7]}
   );
   gpc207_4 gpc4062 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[5]}
   );
   gpc207_4 gpc4063 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16]},
      {stage3_14[2], stage3_14[3]},
      {stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[6]}
   );
   gpc606_5 gpc4064 (
      {stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22]},
      {stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage4_16[0],stage4_15[2],stage4_14[3],stage4_13[6],stage4_12[7]}
   );
   gpc606_5 gpc4065 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc606_5 gpc4066 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[4],stage4_14[5],stage4_13[8]}
   );
   gpc606_5 gpc4067 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[3],stage4_15[5],stage4_14[6],stage4_13[9]}
   );
   gpc117_4 gpc4068 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[18]},
      {stage3_16[0]},
      {stage4_17[3],stage4_16[4],stage4_15[6],stage4_14[7]}
   );
   gpc117_4 gpc4069 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_15[19]},
      {stage3_16[1]},
      {stage4_17[4],stage4_16[5],stage4_15[7],stage4_14[8]}
   );
   gpc117_4 gpc4070 (
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[20]},
      {stage3_16[2]},
      {stage4_17[5],stage4_16[6],stage4_15[8],stage4_14[9]}
   );
   gpc117_4 gpc4071 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], 1'b0, 1'b0},
      {stage3_15[21]},
      {stage3_16[3]},
      {stage4_17[6],stage4_16[7],stage4_15[9],stage4_14[10]}
   );
   gpc615_5 gpc4072 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[4]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[0],stage4_17[7],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc4073 (
      {stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31]},
      {stage3_16[5]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[1],stage4_17[8],stage4_16[9],stage4_15[11]}
   );
   gpc606_5 gpc4074 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[2],stage4_18[2],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc4075 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[3],stage4_18[3],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc4076 (
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], 1'b0, 1'b0},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[4],stage4_18[4],stage4_17[11],stage4_16[12]}
   );
   gpc615_5 gpc4077 (
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[3],stage4_19[5],stage4_18[5]}
   );
   gpc615_5 gpc4078 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[1],stage4_21[1],stage4_20[4],stage4_19[6]}
   );
   gpc615_5 gpc4079 (
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10]},
      {stage3_20[7]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[2],stage4_21[2],stage4_20[5],stage4_19[7]}
   );
   gpc615_5 gpc4080 (
      {stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15]},
      {stage3_20[8]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[3],stage4_21[3],stage4_20[6],stage4_19[8]}
   );
   gpc615_5 gpc4081 (
      {stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20]},
      {stage3_20[9]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[4],stage4_21[4],stage4_20[7],stage4_19[9]}
   );
   gpc606_5 gpc4082 (
      {stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[4],stage4_22[5],stage4_21[5],stage4_20[8]}
   );
   gpc606_5 gpc4083 (
      {stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[5],stage4_22[6],stage4_21[6],stage4_20[9]}
   );
   gpc615_5 gpc4084 (
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage3_23[0]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[6],stage4_22[7]}
   );
   gpc615_5 gpc4085 (
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21]},
      {stage3_23[1]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[1],stage4_24[3],stage4_23[7],stage4_22[8]}
   );
   gpc615_5 gpc4086 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[2],stage4_24[4],stage4_23[8]}
   );
   gpc615_5 gpc4087 (
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[3],stage4_24[5],stage4_23[9]}
   );
   gpc615_5 gpc4088 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[2],stage4_26[4],stage4_25[4]}
   );
   gpc615_5 gpc4089 (
      {stage3_25[17], stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21]},
      {stage3_26[1]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[3],stage4_26[5],stage4_25[5]}
   );
   gpc117_4 gpc4090 (
      {stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[12]},
      {stage3_28[0]},
      {stage4_29[2],stage4_28[2],stage4_27[4],stage4_26[6]}
   );
   gpc207_4 gpc4091 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15]},
      {stage3_28[1], stage3_28[2]},
      {stage4_29[3],stage4_28[3],stage4_27[5],stage4_26[7]}
   );
   gpc606_5 gpc4092 (
      {stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17], stage3_27[18]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[4],stage4_28[4],stage4_27[6]}
   );
   gpc606_5 gpc4093 (
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[5],stage4_28[5]}
   );
   gpc606_5 gpc4094 (
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[6],stage4_28[6]}
   );
   gpc606_5 gpc4095 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[3],stage4_30[3],stage4_29[7]}
   );
   gpc606_5 gpc4096 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[4],stage4_30[4],stage4_29[8]}
   );
   gpc606_5 gpc4097 (
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[5],stage4_30[5],stage4_29[9]}
   );
   gpc615_5 gpc4098 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16]},
      {stage3_31[18]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[6],stage4_30[6]}
   );
   gpc606_5 gpc4099 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6]}
   );
   gpc606_5 gpc4100 (
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7]}
   );
   gpc606_5 gpc4101 (
      {stage3_32[18], stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc4102 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[3],stage4_35[3],stage4_34[4],stage4_33[7]}
   );
   gpc606_5 gpc4103 (
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[1],stage4_36[4],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1343_5 gpc4104 (
      {stage3_35[12], stage3_35[13], stage3_35[14]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3]},
      {stage3_37[0], stage3_37[1], stage3_37[2]},
      {stage3_38[0]},
      {stage4_39[0],stage4_38[0],stage4_37[2],stage4_36[5],stage4_35[5]}
   );
   gpc1343_5 gpc4105 (
      {stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7]},
      {stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_38[1]},
      {stage4_39[1],stage4_38[1],stage4_37[3],stage4_36[6],stage4_35[6]}
   );
   gpc1343_5 gpc4106 (
      {stage3_35[18], stage3_35[19], stage3_35[20]},
      {stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11]},
      {stage3_37[6], stage3_37[7], stage3_37[8]},
      {stage3_38[2]},
      {stage4_39[2],stage4_38[2],stage4_37[4],stage4_36[7],stage4_35[7]}
   );
   gpc1343_5 gpc4107 (
      {stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15]},
      {stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage3_38[3]},
      {stage4_39[3],stage4_38[3],stage4_37[5],stage4_36[8],stage4_35[8]}
   );
   gpc615_5 gpc4108 (
      {stage3_38[4], stage3_38[5], stage3_38[6], stage3_38[7], stage3_38[8]},
      {stage3_39[0]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[0],stage4_40[0],stage4_39[4],stage4_38[4]}
   );
   gpc615_5 gpc4109 (
      {stage3_38[9], stage3_38[10], stage3_38[11], stage3_38[12], stage3_38[13]},
      {stage3_39[1]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[1],stage4_40[1],stage4_39[5],stage4_38[5]}
   );
   gpc117_4 gpc4110 (
      {stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5], stage3_39[6], stage3_39[7], stage3_39[8]},
      {stage3_40[12]},
      {stage3_41[0]},
      {stage4_42[2],stage4_41[2],stage4_40[2],stage4_39[6]}
   );
   gpc117_4 gpc4111 (
      {stage3_39[9], stage3_39[10], stage3_39[11], stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15]},
      {stage3_40[13]},
      {stage3_41[1]},
      {stage4_42[3],stage4_41[3],stage4_40[3],stage4_39[7]}
   );
   gpc117_4 gpc4112 (
      {stage3_39[16], stage3_39[17], stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22]},
      {stage3_40[14]},
      {stage3_41[2]},
      {stage4_42[4],stage4_41[4],stage4_40[4],stage4_39[8]}
   );
   gpc606_5 gpc4113 (
      {stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], stage3_41[7], stage3_41[8]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[5],stage4_41[5]}
   );
   gpc606_5 gpc4114 (
      {stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13], stage3_41[14]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[6],stage4_41[6]}
   );
   gpc615_5 gpc4115 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4]},
      {stage3_43[12]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[7]}
   );
   gpc615_5 gpc4116 (
      {stage3_42[5], stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9]},
      {stage3_43[13]},
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11]},
      {stage4_46[1],stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[8]}
   );
   gpc615_5 gpc4117 (
      {stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13], stage3_42[14]},
      {stage3_43[14]},
      {stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15], stage3_44[16], stage3_44[17]},
      {stage4_46[2],stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[9]}
   );
   gpc615_5 gpc4118 (
      {stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19]},
      {stage3_43[15]},
      {stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21], stage3_44[22], stage3_44[23]},
      {stage4_46[3],stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[10]}
   );
   gpc615_5 gpc4119 (
      {stage3_43[16], stage3_43[17], stage3_43[18], stage3_43[19], stage3_43[20]},
      {stage3_44[24]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[4],stage4_45[6],stage4_44[6],stage4_43[6]}
   );
   gpc606_5 gpc4120 (
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage3_47[0], stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5]},
      {stage4_49[0],stage4_48[0],stage4_47[1],stage4_46[5],stage4_45[7]}
   );
   gpc606_5 gpc4121 (
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_47[6], stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], stage3_47[11]},
      {stage4_49[1],stage4_48[1],stage4_47[2],stage4_46[6],stage4_45[8]}
   );
   gpc207_4 gpc4122 (
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_48[0], stage3_48[1]},
      {stage4_49[2],stage4_48[2],stage4_47[3],stage4_46[7]}
   );
   gpc606_5 gpc4123 (
      {stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5], stage3_48[6], stage3_48[7]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[0],stage4_50[0],stage4_49[3],stage4_48[3]}
   );
   gpc606_5 gpc4124 (
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[1],stage4_51[1],stage4_50[1],stage4_49[4]}
   );
   gpc7_3 gpc4125 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12]},
      {stage4_52[2],stage4_51[2],stage4_50[2]}
   );
   gpc606_5 gpc4126 (
      {stage3_50[13], stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[1],stage4_52[3],stage4_51[3],stage4_50[3]}
   );
   gpc606_5 gpc4127 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24]},
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage4_54[1],stage4_53[2],stage4_52[4],stage4_51[4],stage4_50[4]}
   );
   gpc606_5 gpc4128 (
      {stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28], stage3_50[29], stage3_50[30]},
      {stage3_52[12], stage3_52[13], stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage4_54[2],stage4_53[3],stage4_52[5],stage4_51[5],stage4_50[5]}
   );
   gpc606_5 gpc4129 (
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[3],stage4_53[4],stage4_52[6],stage4_51[6]}
   );
   gpc615_5 gpc4130 (
      {stage3_52[18], stage3_52[19], stage3_52[20], stage3_52[21], stage3_52[22]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[4],stage4_53[5],stage4_52[7]}
   );
   gpc606_5 gpc4131 (
      {stage3_54[6], stage3_54[7], stage3_54[8], stage3_54[9], stage3_54[10], stage3_54[11]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2],stage4_54[5]}
   );
   gpc615_5 gpc4132 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4]},
      {stage3_56[6]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc606_5 gpc4133 (
      {stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[1],stage4_58[2],stage4_57[2],stage4_56[3]}
   );
   gpc606_5 gpc4134 (
      {stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[2],stage4_58[3],stage4_57[3],stage4_56[4]}
   );
   gpc615_5 gpc4135 (
      {stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage3_57[6]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[3],stage4_58[4],stage4_57[4],stage4_56[5]}
   );
   gpc606_5 gpc4136 (
      {stage3_57[7], stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[3],stage4_59[4],stage4_58[5],stage4_57[5]}
   );
   gpc606_5 gpc4137 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[4],stage4_59[5]}
   );
   gpc606_5 gpc4138 (
      {stage3_59[12], stage3_59[13], stage3_59[14], stage3_59[15], stage3_59[16], stage3_59[17]},
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[5],stage4_59[6]}
   );
   gpc606_5 gpc4139 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[2],stage4_62[2],stage4_61[3],stage4_60[6]}
   );
   gpc606_5 gpc4140 (
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[0],stage4_64[1],stage4_63[3],stage4_62[3]}
   );
   gpc606_5 gpc4141 (
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage4_66[1],stage4_65[1],stage4_64[2],stage4_63[4],stage4_62[4]}
   );
   gpc606_5 gpc4142 (
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[2],stage4_65[2],stage4_64[3],stage4_63[5]}
   );
   gpc606_5 gpc4143 (
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[3],stage4_65[3],stage4_64[4],stage4_63[6]}
   );
   gpc1_1 gpc4144 (
      {stage3_0[6]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4145 (
      {stage3_0[7]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4146 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4147 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4148 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc4149 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc4150 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc4151 (
      {stage3_2[10]},
      {stage4_2[6]}
   );
   gpc1_1 gpc4152 (
      {stage3_4[11]},
      {stage4_4[6]}
   );
   gpc1_1 gpc4153 (
      {stage3_4[12]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4154 (
      {stage3_4[13]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4155 (
      {stage3_5[13]},
      {stage4_5[4]}
   );
   gpc1_1 gpc4156 (
      {stage3_5[14]},
      {stage4_5[5]}
   );
   gpc1_1 gpc4157 (
      {stage3_5[15]},
      {stage4_5[6]}
   );
   gpc1_1 gpc4158 (
      {stage3_5[16]},
      {stage4_5[7]}
   );
   gpc1_1 gpc4159 (
      {stage3_5[17]},
      {stage4_5[8]}
   );
   gpc1_1 gpc4160 (
      {stage3_6[11]},
      {stage4_6[5]}
   );
   gpc1_1 gpc4161 (
      {stage3_6[12]},
      {stage4_6[6]}
   );
   gpc1_1 gpc4162 (
      {stage3_6[13]},
      {stage4_6[7]}
   );
   gpc1_1 gpc4163 (
      {stage3_6[14]},
      {stage4_6[8]}
   );
   gpc1_1 gpc4164 (
      {stage3_6[15]},
      {stage4_6[9]}
   );
   gpc1_1 gpc4165 (
      {stage3_6[16]},
      {stage4_6[10]}
   );
   gpc1_1 gpc4166 (
      {stage3_6[17]},
      {stage4_6[11]}
   );
   gpc1_1 gpc4167 (
      {stage3_6[18]},
      {stage4_6[12]}
   );
   gpc1_1 gpc4168 (
      {stage3_6[19]},
      {stage4_6[13]}
   );
   gpc1_1 gpc4169 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc4170 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc4171 (
      {stage3_8[12]},
      {stage4_8[5]}
   );
   gpc1_1 gpc4172 (
      {stage3_8[13]},
      {stage4_8[6]}
   );
   gpc1_1 gpc4173 (
      {stage3_8[14]},
      {stage4_8[7]}
   );
   gpc1_1 gpc4174 (
      {stage3_8[15]},
      {stage4_8[8]}
   );
   gpc1_1 gpc4175 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc4176 (
      {stage3_10[14]},
      {stage4_10[8]}
   );
   gpc1_1 gpc4177 (
      {stage3_11[16]},
      {stage4_11[5]}
   );
   gpc1_1 gpc4178 (
      {stage3_11[17]},
      {stage4_11[6]}
   );
   gpc1_1 gpc4179 (
      {stage3_12[23]},
      {stage4_12[8]}
   );
   gpc1_1 gpc4180 (
      {stage3_15[32]},
      {stage4_15[12]}
   );
   gpc1_1 gpc4181 (
      {stage3_15[33]},
      {stage4_15[13]}
   );
   gpc1_1 gpc4182 (
      {stage3_15[34]},
      {stage4_15[14]}
   );
   gpc1_1 gpc4183 (
      {stage3_15[35]},
      {stage4_15[15]}
   );
   gpc1_1 gpc4184 (
      {stage3_15[36]},
      {stage4_15[16]}
   );
   gpc1_1 gpc4185 (
      {stage3_17[12]},
      {stage4_17[12]}
   );
   gpc1_1 gpc4186 (
      {stage3_17[13]},
      {stage4_17[13]}
   );
   gpc1_1 gpc4187 (
      {stage3_17[14]},
      {stage4_17[14]}
   );
   gpc1_1 gpc4188 (
      {stage3_17[15]},
      {stage4_17[15]}
   );
   gpc1_1 gpc4189 (
      {stage3_17[16]},
      {stage4_17[16]}
   );
   gpc1_1 gpc4190 (
      {stage3_19[21]},
      {stage4_19[10]}
   );
   gpc1_1 gpc4191 (
      {stage3_19[22]},
      {stage4_19[11]}
   );
   gpc1_1 gpc4192 (
      {stage3_19[23]},
      {stage4_19[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_19[24]},
      {stage4_19[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_19[25]},
      {stage4_19[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_19[26]},
      {stage4_19[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_20[22]},
      {stage4_20[10]}
   );
   gpc1_1 gpc4197 (
      {stage3_21[24]},
      {stage4_21[7]}
   );
   gpc1_1 gpc4198 (
      {stage3_22[22]},
      {stage4_22[9]}
   );
   gpc1_1 gpc4199 (
      {stage3_22[23]},
      {stage4_22[10]}
   );
   gpc1_1 gpc4200 (
      {stage3_22[24]},
      {stage4_22[11]}
   );
   gpc1_1 gpc4201 (
      {stage3_22[25]},
      {stage4_22[12]}
   );
   gpc1_1 gpc4202 (
      {stage3_22[26]},
      {stage4_22[13]}
   );
   gpc1_1 gpc4203 (
      {stage3_24[14]},
      {stage4_24[6]}
   );
   gpc1_1 gpc4204 (
      {stage3_24[15]},
      {stage4_24[7]}
   );
   gpc1_1 gpc4205 (
      {stage3_24[16]},
      {stage4_24[8]}
   );
   gpc1_1 gpc4206 (
      {stage3_24[17]},
      {stage4_24[9]}
   );
   gpc1_1 gpc4207 (
      {stage3_24[18]},
      {stage4_24[10]}
   );
   gpc1_1 gpc4208 (
      {stage3_24[19]},
      {stage4_24[11]}
   );
   gpc1_1 gpc4209 (
      {stage3_24[20]},
      {stage4_24[12]}
   );
   gpc1_1 gpc4210 (
      {stage3_24[21]},
      {stage4_24[13]}
   );
   gpc1_1 gpc4211 (
      {stage3_24[22]},
      {stage4_24[14]}
   );
   gpc1_1 gpc4212 (
      {stage3_24[23]},
      {stage4_24[15]}
   );
   gpc1_1 gpc4213 (
      {stage3_24[24]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4214 (
      {stage3_24[25]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4215 (
      {stage3_28[15]},
      {stage4_28[7]}
   );
   gpc1_1 gpc4216 (
      {stage3_28[16]},
      {stage4_28[8]}
   );
   gpc1_1 gpc4217 (
      {stage3_28[17]},
      {stage4_28[9]}
   );
   gpc1_1 gpc4218 (
      {stage3_28[18]},
      {stage4_28[10]}
   );
   gpc1_1 gpc4219 (
      {stage3_28[19]},
      {stage4_28[11]}
   );
   gpc1_1 gpc4220 (
      {stage3_30[17]},
      {stage4_30[7]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[18]},
      {stage4_30[8]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[19]},
      {stage4_30[9]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[20]},
      {stage4_30[10]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[21]},
      {stage4_30[11]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[22]},
      {stage4_30[12]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[23]},
      {stage4_30[13]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[24]},
      {stage4_30[14]}
   );
   gpc1_1 gpc4228 (
      {stage3_30[25]},
      {stage4_30[15]}
   );
   gpc1_1 gpc4229 (
      {stage3_31[19]},
      {stage4_31[7]}
   );
   gpc1_1 gpc4230 (
      {stage3_31[20]},
      {stage4_31[8]}
   );
   gpc1_1 gpc4231 (
      {stage3_32[24]},
      {stage4_32[9]}
   );
   gpc1_1 gpc4232 (
      {stage3_32[25]},
      {stage4_32[10]}
   );
   gpc1_1 gpc4233 (
      {stage3_32[26]},
      {stage4_32[11]}
   );
   gpc1_1 gpc4234 (
      {stage3_32[27]},
      {stage4_32[12]}
   );
   gpc1_1 gpc4235 (
      {stage3_32[28]},
      {stage4_32[13]}
   );
   gpc1_1 gpc4236 (
      {stage3_32[29]},
      {stage4_32[14]}
   );
   gpc1_1 gpc4237 (
      {stage3_32[30]},
      {stage4_32[15]}
   );
   gpc1_1 gpc4238 (
      {stage3_32[31]},
      {stage4_32[16]}
   );
   gpc1_1 gpc4239 (
      {stage3_32[32]},
      {stage4_32[17]}
   );
   gpc1_1 gpc4240 (
      {stage3_32[33]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4241 (
      {stage3_32[34]},
      {stage4_32[19]}
   );
   gpc1_1 gpc4242 (
      {stage3_33[12]},
      {stage4_33[9]}
   );
   gpc1_1 gpc4243 (
      {stage3_33[13]},
      {stage4_33[10]}
   );
   gpc1_1 gpc4244 (
      {stage3_33[14]},
      {stage4_33[11]}
   );
   gpc1_1 gpc4245 (
      {stage3_34[18]},
      {stage4_34[6]}
   );
   gpc1_1 gpc4246 (
      {stage3_34[19]},
      {stage4_34[7]}
   );
   gpc1_1 gpc4247 (
      {stage3_34[20]},
      {stage4_34[8]}
   );
   gpc1_1 gpc4248 (
      {stage3_34[21]},
      {stage4_34[9]}
   );
   gpc1_1 gpc4249 (
      {stage3_34[22]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4250 (
      {stage3_35[24]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4251 (
      {stage3_35[25]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4252 (
      {stage3_36[16]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4253 (
      {stage3_39[23]},
      {stage4_39[9]}
   );
   gpc1_1 gpc4254 (
      {stage3_40[15]},
      {stage4_40[5]}
   );
   gpc1_1 gpc4255 (
      {stage3_40[16]},
      {stage4_40[6]}
   );
   gpc1_1 gpc4256 (
      {stage3_40[17]},
      {stage4_40[7]}
   );
   gpc1_1 gpc4257 (
      {stage3_40[18]},
      {stage4_40[8]}
   );
   gpc1_1 gpc4258 (
      {stage3_40[19]},
      {stage4_40[9]}
   );
   gpc1_1 gpc4259 (
      {stage3_40[20]},
      {stage4_40[10]}
   );
   gpc1_1 gpc4260 (
      {stage3_40[21]},
      {stage4_40[11]}
   );
   gpc1_1 gpc4261 (
      {stage3_40[22]},
      {stage4_40[12]}
   );
   gpc1_1 gpc4262 (
      {stage3_40[23]},
      {stage4_40[13]}
   );
   gpc1_1 gpc4263 (
      {stage3_41[15]},
      {stage4_41[7]}
   );
   gpc1_1 gpc4264 (
      {stage3_41[16]},
      {stage4_41[8]}
   );
   gpc1_1 gpc4265 (
      {stage3_41[17]},
      {stage4_41[9]}
   );
   gpc1_1 gpc4266 (
      {stage3_41[18]},
      {stage4_41[10]}
   );
   gpc1_1 gpc4267 (
      {stage3_41[19]},
      {stage4_41[11]}
   );
   gpc1_1 gpc4268 (
      {stage3_41[20]},
      {stage4_41[12]}
   );
   gpc1_1 gpc4269 (
      {stage3_41[21]},
      {stage4_41[13]}
   );
   gpc1_1 gpc4270 (
      {stage3_41[22]},
      {stage4_41[14]}
   );
   gpc1_1 gpc4271 (
      {stage3_41[23]},
      {stage4_41[15]}
   );
   gpc1_1 gpc4272 (
      {stage3_41[24]},
      {stage4_41[16]}
   );
   gpc1_1 gpc4273 (
      {stage3_42[20]},
      {stage4_42[11]}
   );
   gpc1_1 gpc4274 (
      {stage3_42[21]},
      {stage4_42[12]}
   );
   gpc1_1 gpc4275 (
      {stage3_42[22]},
      {stage4_42[13]}
   );
   gpc1_1 gpc4276 (
      {stage3_42[23]},
      {stage4_42[14]}
   );
   gpc1_1 gpc4277 (
      {stage3_42[24]},
      {stage4_42[15]}
   );
   gpc1_1 gpc4278 (
      {stage3_42[25]},
      {stage4_42[16]}
   );
   gpc1_1 gpc4279 (
      {stage3_44[25]},
      {stage4_44[7]}
   );
   gpc1_1 gpc4280 (
      {stage3_44[26]},
      {stage4_44[8]}
   );
   gpc1_1 gpc4281 (
      {stage3_44[27]},
      {stage4_44[9]}
   );
   gpc1_1 gpc4282 (
      {stage3_44[28]},
      {stage4_44[10]}
   );
   gpc1_1 gpc4283 (
      {stage3_44[29]},
      {stage4_44[11]}
   );
   gpc1_1 gpc4284 (
      {stage3_44[30]},
      {stage4_44[12]}
   );
   gpc1_1 gpc4285 (
      {stage3_46[7]},
      {stage4_46[8]}
   );
   gpc1_1 gpc4286 (
      {stage3_46[8]},
      {stage4_46[9]}
   );
   gpc1_1 gpc4287 (
      {stage3_46[9]},
      {stage4_46[10]}
   );
   gpc1_1 gpc4288 (
      {stage3_46[10]},
      {stage4_46[11]}
   );
   gpc1_1 gpc4289 (
      {stage3_46[11]},
      {stage4_46[12]}
   );
   gpc1_1 gpc4290 (
      {stage3_46[12]},
      {stage4_46[13]}
   );
   gpc1_1 gpc4291 (
      {stage3_46[13]},
      {stage4_46[14]}
   );
   gpc1_1 gpc4292 (
      {stage3_46[14]},
      {stage4_46[15]}
   );
   gpc1_1 gpc4293 (
      {stage3_46[15]},
      {stage4_46[16]}
   );
   gpc1_1 gpc4294 (
      {stage3_46[16]},
      {stage4_46[17]}
   );
   gpc1_1 gpc4295 (
      {stage3_47[12]},
      {stage4_47[4]}
   );
   gpc1_1 gpc4296 (
      {stage3_47[13]},
      {stage4_47[5]}
   );
   gpc1_1 gpc4297 (
      {stage3_47[14]},
      {stage4_47[6]}
   );
   gpc1_1 gpc4298 (
      {stage3_47[15]},
      {stage4_47[7]}
   );
   gpc1_1 gpc4299 (
      {stage3_47[16]},
      {stage4_47[8]}
   );
   gpc1_1 gpc4300 (
      {stage3_47[17]},
      {stage4_47[9]}
   );
   gpc1_1 gpc4301 (
      {stage3_47[18]},
      {stage4_47[10]}
   );
   gpc1_1 gpc4302 (
      {stage3_47[19]},
      {stage4_47[11]}
   );
   gpc1_1 gpc4303 (
      {stage3_47[20]},
      {stage4_47[12]}
   );
   gpc1_1 gpc4304 (
      {stage3_47[21]},
      {stage4_47[13]}
   );
   gpc1_1 gpc4305 (
      {stage3_47[22]},
      {stage4_47[14]}
   );
   gpc1_1 gpc4306 (
      {stage3_47[23]},
      {stage4_47[15]}
   );
   gpc1_1 gpc4307 (
      {stage3_48[8]},
      {stage4_48[4]}
   );
   gpc1_1 gpc4308 (
      {stage3_48[9]},
      {stage4_48[5]}
   );
   gpc1_1 gpc4309 (
      {stage3_48[10]},
      {stage4_48[6]}
   );
   gpc1_1 gpc4310 (
      {stage3_48[11]},
      {stage4_48[7]}
   );
   gpc1_1 gpc4311 (
      {stage3_48[12]},
      {stage4_48[8]}
   );
   gpc1_1 gpc4312 (
      {stage3_48[13]},
      {stage4_48[9]}
   );
   gpc1_1 gpc4313 (
      {stage3_48[14]},
      {stage4_48[10]}
   );
   gpc1_1 gpc4314 (
      {stage3_48[15]},
      {stage4_48[11]}
   );
   gpc1_1 gpc4315 (
      {stage3_49[6]},
      {stage4_49[5]}
   );
   gpc1_1 gpc4316 (
      {stage3_49[7]},
      {stage4_49[6]}
   );
   gpc1_1 gpc4317 (
      {stage3_49[8]},
      {stage4_49[7]}
   );
   gpc1_1 gpc4318 (
      {stage3_49[9]},
      {stage4_49[8]}
   );
   gpc1_1 gpc4319 (
      {stage3_49[10]},
      {stage4_49[9]}
   );
   gpc1_1 gpc4320 (
      {stage3_49[11]},
      {stage4_49[10]}
   );
   gpc1_1 gpc4321 (
      {stage3_49[12]},
      {stage4_49[11]}
   );
   gpc1_1 gpc4322 (
      {stage3_49[13]},
      {stage4_49[12]}
   );
   gpc1_1 gpc4323 (
      {stage3_50[31]},
      {stage4_50[6]}
   );
   gpc1_1 gpc4324 (
      {stage3_51[12]},
      {stage4_51[7]}
   );
   gpc1_1 gpc4325 (
      {stage3_51[13]},
      {stage4_51[8]}
   );
   gpc1_1 gpc4326 (
      {stage3_52[23]},
      {stage4_52[8]}
   );
   gpc1_1 gpc4327 (
      {stage3_53[7]},
      {stage4_53[6]}
   );
   gpc1_1 gpc4328 (
      {stage3_53[8]},
      {stage4_53[7]}
   );
   gpc1_1 gpc4329 (
      {stage3_53[9]},
      {stage4_53[8]}
   );
   gpc1_1 gpc4330 (
      {stage3_53[10]},
      {stage4_53[9]}
   );
   gpc1_1 gpc4331 (
      {stage3_53[11]},
      {stage4_53[10]}
   );
   gpc1_1 gpc4332 (
      {stage3_53[12]},
      {stage4_53[11]}
   );
   gpc1_1 gpc4333 (
      {stage3_53[13]},
      {stage4_53[12]}
   );
   gpc1_1 gpc4334 (
      {stage3_53[14]},
      {stage4_53[13]}
   );
   gpc1_1 gpc4335 (
      {stage3_53[15]},
      {stage4_53[14]}
   );
   gpc1_1 gpc4336 (
      {stage3_54[12]},
      {stage4_54[6]}
   );
   gpc1_1 gpc4337 (
      {stage3_54[13]},
      {stage4_54[7]}
   );
   gpc1_1 gpc4338 (
      {stage3_54[14]},
      {stage4_54[8]}
   );
   gpc1_1 gpc4339 (
      {stage3_54[15]},
      {stage4_54[9]}
   );
   gpc1_1 gpc4340 (
      {stage3_55[5]},
      {stage4_55[4]}
   );
   gpc1_1 gpc4341 (
      {stage3_55[6]},
      {stage4_55[5]}
   );
   gpc1_1 gpc4342 (
      {stage3_55[7]},
      {stage4_55[6]}
   );
   gpc1_1 gpc4343 (
      {stage3_55[8]},
      {stage4_55[7]}
   );
   gpc1_1 gpc4344 (
      {stage3_55[9]},
      {stage4_55[8]}
   );
   gpc1_1 gpc4345 (
      {stage3_55[10]},
      {stage4_55[9]}
   );
   gpc1_1 gpc4346 (
      {stage3_55[11]},
      {stage4_55[10]}
   );
   gpc1_1 gpc4347 (
      {stage3_55[12]},
      {stage4_55[11]}
   );
   gpc1_1 gpc4348 (
      {stage3_55[13]},
      {stage4_55[12]}
   );
   gpc1_1 gpc4349 (
      {stage3_55[14]},
      {stage4_55[13]}
   );
   gpc1_1 gpc4350 (
      {stage3_55[15]},
      {stage4_55[14]}
   );
   gpc1_1 gpc4351 (
      {stage3_55[16]},
      {stage4_55[15]}
   );
   gpc1_1 gpc4352 (
      {stage3_55[17]},
      {stage4_55[16]}
   );
   gpc1_1 gpc4353 (
      {stage3_56[24]},
      {stage4_56[6]}
   );
   gpc1_1 gpc4354 (
      {stage3_56[25]},
      {stage4_56[7]}
   );
   gpc1_1 gpc4355 (
      {stage3_56[26]},
      {stage4_56[8]}
   );
   gpc1_1 gpc4356 (
      {stage3_56[27]},
      {stage4_56[9]}
   );
   gpc1_1 gpc4357 (
      {stage3_56[28]},
      {stage4_56[10]}
   );
   gpc1_1 gpc4358 (
      {stage3_56[29]},
      {stage4_56[11]}
   );
   gpc1_1 gpc4359 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc4360 (
      {stage3_58[18]},
      {stage4_58[6]}
   );
   gpc1_1 gpc4361 (
      {stage3_58[19]},
      {stage4_58[7]}
   );
   gpc1_1 gpc4362 (
      {stage3_58[20]},
      {stage4_58[8]}
   );
   gpc1_1 gpc4363 (
      {stage3_58[21]},
      {stage4_58[9]}
   );
   gpc1_1 gpc4364 (
      {stage3_58[22]},
      {stage4_58[10]}
   );
   gpc1_1 gpc4365 (
      {stage3_58[23]},
      {stage4_58[11]}
   );
   gpc1_1 gpc4366 (
      {stage3_58[24]},
      {stage4_58[12]}
   );
   gpc1_1 gpc4367 (
      {stage3_58[25]},
      {stage4_58[13]}
   );
   gpc1_1 gpc4368 (
      {stage3_58[26]},
      {stage4_58[14]}
   );
   gpc1_1 gpc4369 (
      {stage3_58[27]},
      {stage4_58[15]}
   );
   gpc1_1 gpc4370 (
      {stage3_58[28]},
      {stage4_58[16]}
   );
   gpc1_1 gpc4371 (
      {stage3_58[29]},
      {stage4_58[17]}
   );
   gpc1_1 gpc4372 (
      {stage3_58[30]},
      {stage4_58[18]}
   );
   gpc1_1 gpc4373 (
      {stage3_58[31]},
      {stage4_58[19]}
   );
   gpc1_1 gpc4374 (
      {stage3_58[32]},
      {stage4_58[20]}
   );
   gpc1_1 gpc4375 (
      {stage3_59[18]},
      {stage4_59[7]}
   );
   gpc1_1 gpc4376 (
      {stage3_59[19]},
      {stage4_59[8]}
   );
   gpc1_1 gpc4377 (
      {stage3_59[20]},
      {stage4_59[9]}
   );
   gpc1_1 gpc4378 (
      {stage3_59[21]},
      {stage4_59[10]}
   );
   gpc1_1 gpc4379 (
      {stage3_59[22]},
      {stage4_59[11]}
   );
   gpc1_1 gpc4380 (
      {stage3_59[23]},
      {stage4_59[12]}
   );
   gpc1_1 gpc4381 (
      {stage3_59[24]},
      {stage4_59[13]}
   );
   gpc1_1 gpc4382 (
      {stage3_59[25]},
      {stage4_59[14]}
   );
   gpc1_1 gpc4383 (
      {stage3_59[26]},
      {stage4_59[15]}
   );
   gpc1_1 gpc4384 (
      {stage3_59[27]},
      {stage4_59[16]}
   );
   gpc1_1 gpc4385 (
      {stage3_60[6]},
      {stage4_60[7]}
   );
   gpc1_1 gpc4386 (
      {stage3_60[7]},
      {stage4_60[8]}
   );
   gpc1_1 gpc4387 (
      {stage3_60[8]},
      {stage4_60[9]}
   );
   gpc1_1 gpc4388 (
      {stage3_60[9]},
      {stage4_60[10]}
   );
   gpc1_1 gpc4389 (
      {stage3_60[10]},
      {stage4_60[11]}
   );
   gpc1_1 gpc4390 (
      {stage3_60[11]},
      {stage4_60[12]}
   );
   gpc1_1 gpc4391 (
      {stage3_60[12]},
      {stage4_60[13]}
   );
   gpc1_1 gpc4392 (
      {stage3_60[13]},
      {stage4_60[14]}
   );
   gpc1_1 gpc4393 (
      {stage3_60[14]},
      {stage4_60[15]}
   );
   gpc1_1 gpc4394 (
      {stage3_61[12]},
      {stage4_61[4]}
   );
   gpc1_1 gpc4395 (
      {stage3_61[13]},
      {stage4_61[5]}
   );
   gpc1_1 gpc4396 (
      {stage3_61[14]},
      {stage4_61[6]}
   );
   gpc1_1 gpc4397 (
      {stage3_61[15]},
      {stage4_61[7]}
   );
   gpc1_1 gpc4398 (
      {stage3_61[16]},
      {stage4_61[8]}
   );
   gpc1_1 gpc4399 (
      {stage3_61[17]},
      {stage4_61[9]}
   );
   gpc1_1 gpc4400 (
      {stage3_61[18]},
      {stage4_61[10]}
   );
   gpc1_1 gpc4401 (
      {stage3_61[19]},
      {stage4_61[11]}
   );
   gpc1_1 gpc4402 (
      {stage3_61[20]},
      {stage4_61[12]}
   );
   gpc1_1 gpc4403 (
      {stage3_61[21]},
      {stage4_61[13]}
   );
   gpc1_1 gpc4404 (
      {stage3_61[22]},
      {stage4_61[14]}
   );
   gpc1_1 gpc4405 (
      {stage3_61[23]},
      {stage4_61[15]}
   );
   gpc1_1 gpc4406 (
      {stage3_61[24]},
      {stage4_61[16]}
   );
   gpc1_1 gpc4407 (
      {stage3_62[18]},
      {stage4_62[5]}
   );
   gpc1_1 gpc4408 (
      {stage3_62[19]},
      {stage4_62[6]}
   );
   gpc1_1 gpc4409 (
      {stage3_62[20]},
      {stage4_62[7]}
   );
   gpc1_1 gpc4410 (
      {stage3_63[12]},
      {stage4_63[7]}
   );
   gpc1_1 gpc4411 (
      {stage3_63[13]},
      {stage4_63[8]}
   );
   gpc1_1 gpc4412 (
      {stage3_63[14]},
      {stage4_63[9]}
   );
   gpc1_1 gpc4413 (
      {stage3_63[15]},
      {stage4_63[10]}
   );
   gpc1_1 gpc4414 (
      {stage3_63[16]},
      {stage4_63[11]}
   );
   gpc1_1 gpc4415 (
      {stage3_63[17]},
      {stage4_63[12]}
   );
   gpc1_1 gpc4416 (
      {stage3_64[12]},
      {stage4_64[5]}
   );
   gpc1_1 gpc4417 (
      {stage3_64[13]},
      {stage4_64[6]}
   );
   gpc1_1 gpc4418 (
      {stage3_64[14]},
      {stage4_64[7]}
   );
   gpc1_1 gpc4419 (
      {stage3_64[15]},
      {stage4_64[8]}
   );
   gpc1_1 gpc4420 (
      {stage3_64[16]},
      {stage4_64[9]}
   );
   gpc1_1 gpc4421 (
      {stage3_64[17]},
      {stage4_64[10]}
   );
   gpc1_1 gpc4422 (
      {stage3_64[18]},
      {stage4_64[11]}
   );
   gpc1_1 gpc4423 (
      {stage3_64[19]},
      {stage4_64[12]}
   );
   gpc1_1 gpc4424 (
      {stage3_64[20]},
      {stage4_64[13]}
   );
   gpc1_1 gpc4425 (
      {stage3_64[21]},
      {stage4_64[14]}
   );
   gpc1_1 gpc4426 (
      {stage3_64[22]},
      {stage4_64[15]}
   );
   gpc1_1 gpc4427 (
      {stage3_64[23]},
      {stage4_64[16]}
   );
   gpc1_1 gpc4428 (
      {stage3_64[24]},
      {stage4_64[17]}
   );
   gpc1_1 gpc4429 (
      {stage3_64[25]},
      {stage4_64[18]}
   );
   gpc1_1 gpc4430 (
      {stage3_64[26]},
      {stage4_64[19]}
   );
   gpc1_1 gpc4431 (
      {stage3_64[27]},
      {stage4_64[20]}
   );
   gpc1_1 gpc4432 (
      {stage3_64[28]},
      {stage4_64[21]}
   );
   gpc1_1 gpc4433 (
      {stage3_65[12]},
      {stage4_65[4]}
   );
   gpc1_1 gpc4434 (
      {stage3_65[13]},
      {stage4_65[5]}
   );
   gpc1_1 gpc4435 (
      {stage3_66[0]},
      {stage4_66[4]}
   );
   gpc1_1 gpc4436 (
      {stage3_66[1]},
      {stage4_66[5]}
   );
   gpc1_1 gpc4437 (
      {stage3_66[2]},
      {stage4_66[6]}
   );
   gpc1_1 gpc4438 (
      {stage3_66[3]},
      {stage4_66[7]}
   );
   gpc1_1 gpc4439 (
      {stage3_66[4]},
      {stage4_66[8]}
   );
   gpc1_1 gpc4440 (
      {stage3_66[5]},
      {stage4_66[9]}
   );
   gpc1_1 gpc4441 (
      {stage3_66[6]},
      {stage4_66[10]}
   );
   gpc1_1 gpc4442 (
      {stage3_66[7]},
      {stage4_66[11]}
   );
   gpc1_1 gpc4443 (
      {stage3_66[8]},
      {stage4_66[12]}
   );
   gpc1_1 gpc4444 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc1_1 gpc4445 (
      {stage3_67[1]},
      {stage4_67[3]}
   );
   gpc1_1 gpc4446 (
      {stage3_67[2]},
      {stage4_67[4]}
   );
   gpc1_1 gpc4447 (
      {stage3_67[3]},
      {stage4_67[5]}
   );
   gpc1_1 gpc4448 (
      {stage3_67[4]},
      {stage4_67[6]}
   );
   gpc1_1 gpc4449 (
      {stage3_68[0]},
      {stage4_68[0]}
   );
   gpc1_1 gpc4450 (
      {stage3_68[1]},
      {stage4_68[1]}
   );
   gpc1343_5 gpc4451 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3]},
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc4452 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc606_5 gpc4453 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc4454 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[2]}
   );
   gpc606_5 gpc4455 (
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1],stage5_9[2]}
   );
   gpc606_5 gpc4456 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc615_5 gpc4457 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4]},
      {stage4_15[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc615_5 gpc4458 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[6]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[2],stage5_16[2],stage5_15[2]}
   );
   gpc606_5 gpc4459 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[3]}
   );
   gpc606_5 gpc4460 (
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], 1'b0},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[4]}
   );
   gpc615_5 gpc4461 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[12]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[2],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc606_5 gpc4462 (
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[1],stage5_21[3],stage5_20[3]}
   );
   gpc7_3 gpc4463 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[2],stage5_21[4]}
   );
   gpc606_5 gpc4464 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[2]}
   );
   gpc1406_5 gpc4465 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[2]}
   );
   gpc1406_5 gpc4466 (
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage4_27[1]},
      {stage5_28[1],stage5_27[2],stage5_26[2],stage5_25[2],stage5_24[3]}
   );
   gpc615_5 gpc4467 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[2],stage5_27[3]}
   );
   gpc2135_5 gpc4468 (
      {stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage4_29[6], stage4_29[7], stage4_29[8]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[1],stage5_28[3]}
   );
   gpc606_5 gpc4469 (
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[2],stage5_28[4]}
   );
   gpc615_5 gpc4470 (
      {stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[2],stage5_31[3],stage5_30[3]}
   );
   gpc615_5 gpc4471 (
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], 1'b0},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[3],stage5_31[4],stage5_30[4]}
   );
   gpc615_5 gpc4472 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[12]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[2],stage5_33[2],stage5_32[4],stage5_31[5]}
   );
   gpc1343_5 gpc4473 (
      {stage4_33[6], stage4_33[7], stage4_33[8]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[3],stage5_33[3]}
   );
   gpc1343_5 gpc4474 (
      {stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_34[4], stage4_34[5], stage4_34[6], stage4_34[7]},
      {stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage4_36[1]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[4],stage5_33[4]}
   );
   gpc615_5 gpc4475 (
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10]},
      {stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3]}
   );
   gpc606_5 gpc4476 (
      {stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[1],stage5_38[1],stage5_37[3],stage5_36[3]}
   );
   gpc207_4 gpc4477 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_41[0], stage4_41[1]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[2]}
   );
   gpc606_5 gpc4478 (
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1],stage5_40[2]}
   );
   gpc606_5 gpc4479 (
      {stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[1],stage5_42[2],stage5_41[2],stage5_40[3]}
   );
   gpc606_5 gpc4480 (
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[2],stage5_42[3],stage5_41[3]}
   );
   gpc615_5 gpc4481 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[3],stage5_43[3],stage5_42[4]}
   );
   gpc606_5 gpc4482 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[4]}
   );
   gpc23_3 gpc4483 (
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[6], stage4_46[7]},
      {stage5_47[1],stage5_46[2],stage5_45[3]}
   );
   gpc606_5 gpc4484 (
      {stage4_45[3], stage4_45[4], stage4_45[5], stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[1],stage5_47[2],stage5_46[3],stage5_45[4]}
   );
   gpc615_5 gpc4485 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[2],stage5_47[3],stage5_46[4]}
   );
   gpc615_5 gpc4486 (
      {stage4_46[13], stage4_46[14], stage4_46[15], stage4_46[16], stage4_46[17]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[3],stage5_47[4],stage5_46[5]}
   );
   gpc135_4 gpc4487 (
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4]},
      {stage4_50[0], stage4_50[1], stage4_50[2]},
      {stage4_51[0]},
      {stage5_52[0],stage5_51[0],stage5_50[2],stage5_49[3]}
   );
   gpc606_5 gpc4488 (
      {stage4_49[5], stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10]},
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage5_53[0],stage5_52[1],stage5_51[1],stage5_50[3],stage5_49[4]}
   );
   gpc615_5 gpc4489 (
      {stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6], 1'b0},
      {stage4_51[7]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[1],stage5_52[2],stage5_51[2],stage5_50[4]}
   );
   gpc606_5 gpc4490 (
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[0],stage5_54[1],stage5_53[2]}
   );
   gpc606_5 gpc4491 (
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[1],stage5_54[2],stage5_53[3]}
   );
   gpc615_5 gpc4492 (
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4]},
      {stage4_55[12]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[2],stage5_54[3]}
   );
   gpc606_5 gpc4493 (
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[3],stage5_56[3]}
   );
   gpc1343_5 gpc4494 (
      {stage4_57[0], stage4_57[1], stage4_57[2]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9]},
      {stage4_59[0], stage4_59[1], stage4_59[2]},
      {stage4_60[0]},
      {stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[2],stage5_57[4]}
   );
   gpc1343_5 gpc4495 (
      {stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage4_58[10], stage4_58[11], stage4_58[12], stage4_58[13]},
      {stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[1]},
      {stage5_61[1],stage5_60[2],stage5_59[2],stage5_58[3],stage5_57[5]}
   );
   gpc606_5 gpc4496 (
      {stage4_58[14], stage4_58[15], stage4_58[16], stage4_58[17], stage4_58[18], stage4_58[19]},
      {stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5], stage4_60[6], stage4_60[7]},
      {stage5_62[0],stage5_61[2],stage5_60[3],stage5_59[3],stage5_58[4]}
   );
   gpc606_5 gpc4497 (
      {stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[3],stage5_60[4],stage5_59[4]}
   );
   gpc606_5 gpc4498 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16], 1'b0},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[4],stage5_60[5],stage5_59[5]}
   );
   gpc606_5 gpc4499 (
      {stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[3],stage5_61[5],stage5_60[6]}
   );
   gpc135_4 gpc4500 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4]},
      {stage4_64[0], stage4_64[1], stage4_64[2]},
      {stage4_65[0]},
      {stage5_66[0],stage5_65[0],stage5_64[1],stage5_63[3]}
   );
   gpc606_5 gpc4501 (
      {stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6], stage4_64[7], stage4_64[8]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], stage4_66[5]},
      {stage5_68[0],stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[2]}
   );
   gpc606_5 gpc4502 (
      {stage4_64[9], stage4_64[10], stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14]},
      {stage4_66[6], stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], stage4_66[11]},
      {stage5_68[1],stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[3]}
   );
   gpc606_5 gpc4503 (
      {stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5], 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage5_69[0],stage5_68[2],stage5_67[2],stage5_66[3],stage5_65[3]}
   );
   gpc1_1 gpc4504 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4505 (
      {stage4_2[3]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4506 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4507 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4508 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4509 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc4510 (
      {stage4_3[2]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4511 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4512 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4513 (
      {stage4_4[6]},
      {stage5_4[2]}
   );
   gpc1_1 gpc4514 (
      {stage4_4[7]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4515 (
      {stage4_4[8]},
      {stage5_4[4]}
   );
   gpc1_1 gpc4516 (
      {stage4_5[6]},
      {stage5_5[2]}
   );
   gpc1_1 gpc4517 (
      {stage4_5[7]},
      {stage5_5[3]}
   );
   gpc1_1 gpc4518 (
      {stage4_5[8]},
      {stage5_5[4]}
   );
   gpc1_1 gpc4519 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc4520 (
      {stage4_6[7]},
      {stage5_6[3]}
   );
   gpc1_1 gpc4521 (
      {stage4_6[8]},
      {stage5_6[4]}
   );
   gpc1_1 gpc4522 (
      {stage4_6[9]},
      {stage5_6[5]}
   );
   gpc1_1 gpc4523 (
      {stage4_6[10]},
      {stage5_6[6]}
   );
   gpc1_1 gpc4524 (
      {stage4_6[11]},
      {stage5_6[7]}
   );
   gpc1_1 gpc4525 (
      {stage4_6[12]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4526 (
      {stage4_6[13]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4527 (
      {stage4_7[6]},
      {stage5_7[2]}
   );
   gpc1_1 gpc4528 (
      {stage4_7[7]},
      {stage5_7[3]}
   );
   gpc1_1 gpc4529 (
      {stage4_8[5]},
      {stage5_8[3]}
   );
   gpc1_1 gpc4530 (
      {stage4_8[6]},
      {stage5_8[4]}
   );
   gpc1_1 gpc4531 (
      {stage4_8[7]},
      {stage5_8[5]}
   );
   gpc1_1 gpc4532 (
      {stage4_8[8]},
      {stage5_8[6]}
   );
   gpc1_1 gpc4533 (
      {stage4_8[9]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4534 (
      {stage4_10[6]},
      {stage5_10[2]}
   );
   gpc1_1 gpc4535 (
      {stage4_10[7]},
      {stage5_10[3]}
   );
   gpc1_1 gpc4536 (
      {stage4_10[8]},
      {stage5_10[4]}
   );
   gpc1_1 gpc4537 (
      {stage4_11[6]},
      {stage5_11[2]}
   );
   gpc1_1 gpc4538 (
      {stage4_12[0]},
      {stage5_12[2]}
   );
   gpc1_1 gpc4539 (
      {stage4_12[1]},
      {stage5_12[3]}
   );
   gpc1_1 gpc4540 (
      {stage4_12[2]},
      {stage5_12[4]}
   );
   gpc1_1 gpc4541 (
      {stage4_12[3]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4542 (
      {stage4_12[4]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4543 (
      {stage4_12[5]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4544 (
      {stage4_12[6]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4545 (
      {stage4_12[7]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4546 (
      {stage4_12[8]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4547 (
      {stage4_13[6]},
      {stage5_13[2]}
   );
   gpc1_1 gpc4548 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc4549 (
      {stage4_13[8]},
      {stage5_13[4]}
   );
   gpc1_1 gpc4550 (
      {stage4_13[9]},
      {stage5_13[5]}
   );
   gpc1_1 gpc4551 (
      {stage4_14[5]},
      {stage5_14[2]}
   );
   gpc1_1 gpc4552 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc4553 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc4554 (
      {stage4_14[8]},
      {stage5_14[5]}
   );
   gpc1_1 gpc4555 (
      {stage4_14[9]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4556 (
      {stage4_14[10]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4557 (
      {stage4_15[12]},
      {stage5_15[3]}
   );
   gpc1_1 gpc4558 (
      {stage4_15[13]},
      {stage5_15[4]}
   );
   gpc1_1 gpc4559 (
      {stage4_15[14]},
      {stage5_15[5]}
   );
   gpc1_1 gpc4560 (
      {stage4_15[15]},
      {stage5_15[6]}
   );
   gpc1_1 gpc4561 (
      {stage4_15[16]},
      {stage5_15[7]}
   );
   gpc1_1 gpc4562 (
      {stage4_16[7]},
      {stage5_16[3]}
   );
   gpc1_1 gpc4563 (
      {stage4_16[8]},
      {stage5_16[4]}
   );
   gpc1_1 gpc4564 (
      {stage4_16[9]},
      {stage5_16[5]}
   );
   gpc1_1 gpc4565 (
      {stage4_16[10]},
      {stage5_16[6]}
   );
   gpc1_1 gpc4566 (
      {stage4_16[11]},
      {stage5_16[7]}
   );
   gpc1_1 gpc4567 (
      {stage4_16[12]},
      {stage5_16[8]}
   );
   gpc1_1 gpc4568 (
      {stage4_18[5]},
      {stage5_18[5]}
   );
   gpc1_1 gpc4569 (
      {stage4_19[13]},
      {stage5_19[4]}
   );
   gpc1_1 gpc4570 (
      {stage4_19[14]},
      {stage5_19[5]}
   );
   gpc1_1 gpc4571 (
      {stage4_19[15]},
      {stage5_19[6]}
   );
   gpc1_1 gpc4572 (
      {stage4_21[7]},
      {stage5_21[5]}
   );
   gpc1_1 gpc4573 (
      {stage4_22[6]},
      {stage5_22[3]}
   );
   gpc1_1 gpc4574 (
      {stage4_22[7]},
      {stage5_22[4]}
   );
   gpc1_1 gpc4575 (
      {stage4_22[8]},
      {stage5_22[5]}
   );
   gpc1_1 gpc4576 (
      {stage4_22[9]},
      {stage5_22[6]}
   );
   gpc1_1 gpc4577 (
      {stage4_22[10]},
      {stage5_22[7]}
   );
   gpc1_1 gpc4578 (
      {stage4_22[11]},
      {stage5_22[8]}
   );
   gpc1_1 gpc4579 (
      {stage4_22[12]},
      {stage5_22[9]}
   );
   gpc1_1 gpc4580 (
      {stage4_22[13]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4581 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc4582 (
      {stage4_23[7]},
      {stage5_23[4]}
   );
   gpc1_1 gpc4583 (
      {stage4_23[8]},
      {stage5_23[5]}
   );
   gpc1_1 gpc4584 (
      {stage4_23[9]},
      {stage5_23[6]}
   );
   gpc1_1 gpc4585 (
      {stage4_24[12]},
      {stage5_24[4]}
   );
   gpc1_1 gpc4586 (
      {stage4_24[13]},
      {stage5_24[5]}
   );
   gpc1_1 gpc4587 (
      {stage4_24[14]},
      {stage5_24[6]}
   );
   gpc1_1 gpc4588 (
      {stage4_24[15]},
      {stage5_24[7]}
   );
   gpc1_1 gpc4589 (
      {stage4_24[16]},
      {stage5_24[8]}
   );
   gpc1_1 gpc4590 (
      {stage4_24[17]},
      {stage5_24[9]}
   );
   gpc1_1 gpc4591 (
      {stage4_29[9]},
      {stage5_29[3]}
   );
   gpc1_1 gpc4592 (
      {stage4_32[13]},
      {stage5_32[5]}
   );
   gpc1_1 gpc4593 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4594 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4595 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4596 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4597 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4598 (
      {stage4_32[19]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4599 (
      {stage4_34[8]},
      {stage5_34[5]}
   );
   gpc1_1 gpc4600 (
      {stage4_34[9]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4601 (
      {stage4_34[10]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4602 (
      {stage4_36[9]},
      {stage5_36[4]}
   );
   gpc1_1 gpc4603 (
      {stage4_39[7]},
      {stage5_39[3]}
   );
   gpc1_1 gpc4604 (
      {stage4_39[8]},
      {stage5_39[4]}
   );
   gpc1_1 gpc4605 (
      {stage4_39[9]},
      {stage5_39[5]}
   );
   gpc1_1 gpc4606 (
      {stage4_40[12]},
      {stage5_40[4]}
   );
   gpc1_1 gpc4607 (
      {stage4_40[13]},
      {stage5_40[5]}
   );
   gpc1_1 gpc4608 (
      {stage4_41[8]},
      {stage5_41[4]}
   );
   gpc1_1 gpc4609 (
      {stage4_41[9]},
      {stage5_41[5]}
   );
   gpc1_1 gpc4610 (
      {stage4_41[10]},
      {stage5_41[6]}
   );
   gpc1_1 gpc4611 (
      {stage4_41[11]},
      {stage5_41[7]}
   );
   gpc1_1 gpc4612 (
      {stage4_41[12]},
      {stage5_41[8]}
   );
   gpc1_1 gpc4613 (
      {stage4_41[13]},
      {stage5_41[9]}
   );
   gpc1_1 gpc4614 (
      {stage4_41[14]},
      {stage5_41[10]}
   );
   gpc1_1 gpc4615 (
      {stage4_41[15]},
      {stage5_41[11]}
   );
   gpc1_1 gpc4616 (
      {stage4_41[16]},
      {stage5_41[12]}
   );
   gpc1_1 gpc4617 (
      {stage4_44[12]},
      {stage5_44[5]}
   );
   gpc1_1 gpc4618 (
      {stage4_47[8]},
      {stage5_47[5]}
   );
   gpc1_1 gpc4619 (
      {stage4_47[9]},
      {stage5_47[6]}
   );
   gpc1_1 gpc4620 (
      {stage4_47[10]},
      {stage5_47[7]}
   );
   gpc1_1 gpc4621 (
      {stage4_47[11]},
      {stage5_47[8]}
   );
   gpc1_1 gpc4622 (
      {stage4_47[12]},
      {stage5_47[9]}
   );
   gpc1_1 gpc4623 (
      {stage4_47[13]},
      {stage5_47[10]}
   );
   gpc1_1 gpc4624 (
      {stage4_47[14]},
      {stage5_47[11]}
   );
   gpc1_1 gpc4625 (
      {stage4_47[15]},
      {stage5_47[12]}
   );
   gpc1_1 gpc4626 (
      {stage4_49[11]},
      {stage5_49[5]}
   );
   gpc1_1 gpc4627 (
      {stage4_49[12]},
      {stage5_49[6]}
   );
   gpc1_1 gpc4628 (
      {stage4_51[8]},
      {stage5_51[3]}
   );
   gpc1_1 gpc4629 (
      {stage4_52[6]},
      {stage5_52[3]}
   );
   gpc1_1 gpc4630 (
      {stage4_52[7]},
      {stage5_52[4]}
   );
   gpc1_1 gpc4631 (
      {stage4_52[8]},
      {stage5_52[5]}
   );
   gpc1_1 gpc4632 (
      {stage4_53[12]},
      {stage5_53[4]}
   );
   gpc1_1 gpc4633 (
      {stage4_53[13]},
      {stage5_53[5]}
   );
   gpc1_1 gpc4634 (
      {stage4_53[14]},
      {stage5_53[6]}
   );
   gpc1_1 gpc4635 (
      {stage4_54[5]},
      {stage5_54[4]}
   );
   gpc1_1 gpc4636 (
      {stage4_54[6]},
      {stage5_54[5]}
   );
   gpc1_1 gpc4637 (
      {stage4_54[7]},
      {stage5_54[6]}
   );
   gpc1_1 gpc4638 (
      {stage4_54[8]},
      {stage5_54[7]}
   );
   gpc1_1 gpc4639 (
      {stage4_54[9]},
      {stage5_54[8]}
   );
   gpc1_1 gpc4640 (
      {stage4_55[13]},
      {stage5_55[3]}
   );
   gpc1_1 gpc4641 (
      {stage4_55[14]},
      {stage5_55[4]}
   );
   gpc1_1 gpc4642 (
      {stage4_55[15]},
      {stage5_55[5]}
   );
   gpc1_1 gpc4643 (
      {stage4_55[16]},
      {stage5_55[6]}
   );
   gpc1_1 gpc4644 (
      {stage4_56[12]},
      {stage5_56[4]}
   );
   gpc1_1 gpc4645 (
      {stage4_58[20]},
      {stage5_58[5]}
   );
   gpc1_1 gpc4646 (
      {stage4_60[14]},
      {stage5_60[7]}
   );
   gpc1_1 gpc4647 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc4648 (
      {stage4_61[12]},
      {stage5_61[6]}
   );
   gpc1_1 gpc4649 (
      {stage4_61[13]},
      {stage5_61[7]}
   );
   gpc1_1 gpc4650 (
      {stage4_61[14]},
      {stage5_61[8]}
   );
   gpc1_1 gpc4651 (
      {stage4_61[15]},
      {stage5_61[9]}
   );
   gpc1_1 gpc4652 (
      {stage4_61[16]},
      {stage5_61[10]}
   );
   gpc1_1 gpc4653 (
      {stage4_62[6]},
      {stage5_62[4]}
   );
   gpc1_1 gpc4654 (
      {stage4_62[7]},
      {stage5_62[5]}
   );
   gpc1_1 gpc4655 (
      {stage4_63[5]},
      {stage5_63[4]}
   );
   gpc1_1 gpc4656 (
      {stage4_63[6]},
      {stage5_63[5]}
   );
   gpc1_1 gpc4657 (
      {stage4_63[7]},
      {stage5_63[6]}
   );
   gpc1_1 gpc4658 (
      {stage4_63[8]},
      {stage5_63[7]}
   );
   gpc1_1 gpc4659 (
      {stage4_63[9]},
      {stage5_63[8]}
   );
   gpc1_1 gpc4660 (
      {stage4_63[10]},
      {stage5_63[9]}
   );
   gpc1_1 gpc4661 (
      {stage4_63[11]},
      {stage5_63[10]}
   );
   gpc1_1 gpc4662 (
      {stage4_63[12]},
      {stage5_63[11]}
   );
   gpc1_1 gpc4663 (
      {stage4_64[15]},
      {stage5_64[4]}
   );
   gpc1_1 gpc4664 (
      {stage4_64[16]},
      {stage5_64[5]}
   );
   gpc1_1 gpc4665 (
      {stage4_64[17]},
      {stage5_64[6]}
   );
   gpc1_1 gpc4666 (
      {stage4_64[18]},
      {stage5_64[7]}
   );
   gpc1_1 gpc4667 (
      {stage4_64[19]},
      {stage5_64[8]}
   );
   gpc1_1 gpc4668 (
      {stage4_64[20]},
      {stage5_64[9]}
   );
   gpc1_1 gpc4669 (
      {stage4_64[21]},
      {stage5_64[10]}
   );
   gpc1_1 gpc4670 (
      {stage4_66[12]},
      {stage5_66[4]}
   );
   gpc1_1 gpc4671 (
      {stage4_67[6]},
      {stage5_67[3]}
   );
   gpc1_1 gpc4672 (
      {stage4_68[0]},
      {stage5_68[3]}
   );
   gpc1_1 gpc4673 (
      {stage4_68[1]},
      {stage5_68[4]}
   );
   gpc615_5 gpc4674 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], 1'b0},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc1415_5 gpc4675 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1415_5 gpc4676 (
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8], stage5_6[9]},
      {stage5_7[1]},
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2]}
   );
   gpc606_5 gpc4677 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0]}
   );
   gpc606_5 gpc4678 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc4679 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[2]}
   );
   gpc2135_5 gpc4680 (
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[1]}
   );
   gpc1163_5 gpc4681 (
      {stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage5_24[0]},
      {stage5_25[0]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[1],stage6_22[1]}
   );
   gpc615_5 gpc4682 (
      {stage5_22[5], stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9]},
      {stage5_23[6]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[1],stage6_25[1],stage6_24[1],stage6_23[2],stage6_22[2]}
   );
   gpc1343_5 gpc4683 (
      {stage5_24[7], stage5_24[8], stage5_24[9]},
      {stage5_25[1], stage5_25[2], 1'b0, 1'b0},
      {stage5_26[0], stage5_26[1], stage5_26[2]},
      {stage5_27[0]},
      {stage6_28[0],stage6_27[0],stage6_26[2],stage6_25[2],stage6_24[2]}
   );
   gpc3_2 gpc4684 (
      {stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc4685 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], 1'b0},
      {stage6_32[0],stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2]}
   );
   gpc606_5 gpc4686 (
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], 1'b0, 1'b0},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc4687 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1],stage6_32[2]}
   );
   gpc615_5 gpc4688 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4]},
      {stage5_34[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], 1'b0, 1'b0},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc4689 (
      {stage5_38[0], stage5_38[1], 1'b0, 1'b0, 1'b0},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage6_42[0],stage6_41[0],stage6_40[0],stage6_39[0],stage6_38[0]}
   );
   gpc606_5 gpc4690 (
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], 1'b0},
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage6_43[0],stage6_42[1],stage6_41[1],stage6_40[1],stage6_39[1]}
   );
   gpc606_5 gpc4691 (
      {stage5_41[6], stage5_41[7], stage5_41[8], stage5_41[9], stage5_41[10], stage5_41[11]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], 1'b0, 1'b0},
      {stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[2],stage6_41[2]}
   );
   gpc606_5 gpc4692 (
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[0],stage6_45[1],stage6_44[1]}
   );
   gpc606_5 gpc4693 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], 1'b0},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[1],stage6_45[2]}
   );
   gpc615_5 gpc4694 (
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10]},
      {stage5_48[0]},
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage6_51[0],stage6_50[0],stage6_49[1],stage6_48[2],stage6_47[2]}
   );
   gpc1343_5 gpc4695 (
      {stage5_50[0], stage5_50[1], stage5_50[2]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3]},
      {stage5_52[0], stage5_52[1], stage5_52[2]},
      {stage5_53[0]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[1],stage6_50[1]}
   );
   gpc223_4 gpc4696 (
      {stage5_53[1], stage5_53[2], stage5_53[3]},
      {stage5_54[0], stage5_54[1]},
      {stage5_55[0], stage5_55[1]},
      {stage6_56[0],stage6_55[0],stage6_54[1],stage6_53[1]}
   );
   gpc207_4 gpc4697 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6], stage5_54[7], stage5_54[8]},
      {stage5_56[0], stage5_56[1]},
      {stage6_57[0],stage6_56[1],stage6_55[1],stage6_54[2]}
   );
   gpc615_5 gpc4698 (
      {stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[2]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[1],stage6_56[2],stage6_55[2]}
   );
   gpc606_5 gpc4699 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1]}
   );
   gpc606_5 gpc4700 (
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_61[0], stage5_61[1], stage5_61[2], stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage6_63[0],stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[2]}
   );
   gpc606_5 gpc4701 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], 1'b0},
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage6_65[0],stage6_64[0],stage6_63[1],stage6_62[2],stage6_61[2]}
   );
   gpc606_5 gpc4702 (
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage6_66[0],stage6_65[1],stage6_64[1],stage6_63[2],stage6_62[3]}
   );
   gpc606_5 gpc4703 (
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], stage5_63[11]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], 1'b0, 1'b0},
      {stage6_67[0],stage6_66[1],stage6_65[2],stage6_64[2],stage6_63[3]}
   );
   gpc606_5 gpc4704 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], 1'b0},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], 1'b0},
      {stage6_68[0],stage6_67[1],stage6_66[2],stage6_65[3],stage6_64[3]}
   );
   gpc1_1 gpc4705 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4706 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4707 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc4708 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc4709 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc4710 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc4711 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc4712 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc4713 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc4714 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc4715 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc4716 (
      {stage5_4[4]},
      {stage6_4[4]}
   );
   gpc1_1 gpc4717 (
      {stage5_7[2]},
      {stage6_7[3]}
   );
   gpc1_1 gpc4718 (
      {stage5_7[3]},
      {stage6_7[4]}
   );
   gpc1_1 gpc4719 (
      {stage5_9[2]},
      {stage6_9[2]}
   );
   gpc1_1 gpc4720 (
      {stage5_10[0]},
      {stage6_10[2]}
   );
   gpc1_1 gpc4721 (
      {stage5_10[1]},
      {stage6_10[3]}
   );
   gpc1_1 gpc4722 (
      {stage5_10[2]},
      {stage6_10[4]}
   );
   gpc1_1 gpc4723 (
      {stage5_10[3]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4724 (
      {stage5_10[4]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4725 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc4726 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc4727 (
      {stage5_11[2]},
      {stage6_11[2]}
   );
   gpc1_1 gpc4728 (
      {stage5_12[6]},
      {stage6_12[1]}
   );
   gpc1_1 gpc4729 (
      {stage5_12[7]},
      {stage6_12[2]}
   );
   gpc1_1 gpc4730 (
      {stage5_12[8]},
      {stage6_12[3]}
   );
   gpc1_1 gpc4731 (
      {stage5_12[9]},
      {stage6_12[4]}
   );
   gpc1_1 gpc4732 (
      {stage5_12[10]},
      {stage6_12[5]}
   );
   gpc1_1 gpc4733 (
      {stage5_14[6]},
      {stage6_14[2]}
   );
   gpc1_1 gpc4734 (
      {stage5_14[7]},
      {stage6_14[3]}
   );
   gpc1_1 gpc4735 (
      {stage5_15[6]},
      {stage6_15[2]}
   );
   gpc1_1 gpc4736 (
      {stage5_15[7]},
      {stage6_15[3]}
   );
   gpc1_1 gpc4737 (
      {stage5_16[6]},
      {stage6_16[3]}
   );
   gpc1_1 gpc4738 (
      {stage5_16[7]},
      {stage6_16[4]}
   );
   gpc1_1 gpc4739 (
      {stage5_16[8]},
      {stage6_16[5]}
   );
   gpc1_1 gpc4740 (
      {stage5_17[0]},
      {stage6_17[2]}
   );
   gpc1_1 gpc4741 (
      {stage5_17[1]},
      {stage6_17[3]}
   );
   gpc1_1 gpc4742 (
      {stage5_17[2]},
      {stage6_17[4]}
   );
   gpc1_1 gpc4743 (
      {stage5_17[3]},
      {stage6_17[5]}
   );
   gpc1_1 gpc4744 (
      {stage5_17[4]},
      {stage6_17[6]}
   );
   gpc1_1 gpc4745 (
      {stage5_19[5]},
      {stage6_19[2]}
   );
   gpc1_1 gpc4746 (
      {stage5_19[6]},
      {stage6_19[3]}
   );
   gpc1_1 gpc4747 (
      {stage5_20[3]},
      {stage6_20[2]}
   );
   gpc1_1 gpc4748 (
      {stage5_21[1]},
      {stage6_21[1]}
   );
   gpc1_1 gpc4749 (
      {stage5_21[2]},
      {stage6_21[2]}
   );
   gpc1_1 gpc4750 (
      {stage5_21[3]},
      {stage6_21[3]}
   );
   gpc1_1 gpc4751 (
      {stage5_21[4]},
      {stage6_21[4]}
   );
   gpc1_1 gpc4752 (
      {stage5_21[5]},
      {stage6_21[5]}
   );
   gpc1_1 gpc4753 (
      {stage5_22[10]},
      {stage6_22[3]}
   );
   gpc1_1 gpc4754 (
      {stage5_32[6]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4755 (
      {stage5_32[7]},
      {stage6_32[4]}
   );
   gpc1_1 gpc4756 (
      {stage5_32[8]},
      {stage6_32[5]}
   );
   gpc1_1 gpc4757 (
      {stage5_32[9]},
      {stage6_32[6]}
   );
   gpc1_1 gpc4758 (
      {stage5_32[10]},
      {stage6_32[7]}
   );
   gpc1_1 gpc4759 (
      {stage5_32[11]},
      {stage6_32[8]}
   );
   gpc1_1 gpc4760 (
      {stage5_34[7]},
      {stage6_34[2]}
   );
   gpc1_1 gpc4761 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4762 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4763 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4764 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4765 (
      {stage5_36[4]},
      {stage6_36[6]}
   );
   gpc1_1 gpc4766 (
      {stage5_37[0]},
      {stage6_37[1]}
   );
   gpc1_1 gpc4767 (
      {stage5_37[1]},
      {stage6_37[2]}
   );
   gpc1_1 gpc4768 (
      {stage5_37[2]},
      {stage6_37[3]}
   );
   gpc1_1 gpc4769 (
      {stage5_37[3]},
      {stage6_37[4]}
   );
   gpc1_1 gpc4770 (
      {stage5_41[12]},
      {stage6_41[3]}
   );
   gpc1_1 gpc4771 (
      {stage5_42[0]},
      {stage6_42[3]}
   );
   gpc1_1 gpc4772 (
      {stage5_42[1]},
      {stage6_42[4]}
   );
   gpc1_1 gpc4773 (
      {stage5_42[2]},
      {stage6_42[5]}
   );
   gpc1_1 gpc4774 (
      {stage5_42[3]},
      {stage6_42[6]}
   );
   gpc1_1 gpc4775 (
      {stage5_42[4]},
      {stage6_42[7]}
   );
   gpc1_1 gpc4776 (
      {stage5_47[11]},
      {stage6_47[3]}
   );
   gpc1_1 gpc4777 (
      {stage5_47[12]},
      {stage6_47[4]}
   );
   gpc1_1 gpc4778 (
      {stage5_48[1]},
      {stage6_48[3]}
   );
   gpc1_1 gpc4779 (
      {stage5_48[2]},
      {stage6_48[4]}
   );
   gpc1_1 gpc4780 (
      {stage5_48[3]},
      {stage6_48[5]}
   );
   gpc1_1 gpc4781 (
      {stage5_49[6]},
      {stage6_49[2]}
   );
   gpc1_1 gpc4782 (
      {stage5_50[3]},
      {stage6_50[2]}
   );
   gpc1_1 gpc4783 (
      {stage5_50[4]},
      {stage6_50[3]}
   );
   gpc1_1 gpc4784 (
      {stage5_52[3]},
      {stage6_52[1]}
   );
   gpc1_1 gpc4785 (
      {stage5_52[4]},
      {stage6_52[2]}
   );
   gpc1_1 gpc4786 (
      {stage5_52[5]},
      {stage6_52[3]}
   );
   gpc1_1 gpc4787 (
      {stage5_53[4]},
      {stage6_53[2]}
   );
   gpc1_1 gpc4788 (
      {stage5_53[5]},
      {stage6_53[3]}
   );
   gpc1_1 gpc4789 (
      {stage5_53[6]},
      {stage6_53[4]}
   );
   gpc1_1 gpc4790 (
      {stage5_56[3]},
      {stage6_56[3]}
   );
   gpc1_1 gpc4791 (
      {stage5_56[4]},
      {stage6_56[4]}
   );
   gpc1_1 gpc4792 (
      {stage5_60[6]},
      {stage6_60[2]}
   );
   gpc1_1 gpc4793 (
      {stage5_60[7]},
      {stage6_60[3]}
   );
   gpc1_1 gpc4794 (
      {stage5_60[8]},
      {stage6_60[4]}
   );
   gpc1_1 gpc4795 (
      {stage5_67[0]},
      {stage6_67[2]}
   );
   gpc1_1 gpc4796 (
      {stage5_67[1]},
      {stage6_67[3]}
   );
   gpc1_1 gpc4797 (
      {stage5_67[2]},
      {stage6_67[4]}
   );
   gpc1_1 gpc4798 (
      {stage5_67[3]},
      {stage6_67[5]}
   );
   gpc1_1 gpc4799 (
      {stage5_68[0]},
      {stage6_68[1]}
   );
   gpc1_1 gpc4800 (
      {stage5_68[1]},
      {stage6_68[2]}
   );
   gpc1_1 gpc4801 (
      {stage5_68[2]},
      {stage6_68[3]}
   );
   gpc1_1 gpc4802 (
      {stage5_68[3]},
      {stage6_68[4]}
   );
   gpc1_1 gpc4803 (
      {stage5_68[4]},
      {stage6_68[5]}
   );
   gpc1_1 gpc4804 (
      {stage5_69[0]},
      {stage6_69[0]}
   );
   gpc1415_5 gpc4805 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[0]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0]}
   );
   gpc23_3 gpc4806 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc223_4 gpc4807 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[0], stage6_8[1]},
      {stage6_9[0], stage6_9[1]},
      {stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc207_4 gpc4808 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5], stage6_10[6]},
      {stage6_12[0], stage6_12[1]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1]}
   );
   gpc1343_5 gpc4809 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[0], stage6_13[1], 1'b0},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[1],stage7_12[1],stage7_11[1]}
   );
   gpc1343_5 gpc4810 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3]},
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[0],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc4811 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6]},
      {stage6_18[0]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc1343_5 gpc4812 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[0], stage6_20[1], stage6_20[2], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[1]}
   );
   gpc1343_5 gpc4813 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[1], stage6_22[2], stage6_22[3], 1'b0},
      {stage6_23[0], stage6_23[1], stage6_23[2]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[1],stage7_22[1],stage7_21[1]}
   );
   gpc1343_5 gpc4814 (
      {stage6_24[1], stage6_24[2], 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2], 1'b0},
      {stage6_26[0], stage6_26[1], stage6_26[2]},
      {stage6_27[0]},
      {stage7_28[0],stage7_27[0],stage7_26[0],stage7_25[1],stage7_24[1]}
   );
   gpc15_3 gpc4815 (
      {stage6_28[0], stage6_28[1], stage6_28[2], 1'b0, 1'b0},
      {stage6_29[0]},
      {stage7_30[0],stage7_29[0],stage7_28[1]}
   );
   gpc615_5 gpc4816 (
      {stage6_30[0], stage6_30[1], 1'b0, 1'b0, 1'b0},
      {stage6_31[0]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[1]}
   );
   gpc1343_5 gpc4817 (
      {stage6_32[6], stage6_32[7], stage6_32[8]},
      {stage6_33[0], stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[0], stage6_34[1], stage6_34[2]},
      {stage6_35[0]},
      {stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1],stage7_32[1]}
   );
   gpc7_3 gpc4818 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage7_38[0],stage7_37[0],stage7_36[1]}
   );
   gpc2135_5 gpc4819 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4]},
      {stage6_38[0], 1'b0, 1'b0},
      {stage6_39[0]},
      {stage6_40[0], stage6_40[1]},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc135_4 gpc4820 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], 1'b0},
      {stage6_42[0], stage6_42[1], stage6_42[2]},
      {stage6_43[0]},
      {stage7_44[0],stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc4821 (
      {stage6_42[3], stage6_42[4], stage6_42[5], stage6_42[6], stage6_42[7]},
      {stage6_43[1]},
      {stage6_44[0], stage6_44[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[1],stage7_43[1],stage7_42[1]}
   );
   gpc2223_5 gpc4822 (
      {stage6_45[0], stage6_45[1], stage6_45[2]},
      {stage6_46[0], stage6_46[1]},
      {stage6_47[0], stage6_47[1]},
      {stage6_48[0], stage6_48[1]},
      {stage7_49[0],stage7_48[0],stage7_47[0],stage7_46[1],stage7_45[1]}
   );
   gpc1343_5 gpc4823 (
      {stage6_47[2], stage6_47[3], stage6_47[4]},
      {stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5]},
      {stage6_49[0], stage6_49[1], stage6_49[2]},
      {stage6_50[0]},
      {stage7_51[0],stage7_50[0],stage7_49[1],stage7_48[1],stage7_47[1]}
   );
   gpc1343_5 gpc4824 (
      {stage6_50[1], stage6_50[2], stage6_50[3]},
      {stage6_51[0], stage6_51[1], 1'b0, 1'b0},
      {stage6_52[0], stage6_52[1], stage6_52[2]},
      {stage6_53[0]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[1]}
   );
   gpc1343_5 gpc4825 (
      {stage6_52[3], 1'b0, 1'b0},
      {stage6_53[1], stage6_53[2], stage6_53[3], stage6_53[4]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc1163_5 gpc4826 (
      {stage6_55[1], stage6_55[2], 1'b0},
      {stage6_56[0], stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], 1'b0},
      {stage6_57[0]},
      {stage6_58[0]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1343_5 gpc4827 (
      {stage6_59[0], stage6_59[1], stage6_59[2]},
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3]},
      {stage6_61[0], stage6_61[1], stage6_61[2]},
      {stage6_62[0]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[0],stage7_59[1]}
   );
   gpc1343_5 gpc4828 (
      {stage6_62[1], stage6_62[2], stage6_62[3]},
      {stage6_63[0], stage6_63[1], stage6_63[2], stage6_63[3]},
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage6_65[0]},
      {stage7_66[0],stage7_65[0],stage7_64[0],stage7_63[1],stage7_62[1]}
   );
   gpc1343_5 gpc4829 (
      {stage6_65[1], stage6_65[2], stage6_65[3]},
      {stage6_66[0], stage6_66[1], stage6_66[2], 1'b0},
      {stage6_67[0], stage6_67[1], stage6_67[2]},
      {stage6_68[0]},
      {stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[1],stage7_65[1]}
   );
   gpc1163_5 gpc4830 (
      {stage6_67[3], stage6_67[4], stage6_67[5]},
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], 1'b0},
      {stage6_69[0]},
      {1'b0},
      {stage7_71[0],stage7_70[0],stage7_69[1],stage7_68[1],stage7_67[1]}
   );
   gpc1_1 gpc4831 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4832 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4833 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4834 (
      {stage6_4[4]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4835 (
      {stage6_9[2]},
      {stage7_9[1]}
   );
   gpc1_1 gpc4836 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc4837 (
      {stage6_29[1]},
      {stage7_29[1]}
   );
   gpc1_1 gpc4838 (
      {stage6_31[1]},
      {stage7_31[1]}
   );
   gpc1_1 gpc4839 (
      {stage6_35[1]},
      {stage7_35[1]}
   );
   gpc1_1 gpc4840 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc4841 (
      {stage6_57[1]},
      {stage7_57[1]}
   );
   gpc1_1 gpc4842 (
      {stage6_58[1]},
      {stage7_58[1]}
   );
   gpc1_1 gpc4843 (
      {stage6_60[4]},
      {stage7_60[1]}
   );
   gpc1_1 gpc4844 (
      {stage6_64[3]},
      {stage7_64[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [71:0] srcsum;
    wire [71:0] dstsum;
    wire test;
    compressor_CLA162_64 compressor_CLA162_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1b2a43e2d6b9e6fc993be8ddd97ec64fc35b0ad82259d8f65ecbd8ab63ac43ae23c327e8443f91c68fda826e9790ca433cf136806d5af54966f04c747e7ae2d54aac27bc47e976c79f09d40f06ee509bd460ec4d0f86577405e848465701dc3a15fcadb9132e40928ee1c62680c220b7da531aac9aade8cedb7f6f028fd7b2634b54ce1a4111c9ebe6d90ef54e02fcb2fa1b4e89644b37635541bed24837596f847e5b49b2c66242ccccaacdf6f16528e8d084c20bad03dbfa0e8cf1ec6d592ee92bac118a71dd13767a0c64cf02baa413c2ab1d46482e030dd2de43afb498a35228298f69dbc6a9e2949b468a6309424ad72b485b57eea66d3f53c6616f9fdd7ce5522d5ee59ab4a796188e1d0c062fe7c71975094065fdf230311be099cefc8a878f3a74c4c919532011c42930ed72c3c91f63ebbf341423127e963f169c934f9335655a6d82bb935dafb5794696ec51b5753e569b9ad800d9290c56bfcf0b570eb950ede4057c89c905a38cb49dbb9c08686f1511cf6220836459c4961bb5f42e6208a022dba2300d4334b9c810e5c420729833775b764ad71e4d195028d16c7ee26246186c3cbbf59d6254c0f640d47c26e7508baa7433b564122650644d25ea5ec20d6dee8d1ec69ade3caff32a83afc2900b398af2929482bcb3d88f74b1a24cd4b2254df27125f8a6560f30b0bfaf58f9b7866e4d97f8f73d9d08d0d53f80b58dd24db9b1d6cebe38dbcb582120df508775cf4d9eaa3caf4cad79efcfdb9db6fbc4f9af32dc725c8d2e4edbf799d7e24d72b8f4ecff9094ab80502a4242163297694d2e2614586f6fa0eeb58621cea7336765c007bb5e3aa2ab804d1293cd95191059bfa141aedd4817aa5049f7da58e860f254f5977b0ee608c6fe4c0f8e81936125a18c2a56a28f3a6f6fd58792471b3ab66035cc99607f889f6999cff8d0130b98aaa83e68276a9aa56a4856cbda2b35aac359c51bf595fa261595e94699238af510c62978567c40ee5c6d5b44536bbf5eaecb93528573b59e4fcc9ce25763527063358e28174e508e79d7c57f5c74f4ec248855193c4edb195a1e0fa02c2731cd8fc0f7087869606e5f211a13fa0997409be6ac088ca9b9315b7c3ef76f7875eca8b9c0cf7fd11814fc747546632ec2a3a3bf1fed1a1a71ea6f439a1831263e8ac56500185e72841f66ed7dccd13e48bf0e7ff2bb6d5b7302d072c3607482d39e65d3a2fef0aaa283b13253d8790af16d8be8b74c194a7e8f4cc7c1bf307613466e4dcf14fc942b3b4fba47e85bd95ace993cd1e5fb2e1faf99ac9375ae0bae893c848cb2c0b9f07f775a48e3efd2f3b5a121fd2c96ba1362596144612678b5bdc43433fed09a6f6454b6916e30ea5e8e3e0c9dd7c61478edc98aec92d40d7992445f014bb356bf748503e1415c5f07bce0b1d8f1f4e465a345c746073a3b5ac6ee14e42769dac5d9d0ba3f30260c0798f61c916357c3ea4eb1378bd7d0169a4586ced546d2c2f0a976069e237fdc1349757b1f3be40c19800219ffaea1d06fcc14bcad1145fa2a590972bbef3d0bade5b31f2bef3c13dd8c4eb170f9f9df10b868ad06691bbb32643e4d2897fa2d50e430c1c89ab5552be7d1a5aa7fd1221538e89e827d0fd23e96751c17fde3f66bb614a20aed94a04adec6f17b5d58dbc5d4caf20da391ee67c7825c128f67089af91bb1207dffe62d4869ca56322f21ea17f5745b5b7b5ec0d42c3ca7954bd12061f2622d960dba8d8e6bff501bb7f90c3d6d48a7102b220e0afcb4cfd6b182d70ee0612a2937f1fceb5f8a88ff981f86b818bd1c7db54d041fe166;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h49a7fd31d7d87f5a11c068c9b163e439968c60fbf82be0a2263cb436ef6cbf51b7fb5254e61bc023edfe5dbc029209424c97f0ecaef55fdff1dc9c07dad4f66a7ca727972d571ad0420efdf0b51482bc6bcaba2a797c31e437dbf87cded45b40092932988b518aa5604fba0dfb2e9804866f299c11c564b305fe6e39056f0fa369aa0a443450af54c2c0bd7659f87203dc45b85c585c8c6baa00297f811d090095f326e8cb9b3cf1a05ac5390a8dd69aab6aeb10d0575550d9ce6f49ac1121a2352ec04b0837a5fb4660fc37253fa198458afeb24f9a62cc9db0c97cfb490153c3e0b152e96d07c7f49f228b5cd89bb8b46261c0fe80f6b2363ef77d7db8ec96aeb7d64c11f9c6c1ef028fc703e4ec850931a6f8d16593a62fce6c7974bdb6303bb98685e239a3159b683d1f8d21386c265e2de52bc733a85310bfb1fe2271c48b3fce950757a741fe171a422eb8ed5f859ac8c9e216cea611518c65523b91417150841c3d153c52a0cda872693e402235c12b3d816db20348faf8e2f9945286d73526cbc6c15849887b6e2b49ee2727881e9c440b5bd68f624486225b4bfd806df88c51c0d0867fe5b2343306d29f55e016a1fa05936448ed766f9e29bc4c4a7a03065ade156cfec7110319eb615066ae2f9d99ab64221d766dd5deb8a8775cb25e40fa5ce1cc316a041f3851024b9d85f18a7273e110c735a10f3759e410eb55ce73f1070525ca298ddc2b4cd1aecd3a7c1256b48ed311f5333934da93504c54e5bf1647b082bd67abe3b53cf2782cef958959d6e2dd4e521e5fc2ee8de1a370878f03d034a2417f80ce921381f7ca7a82bd360d5f38f7bc09c93f82c355de0e5dc443649661673c1961a1dd239fba1bbf36046250c7a9ac466345b136b04114b52fd41e9786021d3526bea32975d2465c83796b9b0c9c3a05923ec05c4fe104f02baae71990784b4a848305f3929818fe41117bfedb227f20efad8f226b6021a35a716bb83aa4633fe7ce1f542873f224b013ce64875e9f65ec654a0345f50774d96127a7c456531367904c110495805dd23d81906f10c90fc9fb11c218627d76de6acfbdedf4f302880e23b92a5eab806e68a04a20b79c09c82c2bc7ad35a97dedb3873aefad95b12fff24596d88737fa8d7ecdf2ab55d763667dc5ceaa2a6f90a5bb176287564cddabdcebf68d28f050fddf4b1548292dbbcb227407193d82514a088d75ca0585e821e0ebeec360f9c43220c5fd789089c7937f10cec591c455be8edd27f142421be447e652700faa5b6363fa508b1494cd83ec84c78cfd95066790964f2035a5b14180b1a670cf337a77bfe18ef83954ac96263301409bc31cce8c00e00fd4c9724e42d7d2a5f19b12087738b9031fc16d544fc3f80dc165c708bf66b952de4fac57a390ab2cbf4abf324143b47fb0723cd931747b0ffe2196e845862d01fb801bc7f0821375f4504e584cf1de2e3b2979b5460d2475d7225b239f004d4a48fcd2e23d526b15b87cb7501811a16457e1961bd239b17f2fecaf65107b6ed0e9599e3633750efdeacd4e55d81a655bb530d0cbe6e063774f3a7da8c23a732330ee6a624569d4a7f7f65dbeb16a9b74da629daa3ce2e0f0db9bc0c1c5256003723e3b78e759b9eb6ec949992cf54afaa470cd51488acbd26e0cb7bfbfb060548bd1533e89d6363abdedae994265b8e0908df33b79d35bd383906436525a56ae7954065aac335871f5cc667b78fac0e0baabfb39c6ba008e86414e617cc018f15d0ff704ea482a4d876af5ff177a33fea355bb4b1511f40854ce1345cae7598f743cecd521633b955;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2f90627c33ac3e0dfe219a66fec8fbd4ec4e05d8ba9aac22998fe6927478eec239ea815fc8682bf9ddb514d0d95ecdee61b8ab64bedc99f00b29d2f40eb13cdfbdda19a40c1a7af2a36337cf0132f3cd1ccf7bf949c019a68aae5576bfd81bcd59c881c5f75bcc5f7e2d09b8d106faefeb35823b803ef19102365d4f5ada9875d45eef167d517e81a981890983b5f285fe586063c4847713ab71bdfd94060d00237f250f2e4e23545a028b9c0014883f622baf377d4e18c24de1a1153eab11cd81f6da1bf1f2b8bcddd314b69163c9fb1ceed12093ac015d22dbac3f4c781aa0a92d61b7231cf2c5db600763c8360eb061dcd5dc04a8930222f63343a7562a026b2fbca0c8ea6cd0c1f37a1d6d458049898d439824bb918dd06bb1eb40ba4b2a014735b1612aa6834749d71128e488ba830a030f26e527747e30747ac6cec02df541d3297e9fbf1ee23b7c22a097f4571ab5ba4e852c3ed16c9e1bf73f3188e48f255aa759763dd7a92eaf4e24219a5bf8aa0a5647562cf4eb8310c231387e11c04a522d9c4297d3d7ef1d469d0d475b16f8c6389463dd1aa20c4c66f08012fc331956fb0d48f04e44ba291cd38246d49c4d52f9cf9fb401927fead4d9de5f83077962be24851ab2ae2ee4ad3e1f1473d685f5c64ab7787423467bb53917e6dc0a1232512a6266d98cd5553876295aba95d6cc454a0fc7ff9881b1edf8cb291bd5e4481b7b64ae32277e605d1dbd62cc5b5f7ce63b666a57711ab90b3d804d5d8dc6c433ed48f64d465a3ff2469f93343eec78155b5d4287556e5e134f1c33b4f9c9fe6eb8bc6c98ebdf9c5b6dd88ef2fcc1246dcfdfc7636e8afebe4f4486102a9f2cdd4c59e66fbc2cfc5b7b8523debae92befc11b857e4ea054891c983bb70094b9ab0ac9d954d70c369ecab08f3aaeadd78cb0631d0324beeba0ae49fc6babbea759e809461f266c671b324fed8414f993c0455cd78bc400291a34939579d3b38362c7bbb5047268bdb94b368fa226e0fef022b68b984b4fe3fb62ab2f39949e23046ffbc23ad55184ceada08b310c5ec325ddd416ba9d689a40cc5beee38d8d2f9ce038dc8ff6bde10378371152c9fbaffec81ec894fdcd8265cac57d2ad4e47ce8dd99e4e311ce059572ffc59ebaa4a899522820f128922b977ce2f8391a6fc14111ca7372153a528613d0c4ee35bbb8f8470bebec434fb0661e68f2b022e320070607445d8ae76927ff2b0bbcc933a4615be86bc2cce88aeb0a8ae510978e878bd90ed392bf9236f69aae1d6cdb766fcb52b6d6d272b78b8d4591d76f3a377c73c900486a7054eac72e2e985366397a4de83f0071aebabee7141916554d04ac063fca318c218ecc5ade299f2066c55ab9c4e89b80722b7e8a25a1f091963861f064407136a61549c2cebd82889653cb7895f4551a9a5b127939405ee3909c34b6b685bb05da88947e2de47995d82c6ff3f5152a5d69c948e963b04ce02018a0e7426a8bbc1284770eeebf09f436e3b2e065fc1c5037b4aa19bc14e6ce59ff0e6b32eb1a85a3c64e518982ee8f5f9ef43c32d2afc520a0b6fad1b04f39d2b2375a3636d33682d210606f72bfe9336f3e7fd414eca140cd5c2b50ecbcb7be84bfc37c84226539bc73bca7664338539494e0e27a99a548c68cd989723f884e8f5ccfaeb4ce719c76d7dbb84502e2a84c2e20e7b7554ae90931517d37991703090e97ec04c875f854951405c146b36009a55e9a3675bd1ddada5210412af8b814072bfadadf7aa00407971421a8e150bcec2f311b21001cc364f34a246f7e31f1a729497aa24c89097d7fb87866b0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hdffb68ef5f098e99857dcf613d626bee98d4ae8c9832be4fadaa63b0bbac34662be3af19164c14fd77c0c0587f83879314d4564ad7f4e0c33dad9e995d33efd37f1eb0343cc85e711069cb4f59f2f446ee91687df8714957720a43ee5188f4d139a80f7f7216843c634142605d6e76c2761890df91b3f7dfca73e73cd77ade4d6a7b62883f577bfef318832c316c21b333dce29bf9df10344b7e09dccaa7d94fc898657c394250dc8cb3eaafda10e8c7c38a188df93ded3ab4c405682d6b7b75d0d5f0e12af07bd75ce1699b44618f23435c21bbb2878013aa79eb037e09040dcbea10a3a6b1b8fe993afa4a70686f72015cb5acd255b7b89af9dedf17ec0b11990e4999caa738edb1d1ae480d76dfe38c0f84a2112cb2c5cd45cf52e7cfd9588c328e2ff1b409af140fb5bbf3e176cf6aa680d9a02f5caab2d1d7a15e6104d680afb97deac5a02f74e052154cb80750eec7c2340ebaf084ba468d6ea80d4479daa802feffd5e377ffd03ac905ec3cce8e59e5d0094780d793e5e0f334d5d871709cf9a59d17aa174dee9f0242c9e7e2095101a90cf0e31a4bc44c6d671123c6756ad982f4f436c1f79f52cd89a44eb51095bc9de67a52c69eeaab4f7701239af9766cf9f2939ba019a3b29951fdb92b8df106d76cd8281d4b8711bc583b214d2073dcdcd5c53da88f58df3fad2910646d7a4b24ecbea82b3c8f1f2dec8cdef84b0008783feb030239fefb68fab47f3a06c744c9e1acd8aceaa2bddfcaa1c6a44aad541b6b13a88c125ef93e9a79bf66985cb5599c9cb9d799207a0e29bfcf36c2f4f9d72a7ff14aa58b9e525384df637cc0603ea26371c174ae9e1ee3bdd8f8d3572345f0ac8abe8438962943be8f9c8f1ad93a9b8ec8ce132b24ab0aa27e5d771bb85528375e032b589ed42e21d3d3f8565865d63699975ad55a086435befa00a4e3641d0164371a27db99a69d2d31b86c44306b3e51c43932931a1b1378bfd91de6985a80e4705e7fa357fa73ae53fff46fe3c355044a1dd80c5f5f88eb52bc15ecb849260be5157ccfa74d8f4e6d2319c21a471d5d6fa4cf1360f92371d417b13dcc12f11c986c6a6ecad290b31d749209c4387f82fea4f362a1d390d0e9d54d1f99229f42d074a910a497c7f35cfea851fd5317bae7e3e2affa0132c2f01836b572cd52acf82f93bc102b09c48d5cdc8d5645a5dd8c8544c0ac977e8a194cc24445a570c201ef014b83acabcd46e88a18132ade14c71e8e0f62d191e29b8f666cfcbdd8ad8c07044618c2ae061b4f9d201ab4c7ecb4b2243bb48ab7e98d98663ddf0c26272032448d22e95baa3942213c40369168e996f53945a227cbc5ef4d4271d0fe84a391459ebf379e3b662850930f5b697df441a85eb55ea924a6ff209df08713464a44c2ebb200a2746dc690feedfc0370d4e8febb12b0ce99d2c8a44d252bd00bb90561a6f2c7be41168c3d7b2a1e9aac88ab38892ed749ac113cc605117d09a50da0f369cfb8233a97fa4a2f571d0064676bd0c008bf52519de705487b80bce812ac2730dc668f526b426fdec5a4e44c32f083c34237a27521719b384b030bcad7ed4a90000a8bf974c9a1ff40954d4fddb70bb781e1b7534fdb8fc67e228a55bc570424d184662e2337ce75356191c2a288c582bcd626672c91bc5c3b7bfac41870dd5c1af19315299748427747398b2445e0ee45e7bb2a83a5c5ab8b3494a77f22f6fa976d6e38b88e2cbb16e6994c3d477035a479e216105ef4d06ba5c078fb76f34475548a887bf1515e0caa1075682f7ae71ffb59e07701a91aae2cfa6ccee8b48f5f01016af9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6722268ec2e49d3a07033ab23c6b732b596ff7bf3d2ae8ac84e56975a29051a5a6715de26e23f6030e73a02353fdcd72cac53fb1c05348877267c34155f833cd5d9713beb4c80d6d7ec03dddf5ff4fc240cefb6d41da66c72d63c0f74caaf6eaf860f9f846edff6bf73ddeaaca7bb80d6c0ea9ce60834003a5ecd62a444fa6da371ce2bd8fae3135f2b39c1ad510748036c10165d837a17a4da96923d88e7341ae7edc250423e17a61286de237bc04f7e29a0a92caa2069f23c56e7e991cfca9896649687c72e68d583b5d8db9e7aaa76fe49e22dc2a4296dece52c495e214c87fbecd599f012fc53fd75574c1656af70fbe02dcbb3dc8e5af471c2f7e3937fbd5b69aad0b3b3544c064b259ad1fa363c4e367f8c378b964b472e44604647237d4a04a0e6cf3185114d3a0f33cff2f432173063e5fd448b6d667e11e0a0d11ea64dbd5fc66bade736911cdaa881602102ca9e054509e668270a9ebcbd427e202d3d77c832a185dc68ad0e1c9eb4923e5b8570d5b1d6a98eb7cc05d4e932334770a4eaf78f543e325d9e16f057d1900776027b825666e6bb43417d65414f227bbbe60a8fecc66c2d0f0e73f53fc99405301e1411b2776506d4bcbe1766b69d7f44d7955a494a02365b0f9721ee395a936d289bea50a7f2e2d519c793c843060703ddc1e129f15b2657da7e1208fda40b820b124c0e0ffa0645c7bc1a44cff0b29caa98fb709e947b0137ab3ea2ddcae3f47870810767d192cc1d6e091c5b177815986f42c817b30477a4b268ba15574b8b072002aa4aad6b2e11b389af3921e07de6016cce29befe2f6bdefbf68254db785ff488f75ffb00390b0450f5c7f244ff7ca88dbc40c5aa6455870dd06680ff7ca15b655dd71d10adb778eb35cf8a46412b2e805cca70286d88b1565dd3533dabeedec67ffc5f3c4604fb3c8037e82384ec7f55a607a902c88037f50056053fbadfcb0eb2f9bcfc595cd8851c987e6245c77e0a6515925b73a5bf61a035f2104e3ca23e67c3e90145764c8ed5a697a157c0aa646cb8646f69fcff27138d56afe6a443d7534c41c7eab5d0f272e375b672dfe4cd37602784ad40559749871289934b676c7ac01b898e7dd11e61f082e4a8c2b3d8ed11f9a7cc95af4b6358070351e4a78e7ce68714a22218bfd9b82d98a53bc0e61f35b4efe599616b3133de3d338a9a5715a3526ef49b714616b20be22dbb0c2894937084a2d6e51f1db82c2eb224b362f7d59773a70cee2220443f4b91ee5aa50a3ebce75ad72382d43e3a4da63ad307b534fdf99c71aeb79e9d2c886ba96605167de9b86c407262e66f5f9d34ac7c2e2dddb2c508dba154028d41d2231b004f8e5c0a2f4451d25a7ba0eda35967ba5280f57a79ce2d7dc289874944cb6306e42ac7de7197e9dd8f5b0b738091f992443f05a3a47fc9fab35edf431dd6d42b9ec67b0f966492bed9ff4ffaea41595075644d968cf98fe3802bd31a7e769425eba399684d538a91f37d96e33b79936a70fbdf176124462c67090b64e78152676dd3c57c14e0760269a1616a5d1c5736b327aab29b0bfb91bb3fffe2f71c0331181b652e926c2d033e8d1b343c34ab0987969bc71e77f87fcc49cddb4d1f4ebfc65ac5ca754a2ec6ef80514dc2da0c1a7b207f40fce3207fb88f07eb1d0de6ccf698218b63de5726785ab8c14769f10d18c09a736794b98e5f091436a47acdec3e5dcb6d53ea735ae5be1460e42bc04981bdce9f99abc7f2a66d79542b2772fd525d11277588a5a26e98cccc3931ed941cf72c3357182287ad0eb1058e16e309d6a1723d120aca4a006a4162b60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hae48606d37baa29540022098e45ae02a894e35c1bb2bf0ebaa24a806a9bca2c5dfea4943c70d49f6f5472a6cea261990130db3de85583212a3ae6ed3fc3e256597801a967c9582ccf744cbcae5303003fb21bc1337440dcac6c3ca74598ae73d9551365d8cf8d5bd5298c317cd175997f66e370a9f059b7e581bbaf6e4b97f4f05573e056888f07be57ee33e079a94922d0324fa8776a6135be0b086d3c980ee9779c257ec930ea0d12dfd62f472443c97f19ee51ef6c77fe6dc2044f1973425c4e606d8b8aa3973b691e839c09289285df1c655ef8c03d22583a2c1d8dbfecce97c83593aceeeb7931bd782b52ad79e881337d1f4230ce92c35d58df98ce81b3fa5c9cfb31305be8353c6b628ebaa0ffa5528f21685a38383cc258ff87bc1e1d5b71061ec292917cdc50a726077cfcfdd22c9c6e8a462a0b0ff6b56b386705086ada88a3338227268722e32204b55e0f5120bfa9978c749aa1de58fdaef042ce57fd864d64b2097a3b4d0c94d49f1d500b4f0b1e8ec3de8435615891d88ce0054c6797eaa95403694422c4b2213dfad8557bb15e86c4ac68c09abd171f21cec98f8e680d27de5ae4ba74d1ea9b26a95f88a57d2898b89c498a579b343499ab4818b622b1d93e296662e299baf1bfe01918675b1a15e4d1222282689e6462e7b6471d514fd163b66a9faca4d55f70b63d1b6b9eb2f3b5402196349d623bf5db77890d603f2c4dfd027afe02ed14814c26870f95a394a93f1f9a3354015d499a77ab9f7e0aef29e7e43052a4532c8db33cd6ae00246c9fa2723aa1410e0f5c396f5ae6cc230d3719e89e01da3ff98d8ba8749218a1741b06264de2ca2e880fbefbbbf87fd25bdc9674299acc5041a20939ff38e40dbf227eb3fcb0c88a234505562268c9f36c6627d3d5128f34556f86bb11404158f6bc10b77b9f85bc6563606f3a0eb208b0b2b24210364f8e7443301c9dc8798338568c51a2b88a8efa4be37f3229782fd7ee2c13fe3ee606da875f2d9c2c2b338481a181facb1140f52cbfea097b91ee59c479b714558d75f0d5ed531b7603bfcbd586d2067abc7b73e4ecd90fa66d88c0869ec1262283cdd6ac9d7209d9ac41e02fa8b54ee64e70a35a3731f5a47f32aa4db2f73765a3c81a0ab6d66bf4f34802c88a6609a2c7c8398de2fd9d43b6abbe45679bb9105a97e0572069803c9780bf037a1806c166887ce902f65cb546f9a3f7f3a5e74288e69b24cd54fcab7c2661985bd2a6892ad8ddb2f54d3ae27cd43ec738c8cdf8a60fc8b873da20ee5f355dcc988a6fef4e27ac84bffbe37e971abc3532cb42e1c7e7ff52936c00a5d37cd76690c94f80d32fd31d1dbaf2ded969a6db271d8fad32f49010c0fdc6a29b711fd30357d285c50f96b32a1fbfa65dba93db90c4680bad1c1ee4918d035eb43b854744ee337e2986a98cb452e46f1949651d529e11b908ec8aaae2eed00e57aeac32a60e8d0b3da250b5cf7b5bb79cde703454f3de7d6da4817487c6ad177e20ed8706d778acd929372d9c77b4a6d3ae063aa78918039d4fefd726c236bbfd785b416175bd88c255d0746f89ff3d8316618b15321365f6544e2caf27870168c69d9be075fc779d0de752490beed260c2222e77cf5b704512e75feee0aa9cdc000e179128883cf819f58000e96ed16bf8d107e7697a010d08c29cb83ca41e3ff5c410086f9a5078618031f99a939e9bd207a5fb70088e6eb14a43775265c5df18bbccc42775ad8ccd0bd5404be851f4ba7d3ee802ab7593ede0cc4fa8d88af14920da39fa22c64779495995aebf9fedc473536dcc30414912271fc23;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb35abe8b421075f6a8ad7999c29a53153cce3d37087255fb6bdf80609da8cbb5d0eacd2fb20a118690b231cdf9891d8d17c7bc99f149f92f48d9afc768e7b79ead70f3a283678f734fdb252ae4ccc2b48c10bdebf8e0e86ea0d03ff7c3f4d2a8d6bfd62c0d3e164b2c7cca2a53456200fc3db400213ea8648276afacdc934373b8ba4b110a04f171806050f6205b3261b8a5531b0de4b41d17b8b899159d2bee81e35a596893f59bf32536ee4d47e1125721a80c584445692b5cbebba38e14fd292d82f8f73b28d1e865b0d9d22b4ac7e8f8c174eb69d157cf2201e9c4df5f98ec666db66fa1d0c12e20dbebd42ed0ac83a7bc77253ad6ae71025021fc050451e7dfc7b95a1f8366b05956c2cd0cb17166aca59af873a0496a5a902523c4c24a1d8642099b273cea53b44bc28f873a3e4ed69bda0528749b801a5cd2800036d872075061986a1fead11693d4be9ff509c53acad245f1c00c2aa227feb08a450a1f555e39875c089118e598afcbac18774660501b13e6ed134e41c5f694e04ccf265b81970b933d72af6addb69c5b3d8b59c5aeecfbe562a09012b16b568abfb44b708d3257375a266e6211a5221ab8360f77a0d040f6763be880e6e70c64b50f61c584b9e74d114859cf2d371f54833f853a3cb1420ef5a3fb8ec35ae7f4d2db1beeec67775b39347fe66b253a75a59c68fa7f1088dad66e8469032a31001a2b8a1020e226ef7c910ef6ef0e90665663195497b9c75f22900c9ce0bb904b2754f0c83e9bcff3ee41eb1cd8590d6b9867536001e4e666c2e28d486393ad0c93d161ef22d90fa336a6816dbea2773bd395d688d64fcc4f7145547612c6ae11cd7b99ad62e0a000e5cab318adec8f2af0e91c8bc71502c09df1c41bd563594fc85d2d2040b02adc4f7ff5a631eec5f59f12881903a764325e8b1fa3317cae0199ebad7541dc858f8a0ec970c8fbe5b81623daec53b7cc28176d3031f2b4ddbebee980277a39a55b55eb044e133f4e2c08395d8d37dd75d47ef26fe1e63f1826cbc69d0a113484fff97e2af18b5b272085642f0399b052372b4e648e515744626e395410ebee9c8662af8b5c4da88579abdc556b8873a260af652d5ffb477e07dbfde80b7f5c4165b70b27945451608ce244d97c2b7ced9c3c34d5748e517f0de87a99c179b0ef78febf76ff049f3eead59cdf90a4c3385b216240c042159f047d2220d786f7bf5b1a44a6d6bcb08c314314f166f7f65374fd437c18f226adcbbff29b4a761c89f79debba164caf1dde01eda0580ce45000d590d0cc118b1fc1d55dfd2ec7005d4ad56104f0f3bdc8239d2770f990fa9e22aaf470fdd3f2430abf0ab4824d633fd1a8bbcf077a4250ad1fec535b51c581304626d85d988b335b0b5eac0b72e585ab6cc18ccd819bae9196c90a4126f370474a2f1e6b3136de85bc90898377fbe806b3e4a6b02a218cc8c8ffac5c1ae4e7b9abc27d68d946a0ecb4d5e6e508fd3753a6cb884a0112d00449571319203c1df25e5961ea47598455a8c36478f7a4e3140f8aa626726340845f36895e3109c5131c66be5ab76fe44f710066737ca9b04de135bae72d045a0a846f98051ffcc87fd723b5662c7a42dfa285bc3e606c19537a4039bbafeb735aef2d5f5686dcf56dea604a959cc19d6ca8198667032b5ee72b1ccc8161f9432aa31454a55763f32e96c3bbdbe8a9515a54a239d0c59bc326977102a2ba6e19be970e7597ba9359971fa4f52d786397779482e316a8c2395434664c607bf5569fe5f0dfbf71157f209a9a8cd6050b78fa8423158ae32ec9c8daa7c27dce40e0754d46;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h29613b518ba21f4d8d7613407e8f2615c5d4b46b6c20bd37a9fb843f63d149451c83f3da968bb324705003edafb7d6545f70478267f55fa13de6b1dae85da42a1ccd40978e9080592b7d154f4eee1a08bb398315bdaf92516fc86027f84c97f3a6d9eb56b33bd32c8cef5952c81810b307acca6d85bff920f061fd2a66eb9cf3752d0874129f2efa9ce444554677bbce960260e28ada40d106ad7bb441899cdcb5699bd67acdf13ebe822405c570def5c57221e70f3e5d09417cd0fab6a5ac1b7aefeb8106325cbb67f2942337f79d2cb8eee4b63d4a280c9cd7ae6c830cfe4b38c9c3b166d238550a909ca5d1ac11b3fefc74b69ae098af58dd60d180b042eba2cbfe9a61dd260a9f030c08b12b7a1fbf427aa3d57b98301b6bd59f52ce781a4131c9b84c3c8dc8396402e1c7b1faa06dd0f83249c399a6a4d2db6fdd0e8fe760e8aa97f45a69cb862e3b29c44094dccbb721ecf4b8311e6110cf73a5e80b4743319c4b9412d75c84321cb31602eedc8da2fa8dde733b16ab6b1c7c6f9fdcacbd3ee3b3c3f419d66641a808c5b5a5af701b0c839b275b8531f45ca5f30698986f356bb9e3953fc3e5dae333448644806efea6ef64dcbd200da997aa57d697533d15d4dba1cb880de9bd36fd4c904f26ce9db724992a2b01664b3ada72e016e54469aa848bd3aa71a4f784a01159dcf4f8b230a907e74b8a0961812a56871d7948049a29236a69ea631ecda911976d393bdad9696939d3ba4fd3383b9f604b7a06257c792a77b34c2330e1d19e29f915301efd0403828ba28c5c84e68de4c8a2885771b764ef20b4d404ca9c17b8cf804b8ee7725267f1951682582d8899103ab7c72e0c914509e23ba7efdd6220648633ad132704df577959a3823c193cea09434ea3fe6806289ade9e89694123eba87ad0dd69462c7d7668049e15e127ae2adcbf50c7d7ca8733cfdc8cb9bc45e163813614ac72bf1e0a16ee374dfba73b83588fdefed2ec1fb369713d1520c3f935f02b2885409456129587b35e791a23f093de6b38992c44823d93084f7594fcd78465bd658f5dba39f17387f64840592c2fe5f8c47b120f3f85beec4f8016fbeb37f42befa19e8c6e76299118124f6b4915155c8c4df578221172f78ae994313a24223073a8d72c754f769879650031aae7a8c2bdabc4db8d7e88ce2e275b375b4bc1492993cf41d8e19a4c9691b8596b2100adad8ce530d40d9b5334f74cf12768dc38f2ba1bf21b4e3e86691a3e40cac4b9d1c80b41bf4303c7623f421d9ca2e77dfd5cff74be65b2259572d5d466841a28bdcf0f4891a44441aa348a01ba998f7b50e101d164bfc549cd02d1f68eb798bbcd1d710b1e6b50366ea0ecc651a3c8a5897674d148105f12085e9b0040cd69fa1a43b2bc355c49bfdaa554b83d61634d295c404c932f09c0ad9afa14f2c68cd4039648c093a88dd0497230d911cd8f925a06d18f49d647cf2c04eb0afa0d37e80756ca8186af587abc1e304811a60b12a8c3d267bb48c27c292a427f838e609c925b5d57a2543c5545c7f2ff9bf9d582bb62f10c2973b5bb0b9f4d9419db1e27612f8edc9f148cc21e71846e155d1188c6b2115ad9c11636c8cfcadeedeb5efe9323ecd54fea98e61966f265f474330f48d6a4be06bc199d03ab622a2310028999a12e2939185eb2d86818d261606e25b604a62356f5cc33ed5db96927a762f2b396d6fbd0be9c5e5e024cbd74de2a6fe9a6a10e1f1adce0836c0a9a147db40d94f6673834fe66d48eee6d437a2b6125fbfc5c5699a04b4f30d8df0168e0f03dde3f774133574c10c120045a655b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hec68bbe71e343360d0fc5c76fc616e8a36f5ac39d845664001626d692ee5a61cfd1d00bcf9ce22266c469dc0601c37323666e9a2bd5f5db13d13b03e173539468dd7073fb238e127aaed778dfc26348e267071421aedade99612015913797be0b7387988a8b0a77c047fe200fba67a86c7db2778269d5c62d4dfdab41a594daf8124f94d81f71be157c8f4bd097fb35645cdd56e85d439266be7f20b31e9c8c2b05dd480a02fb79adb1356eddbfc87c2ab28843aa1769f70aa3c34e1064ea9749b178655f156ae28086a4e2147d7138df0fa9b7a64fdf10cff9fca6681cf62239ee906e2c69600e453f6ef6b6d1d298b5a19cea950d76e7e363b8047d2cc42604cbac9c530d48768ab5737bfe6dae1df27f8b915980d96d91aac3288db74a4d4e3b17dd2452ecbcc37f29d108a6044788afd979f3e15af504f35e57dfbd0bd06ffd7a5d5d34bae549b86bf2ca118d4775787e9e9a068b385bb150082f310723693277fa5aba6dfc171835df7ec26071f758f7b8aa57866c66a2a1a2d0f05865e1e9728cc12f4b8f8add573e1fff978ef8437b4c1a2165764c16fb9236e2715084953d2bde47b63c57b200017612a10bc274ca39bf8b8d41fc7fca5766bef44698fbdfcbd2054004a028deeda428eb3e15a984c15f854082487d0bc61d0783c6ceb6e9832e982b47a19d6adae493bdca5b0d9ac1466838c6a0b264141205209553a0280977d847c1669108ab961ebd119e21271945b4641952504ed3235d8dfd7559088b1800d065754a128663ba2ca48044a9a3ad91c154cc0805a6e0bdbda469dc3dd45dc63517f676ed0f228d5d205d8a711071ca19897a37982da5a799f9e21993a5a25ab9fb317862ede699323364da0aa350a095dc38a8c995e3a5b817782a3ae2d946c865b2ab0d9eee606dba1ca65bacf3677da4e37df2d13f15103edf5293a3bb0cda5f34de9b2474ca6ed765d7cd0c00a011af0caa30203079ea28731bf9fd623463211f6b561bf7afce8e73a64025e78acb3f2405dd70e56870103a5d515ebe9d30672aa6d489baea4800dab7c458406ad383d02bce2f4e25fec8d79834ac586648dd195d9dd368d74bf76013d1d217c56ff4460dc6e54e2dfe334ed2e952925107e41733949f98f8f50946bc873a9eeb7bb53bd9ef36e2af0c63d30ad3da197750858224a31626b83bc24d9ff33c4c93e22374b1ef9128407f972472528e9a0a7ce07f14d05546591d614f0ca07a14d2f54df03c33efde57700b30bc34a7535032cd92fba7cf8aab2bcb34a5f9599a47a03989df7b411494a68be2ad6835a4af9629a51b7de012322bbb038acfdc697dc3ff8ac90beb4f6ac43f367fe74b46d8df0eab5309e16c6c92a95655d1883336aed765282553d590fdf58fae0a733f538e48be1b2d1d1050135146d1c957121f34de77db6276c96875d16e9387f9b9b6eb441a320aeba877b5fa036dffea0e7d46e5cb43250868fdc6d21f52577aae24a18574ba852e6a3d44f9c214d157a41abef50ed940eeefbd6fa198526380a60013a6da29203bd558d1e11b5c931672abd02fe4358a3af17e4e93f95e6c0907d9e90875ca2f13fb811a2c08984edb117eda4cf701aa4dc0288083cc58e4adf8d5edb2c8a5f731485fe2c6fda7f9eb9c4246e2ed13eac3f45f1cec1e3c424f8bbefd33943ff2d141b18e30d383e42f7d36d6af1722f67bb6c22942efca2bfd432a3747eabde8420b47003ba42dd6e28601a3f5cb94525be927d554391873a467cdb0a62e3149df8aa306610c8add973d51068329e32f53da700dd99d4e427824fc05ece7465eade0186002b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h64be95803ce6a8c74e2eccff136b9a30109f17cfb91d5707933ca7c2eddc03bc919e48f3723d3aac6569bbfa4a8550a2b3032a501ebc7a5a0935af1fd2639b8c9cc2a076e495f6bd5f3307b02cd1045b58f439f1fe4f30f52aa9b5444e2f8d838ad5d7bcf36b9d49b48cce31833d8e045695fff74b0cb8aced20108687f2ddce7db93b5a323e6c16044e4670fc414cbe39043247ced637011211b6c078e54902000e73fd1c528da50c172b123029c5c7bd6993fbe75a0127dd78b76a88e421eb898872a8a9c19bb8734ac7d65d0fe71321a32e8e53ab5a19b483dfa4a1284676457a3d670fca3c6ee9d217b7bb2aa1bae856e79c2aa773de2e0d2802360e52b0e298650299666858487830ead51c64fc32512e80b11450557f6cba56e46feb652f9aef77691a49ea61cd56b4f4dd60524bd543983d2a86f48e61694088fc5f6c78e7ef40642c13cfa4637b311fa87abad8373badb216831bab0ca27d6f1e88c4e1dd169556c2d4a2e68b6957baa1de5060dc7a97ecd6669c11985004b5454ae04f6b1135fd59b82218b5b8c4d5a3907f543ef6acdb72985bd389f489f043992bf0c33423b968ce12cd0179e9fc2ca6017349706471f116987157db8845835f0f3ede6f9ceb47d54844360919fc74e07e71582c4cfe47b2406551946d8b306965834677804835dfe08480334a39a8d84420404213619ae0c580c619170e31df4b1440d07c5a8741f4848c4b02a170b6fac1431b0c8ca61b0b023ea602400502fa44fc8e0611baefff1c67975d1bea1124dc0bbad43b5c1d23e0a56d11917051f0cc7b5b15bc7c931502ef450c87aade91c808bb3bbe23be7e5183a2bc3790369c0a35bbbc03840ac1ee1caab31b21aed4d64067d7666b1861dfdadb3ec470b011ada03f5b11c6b685e6ff28cc51e05ddddee2a27acd6dfafc50249b24877d5c0dc810c64fc0c978cad2155096f0ed27ed2c6e46f037ea84dd67cd052df446a34cf420ad772cb5321030960a0b9e92b4d57b425d04057e40f406531752408d755a8f3c6266176494017355f55334b8c8d0dd6c6b41d2b2665db094cf3c199aa8197094e2f57822dc9d996b2f8ba6948b5d782fdaf62d74426b16636bedb32d511a69991b0ce4a51353de482d4e7b346071ad54600ee48ad230598c25e9114c65e50c644c021d466a554ecfbfba52486aea082bcd578108bd1cf389af41a149cd5d55b2e8c7fe8457cf6b59d0a1905d3ed35fb3e80a85c914409d11b311dcaa6020afc6cf740a10e10c38549626e2ab723052329157599fd36f3987371eeb810dd9967887840e6f28a17562ac78c4be1f10d9e9fbc39b703ef31f4c02fd00c2da9761a7a872812d2bcaa81c8ff0fbea532b37a2c13eb4cc49aa879988fb55715f88027494def82851308990d7733921842b3f60beeebc919691ec956d2a90784c97112293696e98c1336de2350cfc4bb0b08fe671493d0579f30f5363cedc07348d5cd0403c14c3d0a1a09f97fa437e00460a63dfb8d7912ae40b6e01c4cf2c83d42e450de19ce9ef171fa9535c402e0795ed1ae224d5e117c5d2631db8dbfc976828c914fc4ea2fd36c0bd5a501a4ef74dad196d8a651f86601f76babb648e64c43c5bcb9ea5573e7483df05f527345c9a817ff6917eebd691c6b19a51f024a89ba369cd11a3ceb2eabbad2d4120e6f24b2222e77f715c2b80dbc108c13b031cf66414839426814a19871838936d10795b2f6664b8e4e72454b09ef77673618c81b064ecc7cd71084749fd11f1cb45b3b16dc5589062a268fe92e3e21dbfb23a7b97e59db469170504442020c0d13db997;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7d8b7636a07c4152525a3d1aedaed2b9501126b709e631842a017e5bc17380eafa901224bf5b084451d9df720d9a14809991703ca4ce09c9d72a32ac5e4842ddc48f1b88d6003e92533de08a6dad19020650a27895dec45a11adc6521818693fc08a0a5f4bb444db3128413f5a787a2448cda3f55e6126926a1282a74b8f71bcfa98073bddae4c0f00228da912b1fd24511d2fd5dba415177b5145517172050a357526113df05f5e3be6fb918ca1099fef62a48af738917fc6b753050144460bbca1e289751cbe8a9988259bb80de4a7d52839c3a06e065d3b4289f4f46fec3d3e5ddb7392fd0b0829341523d4fc39e42f9400e2728859a10c95e45f72573c44a4a9ec808ff8e62a4c6b1d34c96885251e4bcbb0d4df1c34694b59d2670c1ef5c7899d18dfdb32956646b641cc28f06c06450b6a59dc080170858bdecf8c8ead6cf98a222f035628cf98c7d9cddc272ae329e2380d4cbcb2fc338c5693053cb3b3acefcf0a8fc24c83affb98a30d7158a7993eedf8f858ddbe4733a82eff15dfdbebde07ac04f76734e21d4f3a9c7c1a4046afd0cb46fdea4bdf4f7fe4d249dd298df95b2d4ccadf0044e0446a5ead67fb69d5f996716c03ebc3d96fd182725e990fe1e95407c6b24098e695c7fa78c0702c91c2bd83b775b1c42657f0d0c7b162fc4a488e4a6aadeada8a165d22d0c038a6f904a9dae5ea2841b07f840b95f00e5440becfd3204cfe8eed3f67be5c2680ba5876f20721352755de210101b003ea8b196167ba01b7b5ab58783fc6e1ea2ae66efebf6ac7b1c2796a2a1936db0729293e505b9733c4bc9ab4d587da29dbfc1e43b064e4178bebca0311d620b52277d203bbd1595a7414e8a14dfc008ba23597aa8389dda36748c086c6adc36cff0e88b468a9cc7948cd032b6056320439da11e90f52997629ef0b4b2f231bb9682efc66cf795569a41916011cc27d11e205f4e5022d2a6182ac80a61b521c91f0cd48a67843701ebfdfe4e1a7bf23f5105edbd6e1b10c4e5c151e6239bddaa313132e3dd1d1e296de5741367b53d1b7119e1546857239e16aa9a948f2c98fd879f976ffd3bb1ad925b347ef4e14eec3fa992764b207182da0b28173ddd6562cbf36e0a261f396da275eefe238696f2220ddf56a8d9cd72a863bff65baff3d8a53704e8e97e8ce10ed15796d67143446ed23bee146034161663a0d4c6db124d4d930506f18155b2445839e4155136e15c2accd87a6c5ede3bdcb1bacd36a80abd14a943179968c7f3d91396c289022838eb8574d683840752c961811c38c702338339656f605f51cefbb035a2ef57621e0fe07c6d7a1635eeb1a6adcde2d094dc25cf9b62dccf349e0f838e3512556e1829f331e04665e99bb34c53e10d284ec148486b021f609788bbf030384c80860bc9edd3874d7f34f734f1bf86659d9e412a3dccf2979ee808509a321a2ac31886b7b8a43f97d1672f1f5e0174c52480da9fdfeb8f8641747d57befe224c197b55a3421836ee4f500b1856c47da5141918573680c9c704bf341784a995d2d94710d8e76d2b18efebf0a874a2480fb9cb80cbcc3c27afc3a4212bcab5f4b95483d9cfbd83ef2e10027c604c2dabc707fd9264c751751562a44952a9b6c96baddf4f545bc0cdbe2360ca3396aabdf86f74b82ca30eac1bd9aa19d01fbb8e718c35d8469995aa01c38c896e1a83d0d7c36df9b98119a787f69247456a61ae0599ca63fc275993590b4c20646dfcf270dd0703dfffe3caabdb369394020f57c89cc543ffa2a71a4611c871e5d10e13c1ffdd0f58aa5767ccef75d94fef02a3cfcab4770;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfe5cce82c0abfb976e8c26d3db2b0cd058f2a78088cbd8e97c037975edf813c965a2734621deaa41fbff2a362f003451ac34ae5d2d4e058a9b9bc239dba3e83a232c4ba353d783aad4a3c9d962b5a7d9dcf97e6b6e495f94ad17422e743dd7a88cbb2e17a2667acbaf80cac51d9df20208c60abfd14aff2f78194111cf625c9766921c3a1422a02de0a01bc813b5ec78c4c2f5b16849f70d5507e93ab269eff9f7ff3a82b520d6def88a97c36cf3006c94c0488a0a1ab905a9723766d9afc0938af6c08d5406fe1634596a4d91de1a3e5b428890572857e70e522b59b1ac6cb11c782c003dce459bc7e5381d2d9f722befef2069d5e2880d789f8c8969c26f2733a378931d6bb831792b9dd95120620d2b7a5c7dfa8646e1a2337e27cb80784b463e1de6201655da894667c3b04806da9f45bcd9c84a4a612ea4341b3b39b6d6ea026796fddccd23b3b9ef0720c18d46edd8ce87dc4029cd4d7fe9a8c52af52cc1e4efb8517f156feae367c0852a7f42160666e81dd85b36d600521864d2a0ef6e8a5bfc80eefb5ebd8aa48dbbe5362072d4ab46e1d2685d82cd801eebc5415c9fc280c8cb5a3762a6b9ea9129d8de732a840337177ebf7425811fdd82180c4770f94556ae7776591e3641fc989d9003fde5a1c730fbc39040454293e3c5575eadfa3d1f0795eae597c370f90370c2fd1f9b774627a8f4f7d09e04b454ae577f2ac2d1970b5723712aa050b40b91c54f79d3b3ef92e395feec1ad18ef22268955c58e22d9aa189e57b6c5baea919f9585e88533dd079039a631d5cf10ad15b54fe7569388bb96f68067dadfffce0c29534289f8a6e362a06a5bfbd080c8dbd8dbbd5befa3c5578250993154c089faf8d1815dca5f829a9008fedf8c694d1b62a0000d10db87be78b33742bb1f255987e7b5f3166cea940812f1adec78991f5d98ea6d3b91f7a84fefc57f852a941900f530737531933fd760033cbe0fe446a8676ab3a85c8d4fb8cf6cd8261a2c0e9e35c05f6e1e1d9d87b04741639287d116942d492bbd826d54d758240d6d2ab8f724b42807bc363818d24bc72ab676c27f7760df458626f39a204eb086c20a4cd9e8b74cea1d0af9c2066fadc3e85813d7e3bc4667d24bea7e9566ef734b9ec941a497440a7919da7a7b7083970d04c3036b14ca525a45df31df26c415d22ee72a4893f691b48440a9ba542770c462ace8c437757b28b89c2cb0d9e219b0bb598f109324b4014bbcec3f802d4b790426dc26c2f40c930b0e690b30acbba3027251001f2de522eb672773531349abee8303c0f8a69bbccbb432c42a01901a36b35100b34ecd7cb484f8603adb1e6a742b2814ca6541419f9964ba560b4a933096010a9bf425f23f24f53f90dbadb21452638bf50159e6578cf1f2653892ed1f35385f07a13a81a801caad61c501eba588ddf4fa52c8ba9deb572630e86ef71591f84c23cc35a2ed67b28437ec3998e1c3f4cea6b8fa0253ce01bbd959ab64f7e74392e0d598acae688ec79ea9374d93c494bf9068b5a0b117d0fb7242784431998285b2426d6d3fefd5f0ccbb8a105d8db5d86fde4844bfb162805768f9f3957b90457b0529a3f081091f4b3261f17988c7c560754f87e25fe2c00db757d57cb47e80342a03bd5b03150d92e6644506de603ebc22a7080289e9e421c77e326c0b84e2487d685049910a957d30820a923d10816b413ff36a5019ced99b2013a02d3fab5173c24a90e4eb207ead1287bb042ef249c349ccf9239af5d6d5161b7f08d3e86edf65bada19d3630b43aa1f14f28858da21fe85b49a85dc804fb5365658597;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he63e71355c01fecb91610a69d50024680469994e9f2b7fb2f1df6668fc010be638a87456e90b6de51ab0bd1e961ec3990b9a805674428abcf09eaf2d85fa1a76926ab6076ba42221142ae24718b636cec8a33fa6e952c93b73d4765177d9a2cf315e2fa086c414f8418d130da38f21aac925f91204db0a1a7342718c5cc28fff2dbf5ac47f1ba9077ec6183fa23132634893ea24141f16540bbc0e4a31491567d9e92dee374acd81695fe00056411f7556c9962c1f0a4e5a1967cea383589b5c0b79da31e4338946f457f5f1232118c0345a14a1d2e5c4e0afbf62ddd7a12bfe136aecbd4ace8c62f680a372f8485d44aeb3614f3b94f56263c1a2020718a440a6fe66fa70dd628b0ff274cf5e644555db7c60f646f00b4e873096490da9322c65d1f4092256f0074e517976b3e6f5a74c0f74bac3183ad20dbf487896e32436183a7c821dee0ba1f7f5668175506ddc3e2f195165f7aa1c6f4f0ff72e7da66ffeb60ee3dde722be0474757895adcedafdab80b777266a7e89208b2ed6dbcd7325a19fba8b938aa82a9fb5a9b1390d0ebdb1e86df009f0b9c69fb828028763c70caa77e4ebff84771990b6245e18ed7740dcd20a2b36b7ca94c79f0fd19ceb473b37eda2405e43e81e7701053b38b1035d35120b5f8439ecd4964134e242429abf8cb870021fbd3505469b585d04ac2d5b6655061939c6d019b53afdd3e3f02542c391b3e1b04cae7bdcee1478d00e8d000f222594b288d35471f6650208a58528401764c6ca93970aeb2b5863f0bd76755d11afc4eb5df311ea00df3391748af20cc8f31306feaa0d8dddd1c2923a416f24e084ee237591eac4727c494597e314affa61cf6042bcf43625a3dca4349483b0ccd46ecafbf976807496b9b66e7d372b7cbe856dc2f68fcc6a205ac668fb4060abe77521950445e8c15daa34512e43f3dfeb410c0ffb8fc0c4f5bbc6eda3f582576be95cd4efb2a44fbec42dafaa2637c8af6936e664acddcbbd22711166124778e97cc8f5bff1176e2c8fc5421686228abeeb1789589c6bcf95d9f4c961de492fb798be297ecfb2151fec151d09f435ea1290e63cd47e493bd2f5868cbcc88b8b3c236db2a721ff5272a34d370556f2b07519f3578ce32675c3a409fbea66c4303634c072d33d93df9ed4fe1aff5bddc1cc3e4a4d6c0d30f01f36b1dd2c781e20a5a6ca93ca4c93d061c6e90e949e52f2e404a22e82aa5c18320befe8bc2c967d1d1691b6c3b4e3fbf1e3c77851a8cec05ab3e9bc507023833a36212f806c34d7b967a1b10b262dd1a4fca889ddc6971134f7c978442344976da71feec8b0639ccb57348bc6812de86d56a3cbf15ed08ed9a1293c14eee935578017c84cb40c752a285c7eaa4b03ec8c705ffe965a005a046ab74e49d63e543191bde2f805ba1e8923c7cda11242393a84877ad53dd2a4d7e15355612aa607ffb57eed036b6702b550a2e67dc6431d3fbbca21bbdfc080214d17b8dae4959f3c097a3537701e8667eb329bfc577b57e764100eda592a41f9993e8288a769baa66937db740456a94a425d83af43f3208a82dd1f9bf57696fe627a9e385696a2d07985fb4a3a35f48dd915b9b145b4fefc0868f902b2900cfac093161251e048b741c6e6027a4e8cad0a842cb9f1ddaa1d3b4bad23012ced44a298d2f183fe0a90bfd44dd9b13298c33a30868af03b9e898488463df4f06a94d5bab22bd0c2e6f39ac65a9ec879e11f54a43a0fb57f8ea59d36eb8ce2b908b18c57259c1deccec80b25a48f2fd1b10e8064051dd82682a4465ab9a185d0d85498e9a923580400550f8bb438;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h346a49e61f219677ee74c3bf90d3cfd3b6a3cd6ab0221fc054414f8499aad39ea4228e24cf62894b80ec17e948bb9b865b5c79f7072ac39bdc44d9a20bb6c0ac90dde2539ad89c9d7b8d25905fc163af02b8d700bcb9997ecbba45a14bf05a8ec85395e98a0a7aefa31f1fe0fa73c045c5409577bd1fb9586646f55891cc5d7a2ae40b063ccb08ad2f51e2184fb460413cc1f9f5e2639c22d549467a9d04097b9d067bf5a072527233e240834d68e3d84b162d9bbbc34b27239d85248dc6f36d4839320f1a1405fed45d3e89300a0a5626ca5330cffd20a608ee23f2812bfefc75f6349d87ab24df35f01ff1356c98c6c7b41bb5a5a7722c3e097dc4f3271a576156cdd88ac58de0c4b1f3fead6416f97d8878d1561bee1b14dbf8e335b4efdf0b5fda9226717c0ec08b084f69a32e96a30dd0110a7a8c24439028acaeadd75e651f80c1793c7a982dab612a0d29f2d6704893e5707d71a695cfc801c9a4bae6cb34f8e0b79c0649131115bfea899825aa35960b778fe03bb0be9915541886f67f722a3641699df697c0a1a0bc6c0af3458b7a025c654d7478b44f83541dee4da22be88a1d9416a382a5d618e33e2270adb87aaabf11955e9b97daf60bc73615ae7aa0a878d01118ef634c6c729f448c7cdbd63a11d967c50e7bc28f0215d2c2bdb04587424ec4068e647c945af406c9660c702be60d73f36c0920a9b98dce408f50f9bf1a44a97ff207dfde187172d3cc4ae713dbcd07de70420f3b6ad8a208d215922b3bc9eb73122761530af4ba734422ba7dc9690440df94d18cfab006b75d1bdb57eba44e5490c59ef29b825e76c9874cc5bad03ae886d35d347a25f9d13cc15e6643ddd0e3267647a89c725e12a08508e46093f29601511c610bc2e86e239739b693b402ab519eefd274355ce95088caf545a725c2b58be11d52fb455c966342c586ba7ee3c64733d3700e4f407825af476fcba40abb01609565a8db827b20d1607b9633441aa4b94c66882250955c2220cc92d7b6d2ea745a6c6e24d9f6289bf736d668da452ce5ef81567b46ba562c033122212982065383d51869a7ad246823ad1c5e601609e4594740003f6eabc810594dd32e5a827697004c42b7f5d7db19ff236b36e420a4feb5cec2dd7cb43e401f6c3efb5c2530ecac6fd68d797fa29b52b934ce1895b37ba3fb3e1fa5005ce0e5aacb85344bc90001f9b23a04f28517dd7357378e21e50a3d8a69d8e2210664bfe77876df88f8998f23afb95d6084114b8192b3c36d72f19b5c65aad33345090d17cc1d9e4d4bfa63960e1ff74ce9a01cb07480bd93c4fd392e163df190e866e947d696d997db905cb4e028526504293c4f34b6d671706feb18eb7cb94b77ff0cc64550c8bb8ba9879fcc3762643d44d669aeb7240fd3af0f509976fe0c031ba5bb30f58a82d4a47185c92a9626dd8769c6b62c48dfb21487704516fd7c6546bfb7b09b39688881aabd3e79546d80f882b3250b30ca9a1942b66ecf3cd57c5e8995339a7d477694adfe3845bce89d42be26a2fb1d6c3000197926288342eab06910774fb5d7b25313b83488037acbb072bbc983dedf786c4710f4b2989d40bc555a5a7cc14b45da6cb9fa56be3d168d8de510c1b64b22457a12e329a1a75d639795d3a49838262d2ac139ea9eccc18c30d86dd17b8d581e6074809449936a42d7eae59b724cddda56f425ca9045a2909100940c916799b78c4176faa2aa712d79ab2be87be877dcdfa9e335166313c8f32960da2b90ea93423233ebbbbd31f15453e26569ea3b5671e3e7e9dab29c2dc1a59d353fa69f4d29e3db22;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3956bda81d3f33dcbab1e63b89bc8b55593d9ba14b3af2367423189ce2bfdfb1d5be1e25379a57bd6474807a3dddc45218f707e026d94bbbc3ace90d6c31e174441e187c4ba2633cc215d6d773be611123ebe31aa42ce8e0c8ed0701d16f0e3a372b28afe2dd8ce1490e02b13b17bf5f0ed13f20578665d796ecb7c01b328a57969603e00a1badd9280725b90101b0e360e23d15e99bc2f99cc1b2b6c672287680da83c68ce334b9ae9ab7ca6e6f9a9903fd83dfcc3f1f4978328f4115b4a6ceea7530bce1fdb9d24640452978824b8b8dd526bc7e3d040c7891df83da797bc8f32e1b55a9721cd320d93c4ac70f5b8aeae5d681d4b25b6add19eac8afb8d8edba6cd0033f8cec5191f8c38c242a1a26701ce36d7b881e28182415773eab8f31a2931ba250b22baa92cb14c4eea51121f870090f242993cb561afd3743da350b88d060d9b2ca6b38ca2228e7278202121272f6df404f815fb60547465ea4b546cc868156c054d4766901571eaa85e38781d35e8c258723abc7ce2a34a7c2d315e8378ae2098f11d460a40c975e251268b8a5653fe03e703c111fa79ce76ed54dca295bd0d8525c924d2239e7657ac613884f85c7731bada8e04046d2d6b8b909680a393afe7fffdbcaca28416a6c61e6a72445ae1be7e00b05ec7d38968ae128657d20b651eac9836235cd438b9ecfc2fd59670e41172f2f1857842dc47407a0fee900835f2db3f7cc2b7002c3ca6c3323b60f3e25ed784284f3fa4b3b2a6a11ae55caa19ac25c6b51821af334822f95d36a8cf1fc0f27df172bb4694c872cb809545b79f90f457e776babfb5a3bcbfea0c085397b132cb4fd915c15401ca23d7a1ba7dd059e0baa0d741313c0b316d40e6eaa17fb66949a574b8480dbd74c9ac8fabdc4f67bc7684757f9542c3b44c77d99fae109df46e95877721d7c3ea1ec15f22dc381515e69e5830aebc84f7773e7cdfd328e6b3818bd550fd3b8d5ddd982a491ceb126344634301e2a203378a56c4b75dd655eb7ad0cdb7be446ac0f92b731abf613e3d445110b1a2a3c7373fed58939b19504c8aee956ffaa28de4a45061e7fa608b6b007c79632b8febc65608ef6fdc30fe56173f46c41df449c55da4d97c5b5176aff476cc4f036b061a59eb81253668c57cb476eafdda17a08d18e3ab66e30484ea639d50d292da67f81632191ba230a80bbc658cd6b9b057484903d6265eea58a8375405c852b09ee899ae64e7171d750f9cffb10f907d2fa9ae543889a18a52e3dfb3d7e2fa9caa53f6a2e077316793cb602a8e1d3728e33be86371dc8c4039613382916a47dc24969e688d2aa1a6a453bbc836fc4f608587ed886509c36ae8eb824fc2cba32ff24ae0072f5d053821bd9927f3be5c8d008533d214b703106a1b4db280d668503fe9181a14ff5619888e18e3368b270d38840191efebcf9e199be37eccb56e0fda3fb8f8143a02779dc1849d4f5a6ac480e2812e42082a78d2c9adf120b0fca398ac7fb2f0cb8a16c7e83411489742b747a57b858fed503df6c53ffabb4afaeed94cadd67377f51e9a1a42f95a9d55fe08640cba5b6dfcd4c4f9fab2859da05ea076eca06ed882bfaeb485f96d54603d1616059b14ae95b6a8c1aeb71a4bd0e0236e92cc4354709c408dcb608743a70c50f9598e4fa497cfd25e4556692e67c3298863c1627a7adb435faecf4d3059f4a895bbec799d019b49072b437c856399bec9fc0623a5ea5493a7546da054a93a4ff9352e2b1af16681ddaacbfc466e7291a753ecf30c97d1f0373c3abd0a0cd279b6bb165b3b4ed806c2c9c533ac8ffa4a6936d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hce2fa324cbd252870a37b5258d075c3cf1b2657fde8b8c8222880bf40754e52b7fef222ef6c15e0702ef73bdeda5b6bf37fbfd7bdd7cd774105a7a5b5340b802953b55ad44969904b5ed42d220a8203fa171004f579b187be47ad390b269683aac255a78f238940bd7050264a855c0190c9bc5d82fa188ce14d68854785466f3d58725c35f2127d53034f5b22aee3158c91045d25f05fb0b9e3a4b4affa2a74c8af178f8637b845e8770cbe57652273ac9fc6cf72d2ed1c4f1710815396feaca44d654f53d23f2df9d19ab002b1d8f67dae0b77892b66621f0fbb329f7dd8f325b79552bea79f4f55e971a1b48d98456173c2763bfc9fdd0b2d56bbc844c0afbcfba38614f0dff50887ad5d04dc43cad61259f01216b6e153070f582afe0f21a77264543b4bd4a30f44a63be48ef52a29d8d1a3597a380a100885f17c9338bea38ea7bcb3d2ed057b5b4b467d4b211e95565212131fcc38d9a5da35922411aff80115fb927cfc1b0a6d513f935e6598b74905d9b8beefbb16436e9578d83cee71f282062960e12a5d0570f786aac2613d5ed23a5ef623794008eff7b9cfa0f2f4d57a855ffea0189fc68222375c6ea695997a8a9420dabcf0ff14aa675b2455a00a42353442041490b109b71791b23c4e4a0a32d6bf5463708ee39582b6d34f314acbafda1d40409dbacf33f3c94d906f73657a0904c16e8b0d77a553a46465ecb4ae196799606e0777d43f64db65c3227238a5a0f4f44687a0dee78adf95f4a5b177a8e1357c7f6c08030a22c391494a4f1fbc627735e0429780dabd0e1bdf8f43d841236252ae20e89042903c079a1ce6ddd616224d6ad4535d4f7a4196e516f1eb611288847280c172903d827803a303fc34df67e06f04b33801af237188b8ee60fe166418bc679c0447e3648c1be0893821f754a1d5ac8aa75ee782e363b5d434eeab9de30d157951e2e6f99e62869241d21a085cf087c5e31cfcc413f8368e838ec61867695c7fed4befe605070146e2f378ea9f74b769092e0c12420270b82b1fef384e81de9370dbc4adccff4e1927799504238e5aa7f58dcbc0baa2af9f5b72f67e838e0fba25e76653bcc175b7a5c86da51779dc7f5f6c33e45ce8578fbcb5025e177840b6ae7bdc3c055a230d4ad4366bc15190a7dc43246e0dead3252f1d6e36dac0cc458a806b8c95541f7686c5eb964d33ff9dece108539e3777eef0d08a859979d7a5cc4073928aa86f5656e8d65ce507b4907ce67ad11443a5edc0a718b6fdcf46bee2d9019e09d3b46c0100e8a854d1b3a0dc24e0339cd48754f92b46619b7efbc3a8038dc7977eeb8dea8941cadaab1f6a8c3f8f838a14b262fd89fe8c13669631e5c80e88e2bcbda120850a3fce3074b7675409e38b3882a0c56bc55b6bc2ab03c6f2c101e372e1c5736fbdbc26cd469cdef01344e4ef2d4e1c28f2b642b8b9d5a4a18c0b99c215eb97ab066fb32b2975604a0e76f17c4fc0fbca04ef5d3adba1ec9b36b5fc0b2950fc25a61947675cd9a26b3e075c609b4b616db1bd4bd5325ed3af4d8a6bcc197a0475175b7a992542ecb5c456e85ed1277610b5954726ecf0cfad53d9c77144cc8bb7dc5e4b54a83512ee25223256266fd9b3207b1c37a76a2092b375ff885b02ee445f1290550c5e01dfe75c7be8e0ec3aa4b0a84a3fe113b42cae2a5524121a62c1e4883f4cb987c038fc64ca4f1e665a9d694006c1f35236c66a108a05f616e52aa70e647e8f26ca1e78eb22d4752ba061318715915780ad808ac49884d6c9a7bc67f244603094ba86fbd5b1948196ddfb120295bc91d3b95d064255366;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9ce56296502fbf5842b96449074619fc79019c4b5c09c028211d661192f0fa77e1f93744d063d2081d6263040e0394e58f445a1d90e8394941c29e3330bc6950a011a178f6e2ee97a52e5ff4b6e0829713f32e77ed93229c7ca22a62106ee64830cd01425cfa52de8d13028357290817c66ef8bf5006d773511a5131c447f97268b64646f2950886dc50c362372aec2722c35cc2b34f72fb3562a7a52fda88057d5e62afbe86391ad79d07c9216f6fea83c055c40e05a6338c8845041fd6f68c32300bf53ae89b9fe0b7b03f9678f17fa66c4581a6a698c2b795f61317fafe5ef80ed3473c526f39d2086925a5d76a106dec681a53f646b451221930d884fded97a1e96a6f12e9d3497766d5bb47bcb4b4f173cd4d540fbb0dd69aa4e7f369d18bfff73eba65c90a706787728b3a3a348b7531b3ff5df4cc373fa0dc93aedab13342065681672f4f2aea4e2b19c1bb5e815c677e9773f0b7c333abcaac1349ebd2417835cfdd7604493786b3d8d4023d16d83eacfeb4f728b33bf3191d742e4adf7ed1b4fc8321b3c4b6650f7052a4649d9dee8cea3015031bd2eaa35aefd2d2d3013fff9d506efbc73896ecd30fba0bac621b5b006fb93a1dc48e8d92a58d63b2431e32f6aee093ac20135cdfb70e7e52af31f3d0e83a497cd74f7cfb436578634b57b9796d06d82e571ed6d6e25c8ae627ca3730e514a358a10a663f33b9a8b20fa93b8017ddce0068963a74fc1846fb6106edec03c93de991865dbeb7658d405efde4a27f6a93ca79f200f8f2ff20c961fc0a5ad93da1635ad3e9acfffe436d46e0e1414c2f6a32c4defd68b7230e897a9ca40ed1c83aa78cb7f1e204c2210f259ea291c58ee1c9f9b2dc1784ed1fbb24fc69d95441b1ef6b275611fe81748827b1dc134d6a0917db28d48b8da6a3d5e5eb1ac874cb0127c992a0ecbbfcfd11c844829abd6f5cd25462da150407c8b542a322ade298b1f7b96749c566779d7b8dc4ee3968af4d1080244c62dd6fc6524f4cf6b6dec59cde1779c863c7378c0d8b3604899f7968d2ae1aa893f3028bf6b012520ed7a347b6a84ff8db735c95b03c5b9a16b78f638d629608d0181abf20677463e385dd5c22cd31947d0b346798dee1674b298b18a53412bb2556c31ce7280934cb9f85ec84362fd5e2db255dc01fc7e91aae033d22ec089d1adc996b2be3a31ac18b4f9d15ecccc626c0129adfa8f6f7198cd23d75884b443c513438171791840b5d75533b848d62dcc877766b45dd74aac4b855e339d4b4e84e28b7e6571fb26920941d24dffaaf9c03d3c3fed82fe44c5684a42ab79529c0b9c60300d0876ab76b70be8ec6cd7c4f5d79a5b7c4fa7ef932b411201177f68fe4c90055b3622ca95c81d16210ebceb3762b41d66467a7f1c148062c021072d3120033b5a3f47fc56daa93d790f9ced31d636af496ca95c035b82e91825374f038f95084a6278991fa660704a070a963c8556dc7998ff47530ee2af793bef06d33e6f2b51b2e8e0d240512ecb624e1b82bc39d3c734d0794b00075c136998d087e3d53584d8062e405c12a53ebfea0bef05944a54a7989285db8e563328d6f4818cad9ab503f04b3c0e6935192a02a4c16c20b3e43a6050deade931364b4c35724f58d072b589efc23eabc19beb9f26abf5a97ae25b518f39ef07ee9b2369891bca344535a1fea01fd8205928d4440a11d67f671d6243b6e8ed4a587fbd84902a912641f76a1d8ae819c1aa63c37a7e493b1c3688d9d3fb73633afd45fade497549a9ac51afbf21c1c5ff1207bb2131ccdf4390004c7fdc6afaeea2c97d04e83552312;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4462b1d7a819150d8a8a6436e647ba3033ad8e15409fb914fe274751c1b5f957a286f59728afadf9fbf2852a9c5f9f61fbc78e79888ec6d5c79223e5afa70ab423a1b7b888e4955e580afb7aba0937ac7f5f21bcae70bd467a7b1d535c880adf47ee8434ab6eac8d567d470b83e7dbe6fe6429db80538158c8705786a7ef75247f59afe659ec8006530f102ebcada69ad6c67b27c2f034e9328bc6fa79144c1c18c9ba9eb08cc66615b476ee494f992d75ade898001a6980fdbceb260181f46e5cd4a33ac8c9b6b3fc005e39d1ced93a04848836a0ce90fe91db8c7d63948acc5294a4eb048155fa29539bbedd339aedff59d16532845e2356d85734d6b1aebdb3b8e9d49b0da5b01ce072496f9fda8425899553478f4290e826af18af98ccb18e5e63f0d5ba45e69eeac3fc0b2a1da040a2f47d9750ee59c82a0a93a61589501b1d0115b51744bc33c27a058875a2f548c2d7ddb8d6620eb6f4ba75d4e62c07f167c990f3e8b89a48639b083e7271f32761f97226358d2df29e29ce574618a61e1f9fb92079d844c8c0b6a7685ebd81de3d406e5557de677355ef9bce17facd35e31483e3bba4fff8bb84470235556c4ed5882e8d246d6031bc768192c16ab65de5570a97c3f3e8e8680391224afc6a06b476baf6811ea952ec28c912ae30cc10a70d46f289b25c2548666990c1cf4dedd548a1f0061063aa0ed1fb348d70be7e284ddb092934cc01c2b91a2e94a206cce431ff039f569f8e0b9d350c1fb3498fd0d0e6867c5241eec7b29b9e907c22111afb41a97f993d86b7aad8bb6ee72b1c872aab17e444b87c848f4c46e9aef4a552aa78ac3c3d4d93d1de760ebebeb245481a50bc96b2fc38d6d6d60fd18e3242f7955123f41985f0f01d32cc2411401aee319725d6260477dfb326975b51246334e51471e87b971493b0980460c80ba3c36ecd27f5d2237002a8686f4c458ef3ba99b9bb16f53a950cab8c75bac8c16e890deaabe78fb7e3943141823f0cf2726beb47a996d681582c73b20f01b4c3f548176aabc061bda293f7821f2840159ce5ba25266711168dc7777dc19ec176e48933b8291fa4fbd3701fe69a532d13e03d9fb71c6dbf074e12550834aa79110f27a1039be914b63647842729596712375ca08f575099fc1fe7ad0713dba1c154806eecba5144b51a9825b31e8ac695a570933f9888d809e53cd73fb6098c06d1596f25ebbce8a658eed3c47ff197565e70839bda419f241189bc7911c62dc7d081e8aa0223cdba7487e85aa904b1f4fe28fe9d51a81a6042429bc5ff9315ab0cb894cc9507503e7a9624d51ca46b048a15e8f9a9f8e3ea0edcd9d5114c66865f9bfbea97f9b1718261c33dc1405fb98aaa6ee33d00aa623c6807cfc94e253736f9f728a8ebe240d36596c4ec473bab393a8d7290a3afa3363937069f413d6b834fe7027d74b8392af81e28c121c0a160edda6dc4e87a28e1f57a666f4c7c17d4c91c2d7e0e66b044e76f2b7e17fbfc86bd10c5c5d5f556c1221b87d55cacf4a3debee524f7ec3eb0f8bdb0f9299c821ea802a5b114c72c4e47ef699c0c2e5f726d76c44cca4f3f548b8cbd672d21968ecf9cd07b8d5fb3989ffe1e27438f647f5ea90365451ee224c319239978258193b3a0fdb6a23d8b65fc643e6b31bdf4768ec2c5e1634cd7e0db056c2385f1487e1ac56a6556de5214e948b0497b98492c28c26d122b438a277d99ea2878d8c3c20a2e79b3ba47706163b1438f0bec93e6629efcf627ac3839defa56926ce58a8e8a6406d5e004d551d3fb55b62efae1d7c9bb3549d4b0bbcff4ad2e8d633981;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h90c63a7b9947468f7bff83513e388f26dd60829a3676e8a4bec5b1e0abdaec51f8a6ff935d4c851c634c597bfcce7fdc5513ba1a46313e67fd8000f5b33ac0c9a4c5eaa78225cb83b3072e877a37cde86b4469238ab131d9029b6a19fb19b148ab06936aaaba1b13dd7ccb0af3fda71fc3e73a3b2c7afbc94c605c829158cd57a3156d4136a1064ae3b99d7b246c38c028688cd0130eb4aa87bfe961cc2544223f6c8c7bc5a057c64ca6143b63ee986739cf3e7b4f0c4a99e85e2d835494f026f068987e7a2f2ff808bcefcb51e0cbaf94750a42db7ffae8e7003bf8f97bdb62956791bca82c93cef92a0ea7f41581c3439e91e99874dd9f53f2b4db00300a69211f0f2f03af43dc8089675fcdfd902dce68a8b65dcc23cc6cd63b395118721dc2ddec263f810f609417685d0c7b4a554d074bc33ca564c2d16bd7b906bc4f9244ab67d37e67490e553b16f18597c50bf0bca5babdc9fbe0644b2bc3d45d06933c6955bd9a095a3cd1f121f42a413974c92f3e9e4d9163a8dc1b21053604ce2f2eee3a76dc246d9fb6120c1deee96b58527330489d11c4d96ac6a8b2c3fb9cb39a700a4036dc76c4c638525c4e6a45c24d8e6abea70962f5cb4c154c2828a52821cb8806d7424dc732511b7336f715c8fa0ff88bfad8052e77aaeccc1b5ac901bba59d6fd055468a0d9c32aa0039cdadc74d3d87f064e59711e352025d58df66fb94d8315376dea0da865ce5543b6b2cabd4430ff359ae7620dbb1c446193d323291a7652476b7f3e0c120f9e55562c165c29d2620c75f2cdc0fcfb0c9c19d5ab40917fbb1624032ef489f40eb39b47380d4cd8d3d3518654623e086c387c93a3240d91fbf18f70149a4601555853a2ef415d783b1b817967b338e83eab40c3c81e363ed284f635e40eead58cdfc9a3571d91c485be61255c0da5cc0ec419bca468aa1b1c6450bd0ce0b1112a7089ddbfdc57da2e6ee8bbe9823360c2dac7652019669f24d2a2d5fa6157b07dff7e871cba1601cecd1530d02478c83dadbee94eb7fefe5597f756e8f60f454ce7e2b55ae3cf43b8855826b6d8f39e93e3289943b932203bbccbaad049e2e3032b1c08e91778dbacf3d8ebec49f47c25210840f7cb3308f0c2fbb998af929278f5e7380187a893c89747e8a5ebf4bcc901f2a159da6d41ba449f172e306470577cf08d8d96cc39785cfe24a1f98de0a7dae561d105bd49dddae26a5c3036982c5a2c11cb3c8b72e5c43278ca56094d9a7eba72577d15912e12f65cc6d36b5ced66de1fcdf0036c3ce79fa46e97ab8b59be18036fdabefd155b2964e105f2130ba250a6968fa211660389f520dfc13df21cbc228bc1a93054287f0cffba55676f38aad242e3fe44d2a7c97420771566696981ccd6f563b95a23c94931faae883c4bad32c60a5b0b892ac96993569a8e40f06a86a8f5770b164c7a6b41637d8007a61f80988e75e39f093e614e2d6c273f07a989564bd5b215690ba91463bfe0a34d929a64224d48fdc22aa2c655ed53ce357088a91664b9cb7cad178158775e77c1f4b9f63be63b9c56f99560907f227c6a84405ed1f365388242ed67af7d613449898fa80f313cbab7c138ad9849c52c91bd4d00abe4bdfe9f6b3ec651a70d3fb229eb459991d6f433f9fc27c632bff07cf9d423c43ab38b942248d4072d4940614b60421943276f95877f286e0c246a64252c0708f62087ad05a2e18dc7a87c99fb1a24bead416dfdbf4d0f1b42ae8e11cb884cd2955821921ec6b81ab521e1b1a45052481fa6b14b0044264dbec13dcd4b262378ae76a5801f071f7424d46fba0ed9b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcf1b8f5304e62d9249c42988ab7b3c1defe4a78a2fee95b5152f839c6b8d08b486c214a99732e5be06e7a1d8537635c3f661d03f21e7f7be8cd5644378799dbd5e57dbf59b5c7f495cbb2fc926f884ad18b0e915ad948193d072604eea785932b25e275e7ef7d2a1435715783160a7e3b8003abf904db593208987c983edee3fa46d1e3778823919a79d2988fdabd6506258436dbd0f6a147f9d0b3716fdbc8b34b18f9061e7d82e2967e33ca13e5bc94c3a951ccce7c6d97b67629432c59061ade267025095bbf5408cbd1688df1270652cfe0e78504e000f762bbdbc54b55ad4c4600ee73067f6557f99f1d2ab0a7bbf02d8221b8bde579e437994380fb78428058d33fc3b6425860d9e0d7ca78fe4e046013704bfc41ae7bda035afd5a67e5b5561c4ed0b2db72dca89e5fd72ff94c71dcc57c88cea212bffc075600d4edd334bcc32d3ffb0b89ebfdadfc6ce24b6ff76c578623385bd4bc3d003679ddcaf8121836417564706c971c729c62e052c75dc76daec0a35e33b385680b8971707fa98806bd3d90f3a8df8ee1653a96dc7661d49248d23150a8ca814947a1d699d857e9b88affe201df8a13ab8d32984a562ee64e60d05b0dd1f3950e42356c9c11abae6afc658e675bd79add7369999416844972ee9a869878a2982c60041c3b0bc0e7aa5d6591da502e51720dec512da7cabca9b6f4712f31e153b0c60540b72823dc60c7014886a433b34a7c6beea7011d24ba99a83f20f404a6468912a1d2e562fd2515798663af75f18f4e21ec2d03864334e3fb0d375b96e582f4f84c1b9c099033f69acfdd1447943c019a7ca6defaf2cf0139d5524c2a5424118b006f16356c115235d191e5e818d82f7a34c0c5b5049b3401ea8f450015c56337fc7becaa125b3e46d34ac27f9c73112acafdcf1da3764cd7c1c18e64beefda8a200d431167831fef4e11c1b7317fc0c30f5c976e50001009fed53de18e123e3328ef84e35ebcf2a894c17684b57256f810876c869fe40452e8194a090d39bb22343ec312abf6eabfb9d34a0fc86b51760feb90d1ba87fd120c48452669eb5e382b7c96f41b22c394faf6af12fd8868840f6d86630753393403606144deee03eae1e1422055ff468a1358b03740f160c90e3731db532d14d9b28ec0b0ed0601336341d5b0c762eee0aea3cf2a4d2d5f7e05cf3b52dbb03ecda50191ceeb71cc58d8175e77a457f61bfa9f79e515d93f267efcb868cea30d5cfa1cd6b87d2b6c4f9822580f2af48c5672e66069224e4bea2d17938ec3910155807669c63a94099d9b67a5d51e0b276aa0ca8458105fae815c80dc87c62cf3e93f5b366fd45fbdd9ad0c30a29adecd3f625a62f8b55904e177bdfb82906b5870c4508c3e1e4dcc07c4cf4fc83a2bdc535305becc342ad551a034443d41dd9e7bd4594a8071554405efbed6b3a584d8abdf19d3af9e9cc2ed484c0463fbeda4ca66e126488064ab944078adbb68e98255ddc3c258e48134da40b67fa2102d662bec16d6f5736b23d31ab2d68cb1027fabf52bc2427e765b38e1f743c96a51aec7810dc3d7ef176d7e9515d0443dd4e19fd631966b14d0b1fdb06263864066e1977315c8bb41d6d8bc9a36e6ead5828088401f4ff1c51c2d760858047576e9b5c1460ae844793c36e2366cc6115a471b8f52fd8705f37a570b33e7ef16aa5823673748ccd6988559be6cc2075174cd29e253eae8038579b26af846dff7f9a1491da6d1baded77d98ac593b09f420a94e447b03b43672e08a59456c1ee5a788407175d78e886209b69b919f3007e48068b8837946f65c0a35a0ca87e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha37e9af8616f41524f50e422ab17807bc304827146e23f457fc15d6ecb3046858496094a83cd468392d6c76c2ba25d55590492a6a77f6ab750619414fbcf2d8dafdb7aa8d6219daa5005412d25600d2e3d4c92ea20c003189e24ecd195ed792f5a182d8176ec2aa4f4381f44e8aea91a6b1f92d3d5174aa84406eb81cae0ed25acf3dcca1203ed7f18f1e9c2676fb4e4b15c2e637efc96aa3165ea0bdbfce44006eebba711b9733a867ce45fe8414fc9b7bd27b6f06361b0e9c30ea265e5c03767e7ab963dc8a1d41b21bceda61255033d1dcf47b6ac1daeeab98a2c606203c801292a9952d5b2b95866563ede94a8567fe3ac458adf0b40347082fb7d47428468e8aeb9f7442601a41b6d104ec6e096b00d92c824ff771e4a1eedcaf98b89b5f6e6d9dced5ed1dade985c734d03e3829650924ce8c8c76c57e3feb050d330e81752dc3ba1ca0df4ce5820d45ad3a7696e53b922eaec3709c968147636837384680ece62fb243d959cc16cd342bf4db6d79c5d8fe87d5f396dbbaeef56845c5be26dea2f80e1d119884c4c22779edb443cab41da20793938b984b33ecf87216ed6988b0d4d7f7d7056932ae3f4d35a7ad2beef0c4e0efe82265b0f861121274c007589a2726fc759d94802f0121bf98bddd09c4cad304c9b29a905a1ef33d759cf0c3bbe7a3203a8718acab573b64d1ee92a372c11c5fb46151c8109bbc91818c1140b20e97e8d5a2db40e6e4d1ac258e222acd7804c59097466ac8706e0f8081f56db5e21a9321877505530d130fc6831962982eae04e447349fef323501e3056aac562b3e1813bdd904935cc81f1fa4e4cd7607a30676d7afd82a283f1e3c27a90eeca41eee8c0f9560372a760e4c10ff40264d5ecfac1305a992c459854e761ffa72b332bc07dd4360965aee6207beb7236ec42ed1c529c5c03b25624525e535343c0b79385bfc5d7d9711db645ed37a9a1c8868297a19a11c443cb7f254891652d47bcedc0e2c9c98ff6c7194bcf36f7582770092d39b4ef31f9d47a7cec6329bbc56f62f23ead579771df8d44f3004ae5c82a3ccd1024406698bd34797a507a6706f58adaf2cbec68db44f78371865f94d6d2872d8d8032dbaa1622532a266646657085e2396ea6f3a27f55b07511a33ab2f9dcd290840906d09c6fd5b49bc83ccdb49b2ebb742d199be9849ed67e4a40c38228beabfc165b961ab1579ba0f1908612e9a39620b31a8626e47b703bf1938334555a358c16cd6c4137945c1db5991c81aa913f7c7db119cb38acf9dbfaea5e27ec13a89db87558e754e26b588f59f260b7b7b8e071a906eeb76d48ee41ea83b13698f8b553f256630fcfbc5925ede12a43cd3e3a0691ea4ec6c9c7acc8d5c2bd63ca34dbc344d19af19ad8a131e7eaa10a361f7c6c147486d4ab8f3072ac746765eaf5bb0fa257315901ad71ac1198309d4bba0200f57c5b64fff3ebc0fd2ee35268f045676572478b6b31bb7aef1fad6421f5e905bf98ad0b8b22e8c1c2a7840ab3014d6ee2c9b54a47472021c503d7ee4492e72ba5fdf23daf5348e5d14994fe395d30ccb1e8d5eda0e560a2b60e87caf1c9f3fc4787bf56bde43c1c3f0f8577a0f3d0a8bd529bc1683c430eaebebeb5392ee62b17badd4836ec7758c3c184de633df460e7ef6323699d65602070bb7cb4dc8373da4690a96d2b7ac49af6b32d80169f89495b74049be9889dd08b424cc1f093293730c29df7da574e3d49a3cf51666f76bc7b34d9776b85d82df2e139f181b1a5534ae4e12551482c688413ca73637ab89803db1147be69ab74fb80b6c5cc439b5d8a3e711ffe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5e0eafb12747c24a81d1d5acfe9e2d3df151098cb0d4ced3346f902577a02833466922ea7afbcdfb1f0495164c7e9f37643c8c84f18c0a7bc99ea75bdf515af9bb7e625dfdb94b8761877affa9da2c248feae44d4e1b8c79ab215e5c005b67851bf1ce02eb42751908a2cea6ed398af57a5bbcec95a129bf36cdd5f695b621c667de09941cf1a5fe67c900163bb585156a9a769e4a390690c4a0499b156cd7ce0f5b5ed44558ae4d8fd95bde5c7230ea3e38695f18c696a90cb4d5e1965711e20e29da6f9264b7f685dafa276a3f1130fa2ce3a82be28a181010be01453269e871397ce90fec50ba7b701497c7283c7cc2deff57dcd5665ea15991c8a2ec6ab343339404ad4f8827dafd49d1ac837fb8ea59a8b75520aa346a2cfb1962a02fe4f81b37ed4b98320bef81801eeda66305703c2bdf21a1a448665bc0c769f2b93278ef1e4ab22c1a512563a7d2113ce8a927838da7dec6927c253579db81deeb3bb4025f7e9366ccdb1d322b8dca94b9a6fcfa436cb4390e35e212885aab40db590af5ef28b93934de95d6115721c18eb1a570489007a83a96243debdb4f62a7edb16ad70c37926921406273d186e89fbaa0d8380c6ed43bf90bf2edd90057376f86ce03677c6d2495a22dcb7179982ed2bac59b7d23fd8b7341b29e46e7154e7b4f1c12e62abdbe15140e3f5c653cb53f47700a390668ac1f7cc042f26169c726405f61360b567e5eafa92311167ba4cadd6b709c779cc3d921263ec3b2937b967565928ce33009660a674846fcd3cd6965973add4b6a734e36b8d4440ba9a154362e49ef27d0119c55cf2ecc7eb1271011c4d3c439d368366427337ca865bc84ebd84665cedd632ac85a68b6589343a9d28ad23bc00ed0cd09fc5ca43881557938e8624aa22186a9fd691b228a007b745665c82888b12b5a57e5e3d9b605ed82eb477ad99a3e622b0d189a0f5c91d52cfe9d9e66b0524039f0afb9b8c754f68ff3552fbc0b3e722e8427edc85474f932c9412cff0a6ea39e0fbcb5e2d490bbac873692113b431416a78cb53b01b73935cc98b3de8b10897af8b57e3e61563c7ac3c1365b0e48d81fa68bd3680bffd4e4e72c30eaf438ee747ca23bfac2aa3619f1e3dfd4269a793ba9acc2da06885665c5e2a025ddae4e376b9cf846e644263d5e094c3d11a1c23a9460975c005bcb462965959e77a8426b8ddd58f6010bde493ca79ccd55abb5e91c7720b4971a4455d3915eefc9b880bb360a5a80543d04ee14c9bd97c7b1ae3f2eae75d1fde68bcf1819095d21ca8e49c89036d90a345900ee59774d00bf980ef9e61bd34c1e00435b078e3387c256a3a32e5d693856a1cd97784ee132de6b80fb0933815fe68c2aed4c2c87767596cde01c949463bf954e90c75ff328dd18e2279844c5fc30dd0d96ad2f9a44a19e912facb41373caa01dd26579f2110f92ee42a5b3b22dc245b4cbab4683e7cd49b5c540c46479ff0efe5afaead0e941c2a5910749c7e97bc97fd0f0a05529322e3cf9e3e7bebe66d54e9befe699942104c4222927218cbc923108167a8acdcfb0f418b25837a2e85617927fbaa024eeaa234e576cae180fce6459750f605a1a1fe655801f092d946e107ddd22a2dbede2316fb628d85eee91513722c59de9a4d49d99514bdb914f63999da7c0aea9c546e9005170d1afe8a0e18f3f590d006294c7f3895e33ee60afa02bd09d0e77e56d4bd6da41533e4df7a1e715032f5aa5118d5913bdfdf8d24ca7cf3dac9c215926a1c4002c74c6cf779e9fd461f5836144533bf20ae63425b40e0a6c9fe7c6c05848e7a89d704198a760;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb7d3a2a3ed5fe9ed3bbf769f0127a7f0d64be5699318eeaac4c0635f7f822132c35f0290f6df437f0b9e264e864b97234bc6b1116e944ddf73b632b3e467e7d474f1a63338e3f00eb5e297118c4e6f075069c7aa95e3849701d5ca225bb1c4cb9a2e26ea5c00af00b1136374f82fca9aef4c5189eb268ec92e548c88869338d33f998d18a5afce1ffdcce0ee291f4833a390d7aa559344bbbd3a26d26f7943535a1eeb0a687e1d4ed3d5c0fe55a6ec75934ad716eb2322325257886d90a6f2ee1e8fb485508e06696967e4621f122cb5fe4b7da597f4f78af6f4a0ee3e4b723032c3aaf973763bcbcc4af273eaec002d56fcd41875baf610b9faf6922c51a80c6224d26eacc41a044245e1f0edd9a26967cedda838fe84852052290bca9ea56430e4e97cd4c6339ded633263df742fd0835f9ae07b821ea2bf01d08b1f1c1337fc549e96c1f2eb6dbbab28a7ce179dfa2e7a4b548245fb94127dd11139189f5ad61b3e40613eaa54170ad1aa1ce38fa4a6efa84d8ef227f93fd87eff1891bcce6b6993840d59cb42d40e031a5b9d960eece5bae74e7ab4e7ef8713919ae0ebb22274be8c78e38e47edbdaf71c989d410a518c8d2698d1a235247d9fd4e70d95f2001222c187ba46c473b3e172c81f8f032183ab6dcc0cc535d331a374a5074164cd149fa4a06ef929dd5b7f68f71a84f64fa4560dd8e48c98444e8fac05aa7b96227c496a40b16c692fcbc5b936804c476224ff2372f68500fbd58b9fb23da8e190d68302c5a8bc2efc2b670e42d0f0f34b33d2cbaa63b8e0f9efaf00e088a867c59aff1c6760786ccb8cc88befd85ae63d7517fd82f431fec03921a4c231992880adf1545dd3a742ba5c9bbcf75046eb6761d14ce35893397a6c7065aa6ed648e29e219b002534701da412f753ed0be75f836e032979006eb6510a3fe0acbcd8c79c5f2d72cdbd7258232f9d7da9836d73b08111260579ce7a70e9de7443e0100ee68933d249200a2f5519a9e1570e8984af8056fdb550aac8a78e0c58f056b0612af0612801cb874fe0dc1553e77e7bde73d6a5f9a4f987decc30154063c228a4e0c7956d02a66ce9aa8180a9a23f588e9f6f50b917127d09481e0eb890a46575b590b0233541a09a7e27d886f87d1ab02eaa53580d9eb5b5e9ba9c143de51e03df63ea84d76c1ed8294849c1f79879cc01cf0b790ca422a1742c1161c8066b0f18419b780d8d3b854fca6578b099dbcd8d7e8c2d0b9d4853537c7f0f73b584e975eb84cbbd8017531baf5df5dc4ebf44a1bac78c2eba1764430ce6bbb6f3d49934b5dfe7c5a8ddf149dce401cd43b218f8632a966ab0548106e27215ee762309eb29d3e5e9aa0b3a4789fc3690d261f0573a1058f4d432e19205e20c30844218214ccf9c4e7983660420a0a39a16b50adb62838ce8d3d366989d880ee53ec7ecbadc9a2085740869a98c01c4f8fd3c92a51f171c31cc0288765a25ff592c294fb84048f5e4cd518b20512dfaee69b6ff808e0a868df675301c5ba89a7d875b730d6a0e63d6f856b06ce9a3ce5f18b1a3df02029864f701b4551e37f6023a0eaa8e9789d884aa035f4649c0364956f9ff75dab192deda44a58ae7b05b5bcbcf712898c0b25b43319657c12d3fa0a9a8d9520b0c17170eb7109dd5359073cb004c899681bd91c0c5c5e31b886e8d762e4d3917174e2a924787ee6e56a7f0b327f21ebd85d6c02da52a2e058108c49abd261c20198b38cc0217af2c125a64eeca9b7f8bbb9ee3d8513fbd435359bcf9b5445b939d11e1b851a4001c4cfe41eae0822a1c6f5525c0e6f4abbd4890be905;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h359339a50de79c2102d7dc7db74f4142f6c3246e2a29ba6a8cac5905cbb9eef23941d684ecb02a9e8108a712692c140daa4fb982615414096bc16419845e5e9305e80cf8fb4ad6fee05436bdbd49b3bd7f3529a048a3bf5b8e571cedaa473a039158422ecfa68b8606f934ba759ee476ce72bffc5e471865eb1b2a61b29b8c41e1ca1c45ca6dacd2b0b6d19ef277af1d3b368e3855e4c7bf806296b7bbaebc5d5707d2175aa36a46bd67db5a23094a7451688ce33e2ecf869f6816adf7ec79f37e4dd83127168217ba874ca3fb6a255b850bf2e5e21b7855eedc6e5eb5c1f49f723209c06324a34c0cfbba1c8d0c00e425cf093d3d6c59811eea3f15aefb02f4c8f61af5dcc3bd29c8ee6e7bca4704e4c6ae630881069da0bd3b506dd96df1916d28114bae59f3536d2b8bc6319f2eca5a5738bc62c4e6aeb330f1b3789f6c6e1a18ff91ce66d7b067722da101c0823c539cb6b2f005765a39b6f68fc81fa4989545a501f71bee54b0ed979d1542169dc86ed51d69b971dfc6310f717a9de8ed6b549ae3c16ff22667a56a042727e0ad46a0869abcacb021fd3b0a80e6a4ef55115877a92968c71a20d1cdb67ff7e65873d0415f6b31103decc12244505825af0acb261fa543a94a0a30714ef903193ad105e61d8ee60b6f926e73aec942dc397749ba054c32d70bcb7badf0b911a63aa74ed667042a298dffdc0f1dfd7489ec60662b9206d1ca757d79bc4264e940644e0d1ff56762b59a62ae03aa1a99ff9db6b180cf8d9d869d00e8099db3d607f69a7e6f51c868d3817ac4c9caf30acc80f6b0af64f6dc0fe9a52ff89de6970a4ca73808fb18f04d5ccf7e22d6fc7b4e61edbaefd29412e8f07c3c9d9767de08fb9f02c11b5dff568db31e02a33741b846b1a3a8691bd4b761f26f08d224541db8d7760fe49c677f8ee3834d5199a6b1801af5a6527ab704b8aeecee52b8276167bc9718859cbe8ced8c7b0b2d0da506f072311b9c4276abafa19c9a9ec517396d637c75119667cf10ca1dba062076e441da60158983d1b06c9d3c304c2acecaeab3692b18f088ccc877e573f153d90b371a40be2f3f30f959c5ea112f719af7ac69b478dbc3d767f679b29c83e75d20779222a9c7f2f38acbbd3b0190fad484dbcd78ea939292e60ef3ffe54d17ea0e4590ce8717cb01ce38a88448941bd4e77b2c7459f103b5ef9ba80328f5e2cd0a07d8dc24301fc8fe090edb9da43fb09fd13a885d2e74f736e821b75f35b229312d6a839fb213f4fab922727e6ddc058c7bfdf6905bc5830b3580537ece77be674d2456c3debc64b42db75af22c1d845f2fa2b988f72bfe0736f4a26f6d8bae3b6a863afd432757daa217b6236335d66975a6c45a91996e3958f9e05028607687256e2eda7db31ad48fdd294769151a300278f6869d3b45668baf1fb5f46c1952bbed9941e3d30cbbf83ef58eae4eea9ef2254c87ed1a81d0fa02013be32f64d101cc83fbf2f55489abf9d585337a11eeefda289d8214c70f1419952ddd82e64a9b0afa728e1dd01509efd4fa25e9eaa1a6130c8ab33da978f2057af7e61abe5c4131937266d9579db44339e88cc8017d4cc63bacc5e0657040330206d1c0a59edd7495617151f890ebf3dfeed38bcaf715b6e1c66fab69db9c3044d0ab8f0d0688a2844f8510c097d46449d63a064fbb6fb673d26ceea9d185d13186f2fad00938a306d04ad92782ce8577dfcf5a8fbb4f37f506f43d22382dcd11526caf7d0ac83e885d09b8283b6a2caf61ee67f064da0bf25151237ef3bcd4948f1225199b9aa9bbc12ffc3d7df4c19e90c00e6a3f38;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4fb334330f6fb58e408864c0c45b4647aa7ef412cf449192dbcf266018aa72bb761faf0eb9ba76a11398461d5037b5498fb1db3da8275e8b0a3a6d30414452e27f0fa9975710a962cbe1c3f4362669894a0c836414decfac1b4fd0ccf71ec61c1c34fd3669afa16c5f50718f393961556b97ca6a1069efc69d12fb268af25691b49ec9c49c8262aed2bbf21a6aaea010f278d91e1a895f3908350060b3971bfe89419d29ab9343502952c5612a2b18cdf057f38c443c1d5ea60289a92a2a3404134483c672fe4a3d31c41384fd201ffb5ea19e6180f39088f2e598f0925f228715e58f47a4e96fd9a12c2fad61487b11488e420ed904fe401484714ee333c2413a3244d2357fbecc1755410368557075d3e49963864fbfa1e78210e63f210b21fcbee6920444f4b39ad8860cf3455e5127d94ea3e0af6ee8e8ac5565e1870c550ffab70dddeb659aab27a7779aa253a34fe8bdb425d02b59d3244ae2cbf89767f24f6c8dba1b3f2b9c8be426ddef1c6ba18d8acd7bc8e91c2fbd7b0a8ac5ed57a7561cc74a269dd67ec87c2aad65781623893cbb5c926e672014082efad475a80876a5614b66b6c91d602b84f53955b908948f01c8e6ddbb8c971801c27aa6c1c8ce228e8aa5b7236eb271441642012b61fe33a019ff9764446dbaea4d38800814650aef91edd196ade7964c875c3b57f503777685413cd21933f3933b3861a3c719f8b00017ae7c00b461e62eff7377ce2e2993deb90ef64cf654b65a8098d5e353e05efc4812f4ff96e56a7328729d35a6472350fd36523b91938f60a567891c1f9702a05d628148ee499177b178767a3a5799cfd822a5b73411535b55dd8594f84b3a7c176ee3b88084612945da27fc4e98b1d92fe9ef998086cc8fa68bffc38d0d3e3422bce8d16fefb301a080d0af35b05d1f2cf4313d0e9dc4e04710ddd35b7860b3feee9e97491546a86a184b6d42727884680fca010ca5f84e1edfceb4c8ba31d2f03567dea5fda59b90e059063aee4a68d099e8548fd0ee7dd3579e4dc46ffa8620f6fed8e96b013a2d0622da63548fa0218aa7d18aef7453243cf2b8433d9f5dd101ae436673b5c415f6f33764a754ecd9fa64dba581a0cbb19e04e4d9f326d178f83864e91fd1f9d13d933ca029384b59dd96b41cdf8e0b9350599edecdfab5f3f2dc539b2a4611ea62c1cb61d98137e75b393135180fbb5a4b79d4aab192334b6f379190b9a12af570d269b04bf6f42338d621b9bb8bfb7a596e78725421630d34d302b2ce494f07d22c5b0b6c7ba67217da33ef9a255d954f2fddc1105b2186ea3463f8b1c2e8218775a9e4257488b5aab330d2e18fc85893304926377e52db4a950aa92ecd30e6b33d56f2f5567249bfaf1fc8e3e42c75bfbe50ab1f0658a6bec26d492ca3a7111059d1db5c28c7036b55eb0d9dc5fced0195727fec680fdf12d1ffef2d9f1e2c7bff8374194fb2efe0fd360eba01f5f39d239955b52624cfbff758f95386fab0a016c25e79159360f507729b3af32c0f3ea54a279dd27d5490fd5844b6bebdc0b9cf0bef7f53a2f098fc6cfe49678043185b929dd09e170dd5407c45e98075ba4c879808ceb176f2707020eb8cac2947b135f3bbe006186289b47afbd7cd78134547b8d63b579b05a9e1d669b3e3c0e3e5a611faf38ef530f74a28935f1437ba0834559c33ce1889d1d85ac30be06ef2587259086fe05ceffbcb131ebb921303671b7d036f351149e292e5eca336f052205f15f86de0955b973474f8ee632f82dca9a5dba780051f855eb9a4ea74045cd07443ca79424bd7b460d5aa83f302be9403;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3cf71a49ce96783a63bb844abe57da26bf5ff4d94c9abb2b5d9b49b874cb155a8757bfd799e148b8b4af5fe9f7e010e5cf5524b371f541f47470e18dceca76a89867e80f9084e77d0145619f02ff01ccc5a2fa0120306b8adce152477e2c8c9b0ca845271897f2e25c9cf25c3e94bf9fa97a3ea804390a729a9b3668279f7b66d185fab3b8d5ffc1228bfe3daf8db9842085cf359ede948f4dac0fffd8a8ce835158f2caca47917939ecc911cf9c810ec3021a8c3388d8216d4edac94b18df5fc7a1fd38c88e4bbcba2cd644a86d3bff1a0678f8b9b378b4abf75d4dbf85282692782c326047639570a06331a9778b7747ed382800f7b322d42aadacf336fa997d276694513915b545cb40700e01b12967b0ea88c7ddcee37bed572136a2765fd19ace85341b03eeeeb1518aa1a8f98dc60b4c31bdc21e5b391630ff2f253d15ed53bebe09b4cd760e6c3fb89c9c7cbb3f966a634554fb886c7c761e578cac3e5befb7c72c88c476a096c2d74d98ae4c14157262c7d9feadaec8035a4f6f9f25549452ee230152309593cb5a4778565fec73b7e055e9c40cdcdadad9f34534170f3a01c61153c42fe3dfef3945fb47ee886a11847607d9028e05568a01bae2a00e363f05758db36c5f971de84dd0288909fada797e37671eac3fcbacc96faeb2d2c8d564ec8a5096181132ca41892cd6f3c7a27d77a2b744928024f8bae8f9795265afd8fd2a47e83a9b422803c52c7c68d78b233b9d5cc7715ad3322e4a0df60ac72cde6cf7e17463af180f66560857533b3cfb6eb2b174b9038c2901f4cf4b62611f33701507454780c1a690d95e94862dd7203c6056cd8150ca936421dde46b32e9907afe2583468d7e9562a9d032f5fddcf0c1f3228bcfc575dc0d9f89d209610cd9a777ba72aae8e3fcdc832059e8e15bd7b24aaaff3f23d753c93e47b89b4a6c937da9f4beef0af43857464d7c906a2aa09e9a1933320cff36d302a341f30e5ae50cf85b40e5a91058324d56c898380b430f0379c715f720bcb4031808e5faea78926fe4848c4520b59842c75e8c26a129e8808d6f040ca8aa31442397f3f230597517054cd214d84f07bf8ee6bc36d7048723c37f6cd31cad440d0060c1dee604150d458222ed2112ff7b072f44e2a97f2c093bf5298e07e9a2bd87c3a36b2307208d227290262111f47787d959e6f8483e239d00b7d36db5a8ca7b8b8a84bcdcf7fe2ae54c3ac96e9201c32f7d5b4cc243c6668246b42602b6c28d8046b3b25eb95b6ecd77c9790c5e2ae4669228cc31d55db2e7a1c09ff72fb00a4a8202d8ea5a7d1c10f2a52bf0ac679ff1f39cb70a663c3b7e2944e42c9a0798c8ad999d435c7c2f08e8106be6453ed3b7c67a3c6f66e057c4fe530de231ca551c0d7e70a87835f6e3ead5aae63df1167df1ce7eabee68d7039930526c438dfcaef3babd19ad3a33ca4453ab45df9b8bb28a811bb6c2eb356af0a3aef2d5704cba4d3e2b280d245c04064e0f5ee2f778cc4b6d5a91738a1f7f0e056d02f3b2cf33aa498843312412c9521ba21f0e480202baf21143ca19bd13049a4235e887b62ad3513b3f69074d5af88764d5c0031965c1deda54e38cbf335dcc0ce6b86d2331a767bc3ce5c9952a21ecf02eea974d3d4ce1364e9830eef2785e213cbcc79337a496f8d5daf000a1a3d55b453bbe83590e9e774891001fd34d07d232ae1aaed6fea781721c255cb9a3c492eadb8eb61018ade1ed23f0e8ce8410773f6c1b550aa41e489f88da63a66b67138ea6ba99c56f9ab7d9049a74dde595a90351442cef94bdc86c5eca826331e1c4954a59df91;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h33dcd166638e22d94470255fbb9ed96484a9f70daae1c8affe235a6540453a65f796e334d7f6fe669e31dc7fbbf23e909f028bbd733b3f542e891883e45416313ebfb4be5ddcef72982318b04d730d4886a16d422bf916375cc5a1c4216abca3764935688e79b9f88cd1da01c7744348eabfa37545b2d6200afc36bc68da4fddcb0838e132f190481fb8e9867e9df379191b4d50a79a2812e212dc0294703e36ab21eb1e03a83b71beb0265082f5711b246037c67849c0f18c0dbdb4eeb39aa22fb31d59aa310623cf7074593a6e276ea3ffabc1741e99c170db2c2c8c5297faf562edb4149744053894070c4f1e3fd11c5605e2817cc109d6f4cd6f9b6f001e9311b1792eb66f27389affbcc924e5cefb6dc77ecab304cc9f3bc6222d6ee3b37a471f2bb5c51b6b2cbef41149ae52c0bbc8b49c8f18091a5808af3fa4c9acf2d4ccf2b0425b9e11c52d5c752f83d65d9f09b864d4a2b6501cee9fd498a246a90e1bf27ad0055b467b5851e794ea312876e66dfbee29eb102718d3eb166b2508514f310afc545ae228ff1a321d4a0eb4147eee3592c6fbd30bc3104f409743e8b673308e7f24188559fa9a2dd3183fdb21dde727a459638d1095065ebecf6b723a7bcd56ac8740620e650a997fc3529f15b10239fb7af3c1ad9d48862b523e0cfddb7ecfe9ca1ffa8cb1f993b700784a7d892be007ab1dee146165093b595ec6202c3405c7431410f536a65c790314510f4e82f9067a56bb7d47fb1455669f31ae02a71421ca4f112979f454c69ea6369bde326a4c85366943f64027bcaa5dce1f552fe13638c844e35e595b2c457dba17ec44bfd9a319f42eec40aa1554c356f7c13cf1b364bfe190d4d614e87df0e3f2cac79a981b345262d12cc39d6132e75d4f97f0cdcc60fa65776dad959267fdc2944f689c0a32acecce1b70f328afac5de5ff1b8a441f1556dfe840f2b63bf46fe93be24be7d566dc563426fc22a3c61323a7637315af3461ac3a7f3961fb60b12909e7090656c06279065ebde236dfe0589608336644bd2deacca39097e033275da13fdce61432c5c90e97adad855f466b5138aecd4c6d781d621be98baf1e794364ff28a989766c9b251cc3344f6b5a0a86583686aa7bf3dc130a90fabd6b63a1529074af1b2280da515f9a3dfcc5f19136f51ae18ac88083c411689aa27a3d2e0e830fa5f763cae5b1dffb8d70fbe7dca50d7abb22fd40ae12050912914f40f9c70202f3169f2154c557d6da6e9dac506bb07246355b4d954a1a651f17074c1f6450a88d4351810f3e29288f848a5901739251506e3e560bc3bb1e505a57fc026eb7e852a92764e9cde24ad38a70146cdc435f909f28c03ff02c555070a7ef0510b136cf20fdc0d0324f2be8712c122b1c1f34945cf0de8c693bbd3fe2c482125962aaa92a30716401ff48051fb761dc2a11ac7a6a138d1376db44eecf7f30dbbe323143a17b2a825e6b2dcee2f6b59e6611159849909330c84a17ac2c7431cd17627c5be2a86eb962b40310b4f93476058666b3808d29803422015b464919eddd2a4cd2cc33c6c1e8b21a523f971f42b05862bc21614852994b9d2268d6b62126409feefed627d19b7f6a2cc7d3687353b7b4f50e4dac15e56206de995e2025182ef502990f93b1578ac0d656de6b2dcb63835c1273d4b38b322380e347937656109c636473c4c3d71fe9b1a466e2311cb5a8f44c224c9ae12c6a6bff4ae7244acfef93f4ea160f99c29e7ae08c91c51bc150aa1908a12d4a5ac6f0c4bd0c62f164193fabdd8f5b79b949ebe1e8648add39c717baaf687831a48cd7aec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7cdea35642e0c51ae78f698e0d112ade8b5574dcd871a3e26dfc7abeb91e1d61fccd009710309d8bed24cef86d8bdd35e74b96b313a414b63731fdc7f8caeab15c11757305ed023358ce38ea4c0131bb77d60c24b354d24f6a8250d7b69d3128dab38ac114e3bb28c8c133c1faaffa606b57785cc24add5590529ba138748f74209ca04f30036adf441e09e3add1e945140017994f44b81201e1e5012c2437b520f8ebe31328a4f8523afdbcbf5c2e4a1616f7240f37a322236d820dec0ae593bf37e9cb1e28c007dd5d4679b52f544e0c8d0300a56410dc9f297136f8f9ddd424639dc68c7cebcc3ec561ae1a8d1836995d87b2c014d0a9577c6f83ff434f554127e45a81725376edf313c8663165c674fef2fca88cdd820492ff85ccdfc1f6237d3f422e08f81f034c6bbd67b6c5643df07e5abee2f60cd5df07d53e5674ddee7f28f39bcee14e9f7dfa36dec19b33ba55ceebcbfe735a92f7e2bd80ebaa3bee68d0a00eef4e741f3aa33d6e49846db0a1d7eeaebcfaf18de7f77082224ad663e5a3453e4797ba728757eded1b2d03fc623fe9f83ac1a3e9ed1ca1b5c88bf36a861c79b5c75cb12f4dcfe0884fc515350e1c4c5852c649edd10b74fddde102c08243c5ccdfc836962021d3a08b1c81ad24ef06ac3773711b83f7b2f95b99dcf844938a2c0af94dd72938bc751e269729c81fdc07a5d57e797d4291ffed7e37adb1a16cb53ad789c82bbdf8a7694906e9bacad8d864a8cc38742e0a0943577bf309d908ace4c76fc0b335fc9d001a039ab31bae801a30deb42a860f9a999dc0b04653ab88b595d89510c9561c399ddb5a408616c68a17bf1481d008034d39fbad9f8583e8c7d425280d7199060f1bea793f5ea3d924a5a64e421950912e52380c79f4462b1da2512fd3bbc496453d6c2d5eea02ab4602066daa274c490028668d34c64162a3b34aafbe5222be70ede200eab4d88ffd15d2c00cd3f1a3d993d80d4f8465fb05e7d8de4bcbd332740a30e1113dd2a1b6bb3a9e1763ef205d3d5393ad05894b4ac1f90ceb17db740eccce4a613854c63e81391a9ac4cf77e3bdd49643eb5c7d6b5f3fe1c0f8fee39e89e6b87dd098792c542519a3bb02cacba8b7a37384e657dd6ed33c4fec8e2a699868b3e73acc4d63453e548e2d4b0eaa13636266a43e5cb0357a8ca981bf027f475d1cf52827d2fbec1e6fe7239290eb3fbdc02e23dd2f205b571457948c4c985d9bfe2c1bafe192de9f592ab4c47e4aa44e220ef4a985164e3a9e196bc5614acf2463d6c7d3cf99cbe9393ab921fb192d14568282f0303ef60b805819646aa84db916ef875b7df56886a7c756026b80a994250de647d24587817110f46e7b54d79bf43260807df7edebb21867f73296d8511ebd28e7446e5fb5b051f17e903145cfaccde356df3e580828b8a900498690b0c37fcaf314b20f2561b387344151856c913d523f2d65392eb4560a922f01ab4520c7b8a4e26ac7a9e9b70272344ad4da7aaf67c9efe99c784b37a0c899f84f1f558325f37e3180a329c6ff0717fb7e1e488f8fd91fad5aa229d63df7deba57970b6ce057739a83cea7a4b6c41bc11314379b7495b7e6dcc95212ad8917beae64fba5e5ff05065c72a5879dfc1d6606859362d4d6e7392c6aea62b4d502f22baa1a0ba3e572510c38f25780e25079cdbdda32f32479bfe409fe86d2141dce08f939174fcd9ed9739be23a5a5665e4ed3303efa9cf405c11d9073c3b02ac3aa8b01ac11c955408ff6bc2482144d751cded3febb6b302c50f3dc3129e1f48db8d9d86db986d63a77b15a5aa8130c2ec827d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he75c62ff4e2973f41c8d9e5a8483393dec321e6c89ff561d214fa01cbf699e8d659cf8b54f80ad6ee20d574bf551edd5409a0d6b027c39f77bce697626a2e0d3b74e55893712891f38292eebf12a0ef9f15e40ece0814022966f3e70d413dc26aa652f03a744a476c066aef724c07a74ac2b08c9e72bf72ac300937911ac1f999c3f15a30aee3785491c13d042057a70700c34be77318c110b217dc55a50cdf06568cffae6a96a2d923bfc897c07b0e9a911b9bac6bdc3153dd6665122bdec3aad8288dd674a7fae9760699311d590d29574d7070214053eca5a1fc991f72afd91ae5314b4764e710d1cd9a6135a2547e2fbe5207ac7ce058e9516d54d4ec9018dd639594e128c88b8d9cd706e5fb14d640d4537ebef3c9ab77eaa488fa67bf9cb1a17627cf3cb291a71dd5e29e68505d073fe25116af307f0adf6d8ff1141de1ad9d097caa86a5ffb026e6af7fba5ab9e1f84b6f793b1e4120d92177f6466fc5f729c8c609a9c56cb69457c166177069a8cf9dd1c0a6b07a8b7771730508e7d310a1df368747cfacb727c8ef150fd767ccd3ee6b19ccce7d262dcf09487f5508185ec89e83c278fa0afe8918c5fda73c3998d6434a9d3c12e323e5e7941001c4fde85aaf023102a06fb50d746f0c469da4a0003473b7aff5e8b27cbe852d0a660202aac916b7b045e5e8bdf39748f2f172833becc668c07e795edcefea93e065674d556794df4f9a25c80551d9ab495b802b4d33a4cc33387ad084d863399886f782d0fd90caee7750717c7b4a39480ee9cf25426626b69d5a89b7533b054a9d72be7275978e4e5f01dec7630a54e88b0c99f4f16308c02a90b62c54d191e57c9ce14c05115b592d3500b920f74a1b82bfb2f594998f5c6190397b5ed63797ddbcdc221c3e0a99857bbe899f59ccc39f151c78905329125f96a103ade9f095734a00c9efae9e55e57ecbe7e2320503a40a8af7ef07f013a6c4328d0e9215ac0d3dde73c8aa767e559ca31daebda93f9a0b969d1ac7b83f5af68efeff97e14cbe0aa32c53ce4310c7417a37cb37b2d906c07fdd249c2beec8908834fe77a508179fe9949e24229d845838f6382d156cb898ec54e45d12d3ce90e797593e234a4e93cf4ba4fb03aa3dddd5438d605b6ae5f261b16984cad9c695e52b33de2a5d75ff7a33e1027d064ca7bade68466423312b3cc17c8fe1962bd735f90e1ab7f55a8d64136af7ef4a387cee481c007527e6ff8b2566572cd4977b876356a89c2b227f2dbd4aae28462c1467a84352b315da610fdd322e7d5a93e1577187b92f5ee5ae5dbd1a4d4adb1a6d2b51325c2407e359f882c2e1ea467f24e4d2b0f9f332f7a88f8eb1e58608e00c5c2e7abd115e6180ecc2d7a80b74160189baaf4811529c6d56317e983792e2488bc37e11c24251037bf5d3b2f6cb357ebbef595d74a855357da0642c7d9c185eb6942457445ee5e8eb8aa16e101d0456617ebd6e6a18bdf3c17b56acade4e51ba683c2e24744bd7e7b0a4bf515da2ae7e1a6da514acf9a39c9746eaca7a7ff619db6f5344229d24109e967cb0917fa38129c1610896242fe3b96ba9cd0658d8afa3ed3be1e8f3c2f9796407ee94a0f869346c7818d4d10e9dab80005be350e231cec9f72ef052b19a77d44276a339cc23473ad4924fd7e20eda1258dcbbb1eb2c260872b000edb2396bff0e61bc3e4f7cdfb671c1402a9787742c7723088e83b89a3d1fcb1bb6f86eb3edbed65f7cd595660e6fefc07046785c5efe0d1dcb924a364f04a7967bfe4a638cf6d4233d0776e6b1962ee6c8ac7f70aa8f0dad239ac193cb1a13fcb3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h276c661d5e3566e61ee8a34e68f7f5385ce515c7d9c5aca207c85a95f91a296b9e42672ad5568b4e46823333befad2e3b7d8dd9bc7219d51058808ef4a33f30598e9f4bf92fbaaeafad2cab5b13d540a8b314b39910a28f1608e5d5be6827b00a736844f63a7a96eb3617ee46b56f8d46964997fc59a72baa96368cce0d67f2c0c76a8fa2a623f6e19a948bb5ce0f8e7e9913ba94f9a391e4ee6fe57388717b4859576f4050b3eba5643b8a45a6191ba120b1441cb77c94a59d8623fa0ee34d7c3a1a6b9506eb83964010b2b945b40ef8d88634ec1adf56c0c41c571147dcc05eb20037f4ea551fdaf6504c4b183d65c05275ab131d06c5f2ac743c59cdd04da53d8f173629f8284df34edfd230d476e8b0fab9849972cabd7b23fc27db6c75863dfe9c520150f98c7004ecf9b8f2a05f8c8c7f624dd48017ef3c3184c55d5a2fdeb32b3264915c03f24ac01c0fa82ad88602e8e10a158eca6810834be64128616d8d02ade163509ce8bc8295e0a1e3043ed2f8f0b38a6c8308e4482d7f280c037e490a5ff5131c612dbbf28d657e989f3050666ecfa67450be32380b6967288cdcb0a3e4d84b55e739f2508b98454afed2861f1c34a2dded663c35d65cdd7b641b9ccec3417841924557e44914bfd3991941fd6810db1cdb64c2f9326e36b7623c8df807b89368159e72167a360c93d4e06cb7cd825e36a077ababe3602f3324504dda2fb9b7dfb313fbfa208088246675a35a3fcf30ccb8d7ad2776bfa087fb7a590a97e1102b3cf446080ef66d86b797890bbb481671e5b0def88d6d428a1bf10753883c6144aa7d1a229782bd3051a573f03c19e669a03411a175aed25913e8c3f9bdd7d1cd125596d5eacc6af68f63622ed2e996df28cabb1503e11e8390d0fb36eb650b810ddccaf9ed81542a573b1b7c0bc7ac863351a5d4ba2fe18c68122709e1695c87a287fb9dbbf4010acd3791be613c8201c2cf3b4c98e21c7107fb345d63a2fa8093165b31edc06d295301a2459d0ffbb0e5ab595d466c853d713c341d40cf306f8116733ef52c1092fca9d23b6b02b9aacc61b8642d8af2b5b6a37bff51bfd66c979f01e61c356f9cf8943f480759b750a9cd27e971662298f9a8ff64d5805430493d349cf97fc1da6c6f9d9ba01a995cb0dbeaf5fc30b9edc4a475c939a5446127511308aec17882e0febd06f177294403fcfb6b11b90061ce0cab522623b0445acab38c5f52d3783cfa166bc346a52980f3a448459760f645f12b835bba42c0a531344dd1153951a3a1759eb861b6e6b273097655cdee61c922cd48c50645514ac97ce3d1e9a091bf3bf30d8c17d71ec8ab6c929360a3e2fa57a559b2d92b870da580556191582bd2982f6a9657095a9ddc1efe372eccab1770453f70881cefe5fcce25706fd0be24dc9ef439b3b7e21de31a7bc0258ff528e5d70e9d6d5a8e526bee186a0ad0966ac169406d9766c2913a4f2871977edeea3e22a7d12ec83a814cf1575439026b1bcb581c9604aef687e4c0a3f76c0a3a9e78cff0333d6fad7a2ab531564c2cbcfe5bebacd6eff6cd91fca8a8ea9595da6127b1f0f70e4ccf5fd7c7fa98e4aab08f513b8800f2bcf90eb32b88b81bbf0a0143c3e9be27d36f9cdb0a456447fcc75b1467ee12053765412bd034018f31a0f70e0a7e55b0252a1a1fb877c6cb2292d3ac62554998837ba83ac4d858e43acd4b3e8c447fa72d785242c4718b115b06a10eee54bf495339be3d196ba8a292d0f4f0be38778534f5a853b94d308033d283170e814b76336d138d557a70aba9af34b986cd9cd54cbd467003e1eadda417;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbb775eb20d37db6a4982935d4f6173fdfc83a07ec1f410928fd320e67fb11ed7216c8487e59a695b69c2b5c59e4ca97897705f33ee09e3b4edab3121a38fcb0ecf45dd5cfc0a265dd14beecfb41776b7a9f7a458f4233c21008361fcb37414c27862dfff7578725243aee6f35edf861a5a4b04e2f8127aaea05be76e5566ecfae94b33429484bc1a1794c8acacbf19c4d6a854be3dac07cb0be420d43ab11a8354e3757b5588ee93ecadee4cfedde59da87e3dd0de1fa2d7e9e6cf00a2594908a6ab0b04f509bcff60d77108675401e80abc7c1fc01b925aca47fed763e7d627799acffd53576b97c4708e9297a72c643d1109d14ba4ea68ac4dd0970f62dc456bc442a146b3df4db1ce0d5c84f74a7d3b1be82d465b1605623b275b36c8fd3fe603f952c0ec195b9bf9c2948a29ef4c8b1dc17e1a30ba056fd694feb689fe48a1c27750163e51176fadfe099760ce210bba9db28cb118bfa908e7ec73e01aa7a390144fb46f0728fc84f1fb697f6519788aad9ba9c1f9fac8c02e7c293d666a004a0e8e6385975385907e4d21eccdf7171df0eb8946505ba0b5d2851f3c72f55eec6934aab8574c6ac0930016efd988b6c2cbf9795e2e04c649a6ff121af38e4303183e900055734fb711dffaebe51e206001662319bbbc6face97d3be5f5f7dbfecdc8910d604a03f153b2abcc22ed6e9af4552427279c8504c0832d8638c1dffb9dc8d0cd3d3f9f5011eb5afeda1bd419d6f998e702d750be8194ea8dc495dd3d905c3e255d31fbebfcb712cbf8bd9771af28efe8b7daf7140a8fe99e6453bc322002c49cda728be779e48deaa6e1248b6c9a09ef56deebe5513480fb946ebcd9565b3a856a5c201ede6c2aef1502ba3e6c6e257058f43db897aa2976569379e937e34a3f1a0016e4add9ac7e5a8abdcaef3e3031ab272fe93c3c40d11a11b3ccba7313d64dfbd63da32500a56f2ec0333e2117f28b243f9e8ac0c3ec78937504ce7249a9bd4a29dfddbf144765b95522d21dd042a85d2a921021f3baf5dca4bf77a02357ef32aa4d23f8f8de34296b39064ef6c41e7ffd6c44ca26ea6cb48cd3acd5e4a760c46d053520319327368f6f6a9ecadf54b2256f29d2b983188bdcde122f97b4fdd893d0a2fc06c1f76573fe80e3093e3c2ac7e8333cfb8739cb2fbc5bab88ec3ce537b4fb3287aa624e87b8f245b99697240d8e8589bc5e7ca082b94e49011fc1cf074f7fef07c43f2b13cd7eed8bbfddd8c77391a431e593a72587de22257c354714831742794ec61fd64e740753aa9ef5e40d5a63d2be8502a44b12426c9e4f5d69b3caaf44b826aa2bd6d09bc01b8eca2e55749df6b261dc4646574dd0c4e1d773623b2f285c5eea712c65f96eca4bc09397d1aa05dadd841e63d65026371133624de3aa55e7464bdc78b456155bab5de93666fe219b11a8eabbc1818424875007f1014f88c21e8d677d5ba8c9476f84b3a826e1daa4e9b9927311ef612a90f5f7b6d0e6be945f28e630217500cbd3149383081b0cd2cf284350f2f7a2b05fb583e3299c051c6cfab8ba115639f65f8dea1fd07eb582a6af6a1d07536038d69d5f74693471a602d93970287f8cc7917d8c2a9a1512f8d91ad026303b0c7e7c01e41cffa44a27f8c245b57e4d0f065ea5761fa8967bf32be8fa941430146747c337dea2c14e88736e96b7ef0973b30f440c17a6976bfc920994b78a3b89dc37656cbd4eba896aa812bf41b002765207f0a0777a0392ea538075158470d6911044c061ebcad5fcbece441b2243753a95e8eccfb5d31dd783b6f86ddd1ecceae58a9ebfb2484c564d99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7871d06b5c452d81aca16dbabf84a56becb7c1ea4159ebba90a1be794130609d38daa17ac493bc82c0237f6e374ce98c8b9df84cfb87c8b7c464e329e267d10457908094c4bad1783e8f978a6af776f33dcad23638b9b203ec2218bf54e6129ff395686e682ef85c2c0e6ed0321160dea00ed807397193a02f060aa95fdedf9c909f3e8908a6f6d3f196838fc6f048291337a72450c9c00882c6bb7d7401f5d1a82cbc3831464822180d4f1f41b3061058a2cdcc1f48443d404a1f36ac3f6ec992c87c28fcbf8d176b7aa391004f5ef558388a148cddd1a300db96f9fd944a53e6a65944170f651b0e6ea4025b691e404b65292bf3b9ff3fefec122039f17a5fdb5ecfe9e72b21afc6851703030342a2091480878a62fba190d6846254fec70bc4d7320416be3b31b1680cd6df61511bee52cb5e2cef6cfb65e9e066f54fb5c581a114c75c83c829f2ad750b1d8e3bdb3a6620362ce70d72d4211ed2b4f43746de116f59b6c78148185e73dd65a69691fd49943da09d0b69240938e37fbc5a65ee8548d68ce69b87fd7e98b35a85270b4659d950b245644731a94ce23ed7d119d6b58b606d0ee1eae951c48257397d42760feed12c00ac8e91c4ac236033712ca04906b06a59343ee9be4f6568c7bea118612b461510905b3918ff0406936ef0998a437ce8b424c648e462624835ef9ca98e449c449b2730af5ee2659a9948085966538e08d5b3613448380f15abb1327aa679d71c94b5f2891f0f363bf5d06af5dd624fbbb2c3a3aebcc9027d0b1edcd5ed9072f00314ec89ea6f9a2bd7441833f16541a4805f311e0b45a51e4519a24175a78a5c154b6fb5bfdd1adfb1b34fddc44d42a98d48eef688ce969b240bdfb179d699a5889a03a29a12b6623ff53472f1e541fd8171afacf277487867ae1e5dff9906f7882d4f736b2379db5dda6e355214b52247145a88bbb192c9e625ceb23c47e824cca8b4be94919183336972e25c056c45fb682cae0af2323550fa6707b5770643388ed1970160fa6cac6293aa2e3f7dcdb00da8c026d6baed2693050f7b30506c9fcfc1d37efd9f16a4ee2f0885289d490353949719e82eeabad4f9eb13763c0dee68e5b526a4b3a88c064e21c4d0360e83145160873526c0b529727d49e51bf71ddaad0550371e5a9814c73456df493670fd58b4a064e7f9d4bbddd3dd95534a54b00276022485b8ce0f530bee66e130f32d781a5d3dbcab3ef4b638d0b8a9a0e08c079eac37af0491a40791432f49a6a47699cae1df3d1979d232c6bfdf106571939c0d7abd496ff7823ac06f67458a8affb1080de9926db15baa5a84ce230c4a2254d1e6c41465e4ba14e1b96c6c1cd174de0588d746b071f54ccc4adadcc684942341b111f1fda0c815850d9a867f35acb8621f5879c703f67827393096694ef5dba31d86317e72afa50e9f422d20231aba8a7c5afb76ec2160215997f6bf83392dbd7563af9f4d8e29ad794e101011adfd571d404787d578783c19ccc775cdce9de6a45471326411c3fb01dd66343d5c7c9107bbe541f25a31218792147b6978d127f0273023cac12db84093d7870b74009d6ab4219b7fb04bf30984d547f5c2026ed11c240e005cf46264dd0f84567fb5ca09dd38a5cc420ce682c678f34a26fe57b474c803f2abae7d04bc89748789c6ec1a0a3823508a53884eba81ae284153025e9c7168079b807d71979e0f3efd6651972e20e68b8af499bf414cd31ae7630168171cf987b3a10471d245a6f1773d06de2169b2ab479d78fddc8f8f35d1dd590411a6fdb345026be64b2f4fc3a7b9101e4090506ef04c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h23df2be8a32002438a6c5aacb73c4e80ee502ab4a421b9b7da889d3fca0c8952a59e07f7e6c914047a250eaff2479501f97e89a012bed6731c361ed3b3af03c060cbbe7a05f619d07ab9996c9f93579f37af7d95b044461bbf5fcf106dc71dc013d04c99104c1cdd98c84e638139f26fbec48a02981f6be2a96c765125fbf7fed2e04abe792d87e9adac10b82165cf038730c210c5bc8d360a2eeb55c44d155cc2ab6c4485297802da5779f570718c88d2a808dd863099b1b066f293b5d7d01a62e218d7fab86d4ab7850def588a8552f65a09815e121abc5da3fcddd5532a6d65d11c35e9089ee25dbc9504a027877e656a791070344d92323e46888bbbc5311174c5a7c7bd215a888f5bcaf154ee219fc6eee42fbf3e0de3e73b7fd1610d88de4c567e8a086e2d56dcf95345d99ce851a0aa5cdbaa375a8726d3a6cefde5ed0598284c04ebe570e451b4ddeb7168a6dd9adbabd87eec81083dd0e6e0affdd12934a52eb94d1d78a330525738c7c763af9b29e9ee157c62d4a85ce8305f49a2410f29c95ba0e3b09bdb2d544a774ec205a1822875ec86e8d8fe79591954ba56f72df7f2df1de659e7364268320583c3d4a78e93401fdde5e6c4acc02c3a4a2a11a4577c11db5f78ddb5db6857a094339febc180613691b45c73fbc73137123288566e982b2f2e8fd05018151125ba85439d1d5e1e00f14e189a7f650bbc5c3e148327b23281a0de58417486c7a651aa4c2775abb1d2b1771a460f9c77c70d1566899a0bd6a78ac6dd19bae5b2555aeb3e25e76993303eb5c6fbdb73e87f3998eed3e2d9e599ef0e9a45fc84953c4ed055f0546f41fbe215fc07d7ea1af908ecd85db57d0bb2eddd519e0f70664a695e7d3aacea78452ff6ac29d191143856b5397b7c47cc35ab459ca59355f0e3e59567e9e43f87fef250903893a7d0bdeb0c5aa9e503dbf6b339bc4356aa8cd98f21b13f8465dee6bd5a8915875e4be2f5b45eb01ad087c6f3a4f88e371a5a45cc63e22e2f4d63187fb96a93d3074a06dd659262a3e9eb57308740242f08bbb6e2d6bb5e47d6a6115636845f1c53fa72181615b41bb19a58d888ff5a9ac1003c36d64e94edb00e4c6d77c94ee0a8fcbd2fa2cd39a72e99fe955e7a1591d3efec8266c100939cbaa40f30978a941d944aa70dcdc0dbbdd8a76507de054fed4784a62d9c93e91137bedb8060ef30087e08321ee4f1adf25b4114e8b93d050569cb570d786bd8c563c53b2663c7a2ccadddab6bc3abbddccaa89e4ae4ad33904adbcfe9429765f805ae68f8c16278ab99b510945474c0abc5e6f645948cc0baf9b0189c08e675627160d693c905da5511219863931875e9c4358740100d40a37ce4c2d378369ee2d7699fb50649282302b7f29addedc5fe686e1091a91e7865bb2a0ac2b5aadeca5699761641ec101dfca3fe5432c69e97023a94b87ee63448fc719152ddac3c27ce1dda2557bc4f72e2d9d3fa37ad3c2fb2ba1c3912ec323461c6576f4bb3b83a474ee9cdc9bc62b0d52167ced4a595a7f4f2854b8b34e0002ac8a27cb33f92355078b7e8d1a46b0e3ee57807f681cf5fd2ed59858ef9ac7272c70d9d217a9612091567a1df152477993dfb019e66a25f65a6c5c4e8212691a2d67920571b8337c91f5a34549d65a8c5cd2a73d4daae2dbf23030c6398692eb343b311d43657cf04eb7976f10e22418d481902a3fd1b960699b6e9086f0a3a103f0df81538d4d63050edad678810dff87d388ed7de19a6d2ca9257bf19ce1c9a309a68f3e4d5a9e8e2cd98e4d63d90e88101d21c00a6a195add3e6af939295f513fd03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2d143e73a0b12f3af9715fc1404fbcdd23ab4bd22e457e39e4e8f4331d7bfdaad07acb326f55d284c5ee3de475ebaf5aa5a5aa4031d0ad932dd1bb261a8fb297b0ec478451f352518e597c1ee29a9995625bf707dcd2ac9b02c3ff7244acdb777d7b7ce24da7ccb2c054ae8c4e658b92eee881962e4625270d8f6fe6492395655b7b7574d0fecd8ff6c2baf2fe0ee49271f6d4d9de39c438f0ae833db7767e438c7d07c1fd70fa2eaed902518d55bfcb2d84e22d518bebc3c7f534818b12b5bb1238c37acc5931c4f7cb9b07957f1cf98f523fd444725dafc53c007c1e704f197a43b3a1118412c5991294418da9452d6d1de3d7edd2c30f4cf3c0b73551d8640c48957a1c05ec5eeae1dc066c23ee4eb5ddfdb59eee67cc6909b29449e6b7c27b40fd525fa23ae8f56406cba463a786aa82e48653a2bf53cd15aedfeb582fd88317dd74d38c06b78a4212629d72e42a824bd92870ae9eaf7277e10da103612d540ff4a17dda22d8c27fa0e50d592d9082f01230c96cf7d92577f469871ea79c9b3e651118fd8bbf03f16f490b8983956fab239e88a1139bc32ad1c5d21d86c306054663a5e1882608c94ec8587aa7c61287e217ce2867ba1c934fe6f500a43a2f8c5a16eeb712b8d940fe84e482257c399ec6b4d556c396d2054e00d8191b9c7b1b127f88f7842491106ea41afb03fdaa43a0cfb96ab68b67e593b9ec683e69f547633e9b63a9b80d2a9be5963a47a8f2a13c520aad70d32c1dabc7eac852c10e29233322bdea4e294bdb97d70b1bc30be7c81eb425e9f4b18a61937d8973ad665808f1fed76d03ff4041410ba128975ece2c1b86ea57644e875a1b5b15917d5e41a8f2dd7ee182b5a3fb56a46c89bcb1f50dbf64ecdfc7859700e9c29ce60dbbb1e18f78a2f4950ecee839338291d090c9c92599bdbb886f08db1ba8885b4f5270800afda2f5fcc9344246b16dff8dd2a934a457f59660f1a40905d787ab2bb6f8576b95d1f2322b32524b39fd8523e41f9bfab5740cb95a5a09690ad1dc5a70c32a9464ec97ceedf4ea54d94e45ef93855fb7a5fed529922752b672fb4b61678764c975ffd39ac267723f8497cb28f9bfea13aa7970b3d620d6234cdd9ff9b846a40955d899b83138df90e025305df40249c8cf41feda99f99da732dd2a267965de40206ccbdf098a6a7ced9add72fd5be4161394fe96ff211e432ef952678f830233b996f4be7af71dd43b1f108d0f9ccf96c17637901bb0873bb7a80f0d89f09531ae1f3a293af800f48711caef5052bbed5c205e99e7784b9c7fc3f54ed7ef16795d17d4c5ce57851f5a61dc603605c3ec6f83d5adc0a00c8f05aadff3d0a03baff693e1ec49acd8c63e9d8b9829b42a773c9afc3ba264247063bd4f815440c2a49c5ed63c709ff69bdbde9091e79e2cd229e18685c594dce7182bcd10ef229ce6d43131c833c8518b37ea3d89d3fdb22c7a99a9cf345d8b7d5d412fae155bd940c759ed1fb2e108459a160141c5d10b92f3eec8b908f393532070074c9f22e5ead789d4b77b13f10ce03e179c86b2d14057ace416d39fde6d033029b4c9fb21c40f6a76b70488622c7f12e808596637b43d920a96096ba2e71608254e6f58bb3c8b4d4d739359263b6e554ac843692136aba0109a77a6d712104c3674c9640f000b8a5c810b5e932e5743f35ca8fdce24933c0d564188dfd6c20e56e1947233d70642a09a55ff402055e264f9e147510dd0bc945a5bb0361f4e393177358b943bbefe37633db1f529a215c40848e694cb388512fdba7fa226321c2666ff50f231f3449f4053a2620a863e65f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc265505e5d41aff8e4a26a0f923c6477ef41ab9658bd1d8e5a5004da5a8051d16a2ead5c5de35766a15855a2a95b72bdd1fb25b93b4073ce1133e7f2810768a653b6100f0cb138ca7b4ba2b7d4743ef0e01ee2ff2542098be82e8549c5776d2c0a11f1921ca88cb8fa80ed8ecfbf379f6c51ca483f64a6e23bc8f8bc627e00100c174d5dadcd7a7e516f5d53e1132ec775a4f93d573ee77e05f8d2ebb7af7c08f0a8140b214deb9a8a13d08d5c30dbc32c086f5ef82a3aabc9070d1728aa36414c0dee227ed564209262bda704f3b9442745aca76d852f4650b0aab66df7f4af1527a0a138be19af4ede65863b36d4a88d2e3db2b0b3dbcc27494973fa5a348915251b35f0615f99d0e49f927ffb0e37937bc3bb36a13acc2ea57cdd78e3632f3bbd353726074841cfe4a9272e37e4c8a4f47c307c02d7eba3eaea77e243cc65d532670b8ade09ab667421837e22c602ad969e278997dbe023502458b02aed5a6fb3da6163a89544dab0260ad6495af9ddc57d06233c263a763a950a8e1f71e94e4e98203f094340bff3dad870bf70f549bba56914a78c5ef842e88c39765be519eae65e8455d2d379a0e89cf44efa68f20d48943b04638a3d4c6853291669cfedb3ad1eccfea9d22246fde5907535752115fb385d9d2db020942c36effdb733290ef4e7495afd3b4b371ee652473d284fe67c602cf58097e98dcf3b06e4a3ffc008dc70a2e82fc50f6a8e22227e841605fde8ae36c951802c9d9a8e00f518f95a620d40e3b39a54a7d3c7e7daff515758c21afdbc569ae2d25a4bd47045003183320dbfe8c277060032c52cd697d5fa6aa7acd303b3ccb7cb5fd6b80ccd684e36c71dc964582557a410f9df0e0e8b5634455b9f77129f0b204f0026a87799dc2b84a29adc53b1dd112126658e786f76bfd9c5e5f42dacfcb0f4dd17bfc8c989a7bfa92ef826c757f36331e3153288273329123bbfe5cab10bdcea1b06e8f4a7c4b3248b7e1f98e6b36f604ff07d18afb752be8b2ce7fe234e2c4e92e7b22abff91c7ef6c1f1226f8fa651bea9a7da9b4b2f981759b3e7b43a1494f822c9b4ea355bef25374358c49447410eaba1408ca5901bbe087cc13c08ca6c5d2a11996f7b963854cbee00357d30f7e83cc10e365961a29400bfdeba79b765e79fbe51ed6f8394d9114dea02f8824c5dd8f873d22c1e98fa0db5bc09751e9dea9cd64d56ec6df9483fdff6c5fb8da862b118234b16b5a4fca67d5021690e79413520c6ddbeafd22eba9d727e403babea9ecadf2a502637e8f5ee0be3575f9690493d2a77f02835a070a18ad7403d46754e94fadcaf27a1eed98f127580d9c8d46a7f76d9c263678c738b6af00dad32044a57ffe6b7e6e6d206fdd649e81e265b949204c235c30f3f6d6a60cc6c9b5aeb71e25f29e23e537ecebfc6b4f6786ef51e4c10c4427e996322abcc4a4037e51e271d954b830ca243f0c2600b679539f056bfb45af42ecc351f32d0003dda2208b09ed87cdd56cd7c8af907adbb399a1e8370ced675bb03426c29cd4ce411b6e702aff99d76e13c05939c18bf41eb74dc96d7eea788a15d031a67818f04a8baeef46477634e5d665c776114766b6319e8a340f3b88da512e16ae853d32ebd99aba8e37556d8469ad23bbae90a3db0b94abb2822df40aeea7c97cf6c01218d859b8275799c43675bee1f077e2933b1281acea4d34dbbf5fd657939fcd93668f76fe6f541633f8385ec7c7702010422b7130ef241e5313058c28d52587288a23b3061234c714c9ee2c59cb3445bf1dad56024a0c3308f09d3e8f2d21f138db1a9e38efcb5f7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h356720036ca4decbd821c6d0ffeea4a37122d5b64d858ae47f732bd181c8e99c5f948b35044d6935f984f8b49c5b8f69a6b66a805ca2c485d6f7a39c2fe7ea507c2d7ef8950387f4433370cd9f25cc671efc2bb28983ac2c131f42897807defece621bafcb9ab2efd001302cee2cee728f061dfe02e2a54aeca86d2f709b45d45e414d6143236bbdb9256991657defef52514167f0dbaa212a33cf1e1f8e6d498c8e506525981dc096593ca6956b67175a9f0da75619d8ae57d55e4e6940959939492287b641852ea2aec278f76a83f3f068e21c57159cf9e1973e11c1dc850239fab466581f754baac5f87994762960de5e63b5eaf4b3cca2fad713d810da386338c5a0e905f67c643a1117c303845179e36dd92b3826662d568dc44a0510bb3100958b2b3b0ccbff00aa2c234ed8ac68bb1d230e12d1fc307e9204fdb87e8cad7e2e05ad3a1ecc76e69b5f4fa2e1c43b61d44aec1c49cb94f40a8477e0048a5d82045eacc2e65bf308b27f61ed1103f94ee7cad228d4d3f414d6605ee8d2fd460b312dc7ea08c21e4b05faa391de7362fb9223f087b68a0735f4809aeeef6542124b4b8424768d6dd21c89880511c48394bf6741de95af632f519c98da0b5715f36f7d2fcd2179dee5e00a88d535065cf1ac46ebbbdece22cbe5709622266ab74e785b6f09a0ad4bcf6f5954531460b07ed03aee94f734aeab01841e161d204bd8c289b4d5099b02677fa96de1f21f34b337b22b71587abbc1426890a7a86f2d52cabbe639260f4eb069fa994c2a05305d8b5b05b890eefb80938cacb97efda281ae1b2959ed760fe225b567cc413e400e0fed49280244f8fe4bbff69c4591c62df809e23671f919c5644996d9729d54f3fee0b951e94c32890390e0c60f4b7b49a239bdcc5ffb51f6db209f36cef82e4151e249b49fda26a595d531f5b61e79049dacf7c5d7631bb25b8f583aa1d01411d183c37c5f6fa684a60dc75f2fbf05c6525b532b09dc03e07458766f3e8313e65d108adeb2325869e111c00dfb656479832b35642cd5d6fab108b3a15c7aa459fb6b48723422698596ad90fec779de15134f2d1282917a3768cc0c00eb3918654b844005d39d4a574cddfb4231ec035d0df275a23a7a62d77dcb21742f243a0c4ba0edecdf4097910085eae4f857ae92bbd6f0b424d20fa87970a17472df7fd142973803ed186b279f7feefc160d36b86d8d78bdd269c0b9c98e22b1e3c3cd0186c35594c12002f9f79087c90bc610d78a08ae6d3036b9dfa22895f1026bc27381e39c4fb1b0873803f5ba31ec13085782d8180e58d238a770151f5789ac909f688b7d69042b4e93a818689860f09608b19c813c4bb999310550b3fa34d10e1947762a8bb3e33aed34ced9154f5f2407fabc04996ff4daa2a2811816d05d98045d18a707e68474def9bf356e51dcdab3dbb6af6cf32204045457c220198b609c011622e256947dd7fe69b0a75fc97e9e4a5d59a017508e27777e4ad2e5618a10c21a9b5c55abd6862f7176dcf43ad16227fda6d92086b82a45551f84151380f7ada5e1e5fae2d514f5f48b067547724c43592cd6a0926a564bd6d6d11265a533e2f14107646fcdb564f899e6b71bf02694f2fc49f2c4470ec296377c56620481e16187eab66021e6ef6c8bc70ed2f19d5a3e25f1efcd280e39cae3b5ea6a2dfdfd6fe91b07da5eff890edada3f1de82e263bcffffdc1ce7ce679a3942659ea3c5d380e989e56f3181525ca780e03cb84c3359eae88b8fbb36ea1a53db4f795fe648457e524b5c87a1fdef1138bc5269601a96b0973f7cc39d042e5f4bb22;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8ac09b7678b3bb6e163486ef4bb1f7056980c68c774c735d015b28646f476a9ef2dd4294cc082d4f7ca921c701a8f1b7a6d79a9bbc6185526c7ff9b82e3eb709cf1bd451e047440e116f64e627fe5e5ea8fcbf307ccc305e4f8fbf7ffd35972535cdc4b6310aea673c3bfc35e96ccafe4c962ddbe191f1ac360e9c53cb129a9963785a9fbad01d29daccbda5d9f215f660167f9a4767440a568d3103aa42b20073e577162c9f2674d1d0d8469fbaf1101ab12dcf2b31e0748461c0f0986366f71b3d41b247ebcb5a9dc73deb7426723eca7774b84535a1ad58224cd2a033a27a20d4ee2025ac3b46be19aaa0d8e8df142ffb07145296bc5ba9b612db0f9d30da2d385f8341a139dbe5692e68a59be67ccf31caca4cac7272b83d6ab7aee12e78fec23ed11fc46d6e14de90ac476addac6498fc59ae2e0d6ed9a2d417fc780420ee4b2c010c8c675655cb94cd033b086da278809b4536de920b0eebf18f31d253c607327f32f504b5400f99a57515f287e0e16b07636ac9d14de0e6b5905082b6be881d21d093c251039bb1a279e9d90fa37d5b2c415aca47ae7352d105786f375e96effc72498f5baaec3d377dd49a6521378f4d857dbf30dce7959f311070dd2f4bc795f44cd15d564103441a3e85b82408b869bc17d33470f1a9df759ce9c29ce70a185708d60d0a681d5e561b4c05c542fe779c9fe2d2f19e1f5b9a7106bec102f42c415d8b6043019bf61f5ff4779d9c76bdecf2025cd9e6208c6ee9f16eb68ef883fc3ed1af6731150c7425b5742485719dbdae7d84ac0532a37c2dfce6ae5ff68b2b46fc59380e18e609b85af2f08ca76906f43da6ab01a07e6be9481f46b9478710793ac803f9a4b1fb7d7401bbba0eac081bba3a5a719bf35aad254aa4f27a9480bc02065996b5f0e75e983620a7d2b10cf9d414a075ced6b9342bb93f732cb4979036a4c756a96e554580802388ba84df8301ae2f253e9c94cf22657ea06eea06f92101cfdfd18518fe811b1f2085acba173a37dbf96052dca9a21b461594ec6333c4e5d5fd189bb78066760e123ca2b7c105e35bd77b37d8f1eca3702bb641ab520a448cc7a196a1e990d29fc147e62e642350aa8b64680790bf14f8f9e1edb77f34e6c8f971ea89c0c91690d6278ae6cdfa8ad8f1f309a0ef10392770ef4853cf62f5b7dcf32e6c7288fa3674ed0d10ec785a7b470044690030de5e85afaa8be269c7263a9fdc5c49d2b63a98fd398c35b9013c2daf0e3cfa232dce2f2cce151567f7db1b0d5558db80767761c733b28bf55c9cdde543dc267a48d03bf040a0a29266450f20b8c0da5fd958cf387225e1264a9d6470df02e6446c999fd63b28187440b409c4aee080ca573b89b23f1859409505a670859f35a8813d7ac4a21f57ccfe9131d81d56c309cdf34ce49fda426382aeae2fd347622a90c3d042f5d1d72c2a6c1dd6119d8ff6d8404283011734a3c314bc9dbaa9b93a321736bd254fad1a387b3c9c635930ad19aa7e1dd40666106788ebe279709642f79cb4b9e7a66638ddc998dea3af835c22a64d2ac0323aa28a13feef365ef8fd0f460edf8ad1da3b0c14bded01f514a87177b6157845aae1d1ee937aaacfc8e99145aa299011ec33082fd0cde28c38d268e6414096c2e0f011c2dd8c786b386e41cef4e278985d04ba2535cd191d6010350eebe77f54c61cff25f430b60f3d14ba70a8fa543ccb845291eeb1fe536cb1de1ea44e846f5dadb9f502b87e8bf6f53a437c81db22c1e61278595d5089ee41d1b038c490f13d28ed63f38d001b6f413f6b263ee1b502191c00f7dabf2d3905b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc12ba72770e6a145b4720e129ff9a7c78db64e8441b9935025baf095095b5083925227541f25b0920731ef1bcbd377a29b14e9429fbf24524d6c7c6d09e392996895e61526974aa334016620975e7a8bad04269d10a743e21e58f72a987d9e29a195f85d435531a77b2248bfd35f4449e41880cbbcde172cba809f411d5ac6725650eb89f77cd065deed87944920a6c2dd526e0166d2bd5561495a2713b40d8890345573500223d0e7c9de891fc89ef7a673c395f7f3e1dc0a428cc5b2d8ba4a0b33e3dcc7aa23b16d8432918a76d1f4a0d058d84b3a691ffd0f7cfabae163ddca4730ba7a380a4e9dc95111f8ec890100a92c5117189933bbabc15142925ced00c5f797f9d332ed8837d1e663029be01e396807ffddaf49630e98244f9c0f27d237ea6b26053445bb0b0b6bf1506a403cc53990fe5cfb595c2b17f10af99446b7070fe6b55226e6a48a8a3ac918ed3a2b3550af097dc08adc56d7d7063eec16ebfea02f951a00222cdf3fc7707f7244731dce0e8656f95f29a9e29af31b3e46edd4772b3bdf752f6c2b943cb643a42e4e813a4511aad4116a2bd3dd20c2d01bf1c4bf195e822a82f6c7f8864eb30fad0197efaa124727bf293efa95a8cad5b33fc645e267af978ca42973a52992d961c328a0a9787ae2e6fb1d2f5cce71927bbf7af0c6a9e8f6cda2dfb1405929f04691b085597e8f7a06fbac756a14012c96514ddc684cc1046bf508ebd25fec083fdffb0afba6c9afbc4b019a92b68e11facaa728d49fbad7081563540a18fd217047fae12581e0f6590598d25e829cca51479b3dc2042e064d934c629b6dcb53c7c63b835d4c63bb2c2d9e5f372aa12992919991dfaf58e2308ca6f6f37d8454248cc656b0781f313ebc955ec9cd689da860f98630292666b66fec06ca82261fa3b79cf6e0358b62f6badb3ebcf676d97852d7c52d95e14ac8e350a72b48eb3d15f250af4fbb3b5e83399c42580736b0c77d2167d4871df0be2f5b4867356505965a27c6b0dce06f95b4adb023a51ceb1b311f0d7c5e1a023568365b11a45d2e67f875ee3fb70f188495e3a7d71145d2a29f9697ca2a1610485ae0a5a7a60c791e3e82cb605dc00390c0ebb755698101f46bb580862d6c6c88f5cad91ad68224a1abf8419120adcbe1d1e854551c09cfa0033d2d669cdca7ad6c2b211a9d1d1e5139be3083ed86b43cd4f8f117e823d8e0caf5e554e7e5ec2f138ea6b8a92826abd81d74ac831eacd589a1316747d7c4588b6769fe46c9bcb184200a327ac8b6968ff8807dca1de7a79827dd21e2d1f4ed3959171856d980fda9c09ce3d07c1132afed5ae7eb7b7ebb31232347127baf026d6f747b8506dad76a66330ddc2039be1a332da163f3bb031a6eb43f77b2ecba0fac77eb3f88e9b3157c5eb984e2cd5f01795e23a1299bd99c67b97612373d100b6cd44a4da780b1c63236e43b0a357dea8d5316e4a68b6ef156f92a81b8825223cd7620e95173d7a873130d36c683a132cc63458e90e84caf46ff15877dfbc91716fcc1727c87a0f91e7f1654c4117afc755c22e3bb19932141045d53de5bd0ec0222936421d17693e126d98ac9526953324ea9bddf260254d564d2afe0124c2cefa91e914e7dd1e0eafdb668360209c9cfa2bf90c4869c9c25893edcee462315ced1c26160610bf0a37406f4a5b04d9fa280fc2eff0731c0c2703137bf0201b10a55e5828f04cfadd6678825e0619f571c40d78c4b7451b41903fcab711360926eb942ee4ae886d9a20627abf0c14c2bed8e35d3678dd27d7e4b6348052e96731fa6bb856ec565492e2d1c091a1cfb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4709384ee2cae87dea0681e4ac8ae216d78ae6b6f6e275c678b41f2c95b37065ff1e38d22eb5f0ce0541eb07f3c6c4a19cec4b517f4309572b35dbcdf113cba66e96a1d682ad90b5a51bb66d6d088ac93e7b1b36d62313fcca954d5481e60b6c8695b5c72181e2756cf522f802456397421966c970dcbf6b38684ac15bb6a21db89bd67b26202a14d52b3a7accee2640481f68314d9a673beb6b1514c364cdbb53b0d7c500db8dd5d039cfcceab0cc14ec7e4f8b88000dcd8aa3e0200d8bb197dd89fe1e1a26001c0fa7e04c10e5f35abb8e59fb8632e3d9081f8aefa897573075a1134395c2fe0ec2ae9d52b78603c2dddde2dd4bf4d75f3dc92b1c40db6785b3b65b1cf82110a8b8a6b73ab93d9706fbb951ddfbcbde0ca12b64a4b2ec19128d0f9c14d5df5def627c0ae3183ad02970c0020fcf80fcb7d02b3740d2797d6cc1293c6fcd9f4f0f6bdddac3d2d947ab9a962080c5343583022a5dc98986fca9ef96c549f539ea84fa85ee1ab673dc494f9156b61b23c1027a3be210fc3c386f0b9a455a4a320cb90d8d828c1d276daa6cf331fa2eb77effe1db52643242530cb04c9484a77140b24bac24ded30cc9979bfcf5c18965730ee66428e10ee304ba7a03152fe68d4ebfb0962604d7f2fe43bf08ab29b61f4fefaf597180c30369f0e73f0a9597bfefeba2eb0e539eb9ec10430828ed4a76900bafc3db856bd1244b0656dcd99e44b67966514d691d99c1b6aaa7dabab939185984e622b2d49442adba63fb6a1fe5b11318052306e3ae0b56be34eb8f515b637c89c1fe67b33aaa738128fed498d340d8f5553eee43d4c348b57a984539ae4db5a3236b46d21c2cbb7e518786e29fb54cf65d6cfe2b89fb79574ecebc46865bc5e16e6ebba4d7492b32359db546b8f79bd4fa51e0d3281db5c35003dccb5721ae35b6ccce7fcd4e5991810761f68cd1de8a608c5bf5e8092c0b80a5a140e38d25c531a6f22c3d5777fab19d45b3c99c3eb379811aa894350de1dac5e56b4a9c6814cc3755f6fe3f682d6042dc26a3dfdd49db0c9c1d8b7715e569d18a2008b08887b12927fc261e850c96df996baa103c911adb7b6ec6c555d32a9887fbf863a50da7842dcf075e3bda2c3bafc6b00f718cc0b13c49c0f1095769f5a26462734027760da9305a1d3cf5d0dd12d4c5169378e6e581a47ec2d4fb2e2eba1d17f5908530c46f82eb27842c71c53a3e0661be49c59eb1739ac9bc20b50980788428c8104b52451e995f9079a240b464cfec5205ea9383f645be1177e821f7b24d268be1ea96efba86ff2f2e1cf0b7cb6bc14ef980d7d07f99a08ff55b7207d44b69df9287c1a336a8951693fe151c54c830297df96f5c49bf0e33d513acc26577aaedf6feb10cbb39e2fe450f506d03fdc13b25bb4ed717af38646cfd599d290bb23333f60844cdc54680e9b31c7ea0a080af80482f1f7f226b8a2abcdc4735a46b3aad774fc6dd6e374937c24e4f5ec81a1e902a2a22eec234074832e5f4a6dfd70cfa5bef7f0ee4972e578512f5ea9b8280603ed914fd2a0513480741ca9ff615c3521307fb91ff4a171ff90619ff552af2d40790fb4a8ff10c7c8ac4ec122d55a9ea169ba163b202527afb2acb789e95c5fd6ac44afcc8d7ba0680b37a9f6fc33a077adda81d93d2f6af434453616bac3f17e8305e374c549475ded2ccb605498363177a6ae25ece0c8d7c84f0f5b03fd213304c48799daea355ac849f6331d243a12af282412df9470d98845938af913c4b8466d4c382483fb8a597b7034ec60ccf50505231decb29bfe849056912ef4a678d3c4e3429af69;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h80f24551becb4aa3919808f42665f11a34893b077ea11285ee10dd9701ab1816fa49d43cdf9f0c401436c80266e2dd1227bfbb37fb04f46f32a7108d77a2c5cb4928f766b64046827617c2bcd9fdf307e047a72ad5eb53c72d8ef579c83143b3bdaaa723979759642b1b7dcdfe2f6d0b6a0b695b17a878cf82a80d3aa4d6fd64a5cd8dbd5bfd63c5c72810aefbb15dfb68ef06103355da327a0e0f90d73b1e71ea61c16e8b0328551c264a378c8053b61ccd78264b37254071cd358db511970fb7c55f956364972f2b3a2044dc2b122539e2c3e061ed11aedfe44ec6e3848bd212f6d40d097cac0eb80bff114cfbec496892715388f56347b16e74c72a3d56d9239e9e80cb90a51a0de00dfae38f1a72719f81d5139d4f713a4b4809215363fd61eb7693c7384998348350e1ad5e04b87fe4d2ed7f164cf12a9d516e0b081a5704862bd6d900718fa023e70c372d12e8f1a0dfbff9a9172fbb116656b268b672ea9d72970f9d36fd38e1bed985c393514b622b716e98e73e1a22e7f093077fc98511b6b30b6ce31079a50b55d7d5cf6fa0950d06c6ce0fff2af9b85297ff0e9ae3d5f015ab410b29ffc4469605a8836c516b029ed4bb9fea6f3de1a307f750714198072085d8cef1477d7a49af1adf752dcff7200888913abb8d0c4ff817d8fa49207fd7445720bb3f01f4afbfcb34c4e071a0cde8e1bd50701641b15e62232060cf6ba721b2a190364f2fcfd047f2c99cc46d93795edfc37b4a98a98a01caf4a20b2a931c1144de6ee8dd640731fb2dafbdac8228d09af114551ba5e7049565435227e680eaebc9db6d1e1718c98ef67782e2eef3669f5b5cb1cce73e1b51768a80f54e4512a64eccdfdf17898668c640d13bb74be3c2ad7f34bcdc62a7918583bc0cd96029207e5aa0f1f156de51e7807d1b1f702580c716a7c3dcda9172faa004de43cca7b30f4582e850b8f8002008e32554e9cdf66237bb0212d58b295018a62bb836489697a60d3e0a40eaf82878471c665d971c2d1aea33cdf40d0891994ebac57987f7211b305d846f60954f19c7ae711c8f14b9561b7714c30f5ca6180e2efe26d873f0c29a87665ed120df78174e39d6ca6448a80321da8cc4b233c9718967ca9c8fc3c2fea45bd7ddf3c8e04e3a4ad2f4d19c7c03d4bc5df286c0bfcd0aad0824f2fceea62f0aa2ac66690b205d9e2a2be040a6298daa60bd21b71e627fb8f22774962ec5a2aca11770467b4371e9ba770fc7e991befbda51f37489ef5f5ec6075e8c850abf04253f1ff037b1e0d798a921a52037420f8bfbac4c2fcdac1a3a7027d15091f5ceb6fac252c8d735b97d6232e4e9becf0bfba0d1549e3e8deee981dd52890250280d702463ade1bc8c971243b23e186918ff86f0999b66a3021f98020a07414b68764d4e4c73645ce0c94007182954c6d20cdeaae64b6b9124963e2e7c4f1a7b7fac3687285a451f5a883c2d42567b666ddb56d3197b8f635a6b383d7010d58044ea485b50f02f92f84aafcc6299cf59174131ec5ffa971ac41c8c9d9cdff8374ce7a29e865a0cacc74f9670183fa3bbb7f442a8c0c6f20aac06eee7663f2fc20933695e483f3166a8e0b0e9be81f145fb11f0961468fb4768dd8d371077f212c6a27dd042559cc7cf08a81fc6d8911836d523636d9aa8b94de7bc1447c3e6ebd74eda8d9dd75bf4dc54825098dd26324f92b6eca8b176b429050f2ab8034cf5cb80ffae16fe607cde9f9bbef37e5c58251dbb663739cfe0fefde773d06f1c8f4a14a2b85b6e840509dd0ff641863018749d3de76f38294dcbd8ae6e9e7c6d71b8fb5b4c86;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc6d16074d46c6f2f46bb3cafd4bcb8ba117793cbf93355a4dda62f6c2517c783c63d1e2dcee4a9669d52faf96e38c303a035335966060631cc19481e8b557252846003ed8263275a56cddbb769b289f834dd3b9685595cd06c601de64e95d0fcc86d9b0ccef397f3156f3ed4719059310957b1fab93473ee293374bd6533241b25c34d0a247e484688f97f7440e4aaf1f166410ba2f6dac660ecf38e22ef749fd115e83c752225d132f4dcd47fd5c487ece774e166f7b07bd3429d261c69dd97209c30ec68273144418512329865c8a8e4b88bda2fa962476eaa0b45bb9403a34fe8d261fef668ff7439fad28739b2305c4f03f76bfa91b740b2c70229c50498ae56bf8b05dd5f3f7d2c597a2c132a0b3190528ff111b509a444e3a68564eda924e1af974a494131c373ba6ee83bbacf5ff41afdc051b9a7acd10e2ecf9070f3351804902e9f4d41728bb77c8c2b0cd10f7f1e84b7f7cbbb7b28d61846c0df6fae7e35eae2075cf2ce1f83e92710e704751001a58f5daaab899ea7c01811ba0094c0336bbb62d4631f208c681435fc888cc457b4cf838ab8a21fb654a408d29fbbaf2c04b83b2f196037abaecdb2c6f09aa301811dfa6b030350259372716ee5de7fb20d56037367103493ded55ac244528f2000d80ba42a5e4abd89a939a00c12fb5b5706e7e9cf5bc07bceb62d5714b4e9251c6a393e11e11687a4cc9adbb58ca3d3283461afdb45ca4c97b6c3e149dd39ea273143f0005223a4b5141c2642747aea1b179275539e3d71d0b938eb77fa886f365a1949dc5e047d221beeba9541b7c99ced2e7ea9527e5c7d4b1bbd869f61c8ac00d4ecf333094742578cd079183b28adaaf95eca856211a30b3f791dc41ef550c5ff2e9503558d3b262161aa0db3560096a180b35c196ee1b96391d025a8afea189f0320a41453e1461ccfa5edb7d7927f1a38ab6bbc1dbfe62b4f1a2c225b093769d944a6b31af5fbef3e39dc0e5a5ff38366569429e296fff0add311c8066b92c80d51e6b5e10a1a64834b16a07c69f1234f0cc8b60ad5584636b96e83796b4b77f67192764e148c2d63ad136364da2ce4817d5a869788d9a52233b8c616c01d6fbf3ab4c5b74d1cf9834e0b3420054e6b09edc4943937feb43d8704370ba628998516d718cadcbf2389bd378bb37cedf2a7056410f4e85ce2c87c4e21a85639e44ab9b94710efa55abc74269a5979d4c019e9ffd00c20b565fdc8803b82b39947b0c325792b997f379877acae0346477542c369041be9ff8a4df3a3cf64ab5198c1cf3e72b00af103be0475c133fbec985eb07c743c2e8b6079df3dff86df81c94ab7eed76ece05fce4d4845a54dc97db69173ceb660dc48eae956baaea7d474272cda3542bbe193bdc732815b17085c394806167b9e776f3b6ae4623df7787ed14aa5e8c156e2b60822d9b7ff8d103d000a0c6eca99d8f7f66a67abede61530ce0553fc4a60bdfd1f9a676d4b288640797f5b0dc934c5aa183c76e6e5016cac2bfe1aa820a283c2c50667112ff9e34ef0995d0c253c9c9d05e419f370dd4d27de4bba9d8d0fdbb4b9b3e5dfdac97d73b5ba3514a8a07c0dbeb1aca872b59b60cdddfbb598b252c1bfc6f6814d18e9ce29a6d6a450b3e94dc1b11a80e53f98193f2c1ce5bc79a78b90e7bc66c4ba9af7e5991b52e7fdc0e9982b8b6c6ad8c3e722d2d8dd300e8e8b31ea827d8f00358afab3cb2448766f06ce592328b3b8be26aae290b673315b70db52bc249b9801d69bbafd0a13daecb64b6543a05f655e01d8a97f989b1f9ddcf88ea6cbe16105e2dddf160e97701b4f49d3c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h449fbcf9d8cb5fbaed87f65b321b1af2ff061d15344588df9406dc43cfb58a6b7e1699fdf70cdfffe9be04c7d995d941bb5de0b26e1e07c4c12b552b71cc250a6d3d7449f3ef0f5c1ea2fe69eec7e607c2edf45d8a0d66d922fb746950fafc340679015011549fd6e9ef701b6b160f2888852d9d713ff8030b27f6e1ad9df94ba46811e4acda0baf1a534eda0c6f5ce59f341364e580a931384aca04850a7be0f253323b5a5017a1c1dc5aac683e4a58897217df689482ca9d533ed4b819357a752f3866be3c06ea926757adb7643320798005c9aab435a3ea6c327b7450bfb14a5668f5111042bce0e34fdd0b723735621e1d6b0651f4e61d31f3ec6b76aef2ab4dd2f43972ea1620cbfc731add8ded4004358d6968360eea5046af9b875ced0ab7797d6c81fb88d41fdc6e7f84006827dde0a53ac76ee4ca12e28ab76503eab418b779d20ed72b9bb1667e0fae675cb47d60bb7b329746acd416247e018bf55560f1d8039573302cc65227db75fb1dd34bbec08accd35f7b802a0afc21184df433a4b9b29f69ce741f28176b9d1a7c374b1ea9c19ca0432579cd67cd8e26f1321977fbfa168f394b9ab62a00df09c2de391ac0a2f789ce788c98ede27a6b4d7d763f3cf131b2621d87802ab96ec23fef62970611c6dda268a4aa0064ed9e5529dab38bfa65c0eaef50a0e3b30ce790096b3f69000a990583e43296168c481587446c31a59a6ed2e9e58e45ccc2307ad6d24c14f1b8cb7582067caadc6908f4aded4caa2d16b3d6e528c3b99445e4ed55ae1d57edf033e3aada6a7ab17c81c3ff04cd93e34126c8f16f0a6dab013cfff51c563d62af3a4f35515f65c4e7fc2ecc99db04c6e008afd188e98b67b60e8660d8d098354a78bc4da5d9950c29cc720e91fa6c0b6fb3f57e23b156298ecc61d3c8566113a630cf2ab99f2a2bf01e465686f0a77b25261b896cc4959fda15445316b072686b4319187db571a058dc8833af4e076a2620fac1da58a2f1d3b1639bcb30655928a9a8d4b9266a4f0e26e70229b845d14b8f629da56ba8d9f76985630248eeab8787836f5369444f5d42b3e04840dfa4683714e837f0136a911d1f27b95bd63972c8b07ea9d2de271cc983e0a3644d1a2c9c0db17d3aa2d727190348c15a9f3d6eb8ada45d91aa0176fafc4531ce497beaf66eb5cacb8b9921f8fed398c3a90986260fa02edbc11ce3238d305fe3d85635ace8066850a419bf1dfcee7dc90ff3b37714dd91f63a1323dd06555d3723ebbe2bf006bf172359f59728faead23d6659b9f2df19e9e39252f28e2632ea49f6fde547491d108a037b8e9dbe28e132a1f4304896fb584a185f2194ae82c3975561f0307a77e4def41eb742acc38ed807a731427f4aea65b4f0bf9ecb6ced0db3733b545e0dd37d62dc166d5016f7c61bdbbb559a6a4662cca6349aed12c98b0cbc4b4b832ba25b7541950ea81628dcfc6a1dc1884b04cd153fb04328ad79ab750c2509b52dc4af8b45550b00e041b53ff691a75fbee096f0d117171853662afc8b34601a0055b6553bed6977feb3acce4ca33e58ae4f925aa338364dac6382efce84d4d4daba19a972adb9fbae43c37bf7591201f1e54d2438dd89e87d720b8c9f1daca2915b814435311dfc7ee76d438bc8bdf37ce98adb80edbf41821fc3a13480c9cd792176c910e846f1102ba03586c48f5f7c3282e465bbe6f3d35e87b0b61957b805319ab583a98b9f4f71c3cc9299c93247747c56dc22b4b8ad7f75e9b2f0577863a6f2ec1e08c6ca21880e2e25dd603bebb72104af91aa1c01f4da1321a4a3968959a34608c14a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h58ce6a764fd7079a8775b2c1ac86bf0417dd8768f1b28ca4e294fd936c1176f3bf752e572f99bcdf6ea89f11a31a96d7627184f793637a03ab4398881e94cad7d850d6ade864a1b8e97a5b31f27a6c6060c7754aff95e067b7ede068d368cc7836aaafb7c6b7698ab54bba62646d1de031ae71e4abe0c076096ee9c93d7a35423d6e3aab2d52d2bb4a8409250c010f87d610a48475407e57fcf657b143502b4895d3338bdb65b56f8bb7c44fd0c60dc7ea2c84139040fe3b57959360044c4fa194b96d19ee2d76b8e44537cf982ddfcbef95c4dc70f1068c23b972f886386b3db78d031d56fcf887bacefeb6b9bffc05c3d6a2fdf2131ff928130dddcbbd663cf3587a9ccc23bce26fa4f23aea3cdd2e556567acfbb494f00e6944972f4108b16c13f38191a475eae4251a92002575028ebe866a1c4c437ddec4b4767dbd43649e1a28e266070a093bac711fd719dc17d4765ab089bcf6519ca18814efb19be4c22ba8c9691a82e69a38a9147096f078dae97ca8ac4d9ec066fd21437aea540946db07bad33a8b560b43ac27f6d798d844cd871e8e310dc519be6922fb5c8a3d1684501dc068dc3950c323954f7866a4d876273100f4b487739c5cf68e8295d21b65ae6c11659d5d40a28ab42d8c42200f2a24d0f211fc99467a69fd738b2ed5a72f3f5e1f4db64bfcd2576826084f6ea80015dd3940cd8961342f392f32ebbb2df857adccbebfee6ecec826deca355dc044f4dc5b4ff82eef7c593bdd691b94aa7088834fb34ff486f99c890b38350e82cfa63dd68782477b4c22e9e3b2df076f6c5297155a3ad904e01d609f3dcad51e38ef736db6850937652b2618b8aff061d9ee88ec653ed5f5ac876c9f18c840004630cd62477d2e5e9c6aa96ef463d042e1f83774589e9b8c563bdebe6c471a1f7e9a73111ccb8152bfb53889e96f0079553ba8468b3ce50ab284d1c5b824f71ff7a2eb0c6fa005b65ad629048eefd64a45b8d0dc3e883010d49383d6ea62bf4470ff0706ca9589704a10c7e4f14bb5f4e08fe2e6ff5d063b595b5f8ddbe54b27d168da89dd79d5ffff760b89f79c22a8908422a0029b77fd8349bbb04555e909cae8877474ae2746d4461fb9a73cbe980319641dc3d400016cb999f11209fb5bc097895597f24f4b070b5ff0fbbfc9482efdf6fec78f25b1000cca7cc1e34578f7a0a4e83dfb80df997f4637760ab579e7e98346cbf71543af06941938bdf2509c65706683754e9f599e3decfae8ca1760b0b97c1b878ad836df1ceaf8032a998fbe81651d31e2bc07ac5dede9870cbf330063704dc6b4c5e4ff52c0c495f73f0413ac046fe1b906c1285fabf9e5f2b00586cd8bffc2521d62d7f3ff12c4b5d292350f0dc46e2002d52307d3fe1b57c2ea2f3eaa5a254bd49bd64d124202828f8ee919f9b8d10bb062e6ea933ed8e8279c8f6c050106e3ab92744fded19d0da9d1a7b2ee0b0e34fa4e870575c5868b9661fffb25fee5012bf0ef548e0608f1b3b5e3014ff3b9f818ea68fd36b1052d459d2b64fa29e032b9588579c1bbd8fa5a7e745e9b50a25df54b04b8c71b308a05bd5ba7a693b981a9ee7529d0772f678df9295ece221538a39ac5ce28e116f7707e5d30f7eaf8f84d6aa51dcaac6b306a331cc3916ffca5d072347b9fe8c151ee92d6fd572101585be2bfc3ffe455d2ffbb6d4746d8b24dfb1b150396b08e074c591d74dc094547f0d6330c891aa0dcadc5a3890ac55bed5466688577bc14ced1da5a3d99449a0ef6d82a9fdfa76574339bf53f2633355fe50db97425a1b1399c9073e8320d7495d835d3700de20b1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3b298f433d3a26b4491fc9df49e28ec5ca3515a2fdbb3cb777d78cf3596b66db8d4ce4c1262ec053509017fd991016d0207e33fecc7584130d0ea14560abefe2d5ebb37858ab09106c9405fdcf538dccc7604d4b86aacc3d3d2e17b70924003753022d713a14af40a6cfad3d2bac1388eb646c7a74991a29d707297a87998d51c82ffa85ce26723cbcf41e6cffb3774deede40117a0409fa5303b21b777e02c4e06dc16b5f7bdef4d33f873c84645a8554ad0aaf290aeb18953b2aaa42219ce9503eca9135d620b654d84c7790f0bf0046b97d54ddbafc431cd63c1848afa7a7aed7c6bedd621f2f44ea4a0593506c1d3666e1754f0d47fea68fd3eb361ecea1ec8d50daca20bc81b3021910608007d2f7d8ec53713f96826de46d86a7a3edc9609350627f69ff46efea13918e38abaf0959bee8801f0287fe4fbb2ed44fe19c97df47288d8e5212edea2e3f310077fa0b144fdb62e4a0ee434d814f80f52182b4a5fa9f71eaef75270675a90c488d7214478555925766958b399e0917158de9a3273e4957494312a022c539d68c0aa4a50c7502881a904a7e8d11b58c39329138941a4c8e3f431bc2ef84578b63daadee96564ea0ed47662beab53017230937ac8bcbbff8a2f98cc780a83fda1c6316a55232265cb5bcea7afc50873c50a6cfa3b10dad1df4fe8f79c4c16612695e850d5f598906c272f96ec0e2155c8af1cc85c329d4bcc3f03eb71a683a9353f455dae28135e7268149f79cba4e9cd6d427bd1b170785992128b7de1b5946c29580c2d743f4b717666824a6126ad96898b3ac7b2a35528398eee956ee4ee706a0bf792e0f7d72753c887c5b6d42299b07461b65747178d455167ddbbd90af5ab97b9795d025819f049245cb6f10209fd69f29aec5f0dae0e252b28d3198d2d4f06dfebeaeecf5b847318f82b472658bd97e4276cf34e19ca0954eef9f28282f71bb2e107c95a2c2ce25c6fefaabdf26c96bba56c827c35b55ed2ba6c1ec979760949830e78fd6193521d801af1d1f28b66cf7a6b7dddb4e2f307ab8be5a50072d2249c4188f16b15f3c11802a6fc0e60f9709526ff8f4377f20627a26c70c20406637aa392fa5ed23b4e482dbfc6063b5e0b037a63f3b60d1ffe6f7258f54490079d76c14997cbd09f455eb1ac74d7f371746f22b7777fcc299a0e8834f55423e663c653cfea387eab1e5fccf9f811dfcfd40749159a48d9be3ea1ffa7d822074c47cf9577a829abb2b7387caf9f9056d09e0ebe95f8c96f24bdb248ce102e9e3180cad654fd4224e3cfac180bc1277e93e97a2c6069e1f706ab8af2fde92f656607ab9ae0d5540ddc2da43a2c968ee6fcf0e89fc0bc0d4fa2f660d71af779d58911d16df7718a31017c536082ff8803ef4dd31c8e558cd11547000f18b08455cf4b25460d5bd64c1e2191c3578cc96fab8588d288668452692919965d23e6d7e8c9ae50c7093449709b6e6bd40406bd35b98b0c13dee73eef701d8654efd9e3f89b76e2c48f3df67361b487fbc0456c56d77283b9cad096f235722c225b4a376d832da4357a2140acfb96d383bfa8416f36c6538182d0f0d3471ead3d8a29182c7b9a069351c98183341dec0a244c890491c6ff6eb2a61a7af93445512b21221ac516a1e7aaeaab74109e74c9a9a55d3d550950f43bcc65632f21e840f2aedd0c1fc8f90a2c517db461ab9fcc366e1283c13bd209425ad10f8f5fa66634d5de0aa051bf60cc4b4f5e54d29a1ffe4ec51e06d23df3781a53652e647f5ebd0bcaf75c02839d29b026700da134af5ad9cd08e10fdbb7eda769a820b45851097288848;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbc040b48a4e30d11ac52bbbc2ad51bcf4418b31f3dd325145b7137829929343ab4891583b59840ae3d3edd6dba5e40d925e943e8df317e4745bc5d04f968002b45e008035916d27bb3541e345139bad1b7b17ce1e35c77d237c6eb9f775a3826a07fc0c22fe902b4a25f19e389260d4af7a015c853d08808afad5d4ca59063e1d301f1ad14c86c8d4cfd9b567b3c61292f58c23bc0f4241be24cfaf7493883643fdc343cafbe602b534f1fdce6216d72bc85df9ac6688c29f34062b8ac8a8d1eea0f4dd76aa6a2f5dfb6fc99f2de032293c60b28968ddcb16b2655545ffd90da0b79016ef85f481a986ac7af475d928208544772b9212d7d7497d097b9e7b699f7542e3fc4fa5389d052ee3e3fb2abef59e2db12ee2d07559b1862ea7c9d873643061f52c3b42cacf55606cc930ebd65d905af6db76377e3e5d469a8d6ccdac11a0e2d79f72d4adcfc765b1e5ee3804016159f67ca9f85751c9c0c0ba7a9c957bd3267faa6929da9ea544ad2af7b35296e137eebb178ac8de4a619b74e7280985d038c3fe48e56918946d31974314ff9b127865beec16ed4b0423cc8729af0a0a9f9d287f0662b29371ed6cf732cc93ecc2feea18dbcd88c2adeb9d514725d58b767821161912c4e527159be81ca0f7e3cebc10c9313a79e5b77348e5206fb18ee470319c0cf6d4d65827ee8a17f606cb865566c18fc84cd5c65234ef6c7a64fb04c11f974a0728e891a69fd3edf4c12410d692e3bd5f05ec08bc75f7c612b6a2e790e95af7e2faf2bb4a17f3ddbf98f667b86cf46c1ccc33966856ced14f53f4f3af416a6bdfdca63402682a5fd525eb52b9cb7c1d1ccd442376fa804e8ca43dd3246f0e60750a58c58cd9a763235f5a73e6dce6166772c364b362aceeadd9c7c2bb032a33cff0b7798d61f9dedd2e3ba5eaa82ef772eaa539c2ad2c4f3188fd4ae83268d788661714ac563042f066fafd4cfa9ccf8fc8b82cf3ab862f5322fe09a407ab531b4885c82426e33e2758e250e18d3a607e3e16dd110c8dc26e229cc307200fa33d84a221431b4148bb52af9cdd8d060f9a6584022d3d04ac048799e6571acb75f296d5074e25f54afa640f3a587654d0bea55ebfc7629c0a3e3bc23b9aa245cb0d30942445c87fdaa52bdbb6800151b732fa4bbd0e5e301907e46ebc369d9b6393060eef541d83e1945214cfc7077d7c7df9eee3db08c101c1eb7f5130ed9e8da7c15312efae4fdf5572b7f8b69345f3da5ee5037b25507556b57b84fd34f78b65066283dba379c917f297ce3caac5200c6e190b4e0961b6760b6649aca84ea64607343061ff1566cb0bd99bc3a500a437b97ea9bd3c59b78b856f831572a505f52ca85716db9bf3dcc09e0b13076eb7678d0ca8f19950d36d0382817b5fd751d8180ff09bcb43642a3a45b2f29c432bbfffbaec60a444a5f2467d4e991233833ea89c697b56a67317b18e89e71b39b7408a314c66c510220c025e649e4d1166d4833359a4bb1a6fd84f17a2da69bf2992120bb7b1e7f2b32c4d127345c04f62a1cad7ed860d4c344ecea6e794e8a8c2ad160d7ca9ffdf751ae8a9aae90ec316eba726b25a4a8459c40b4b18f480460ad7e7386aaad9aed23455903a0614257019d0026ac15cddb00596e272153dead3bf65beec7bfc7e7d99734d5694ce1ffcd0539fc560a9b3162fa571a5a0b536dd85309dbfb5511215078f94bbc135328c8fa4764399d31d2a881332cbb7eafd6d4da638add27c6be9d6a6b67c3a39c36c13db4b70d96a0f6f6c230609c38767739b54d4b5793a714433d0846ba036a9e4369a6a41d92c7a539d2f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h821828b71c06c567bdecb9e5d64d723d7b2f487613bf88605947502a34901a3805133207e869b9375ae2e77256a705c13d7f39ae78e96688eba073d4750c740d7ccdaacc9e691b67eb6cb96f7563964b966e25699bc91814e8e4f367915606d6decf628549315dac45ab49f2f09e61f39e428aaa5e5300338fdf50c9be1e11b072c2c3e660bb7d2bb485684a6ee5618236f2d8b68781dff95a44294de3e18cbfb875a6b11b30eef33fe73e6fa9c527de5c167b341ca855dbe53459abc6be935959310b174a9d8ce495f8a3fb91af0618df34ca2fbb83bd0639e60e3ee92e7958954bb7c1daa6c6cd26e1aff1ea62c4b72e075d59c6fab3626354ba3063e35e37527d709074e8bea07336ba777b04e94bc280f4e2b2fa18f1aade1193cddcd40a0210e627c179cd83d5889473e14f8dab85ad3182936367c386e6197c8b622eece765d9210457b15defe0c5c89ad8eb038f74b6a77b436a0f406396ef5e2482561a7d9653df9497355746e8fcd178e5a08728f9bf309d9222926282d2dfa841849bab68b4b813e4c2c3ea0baa73ee58388aeb675cb76dc51d8636efc48fbf2f197e515ac31e1c0fa0b0e82a55d415292b74ea5ea9343a18a213071f0ed373cb11da26c640fadbad095b6017f5da96a189a24802346dbf468d6cb715104a4159fe81eab25d1912395e5241e412535d6390d5d39f60e0910dff70b54a4ed954b4c9ee010501e4062446227000fe7a0590037cd8d75c58da8aa617d9d828aed284ee29aadfa906886aa4963d50b2f06682d37300c85443318850b6b7b39e2f0fe74993c62bf392eaa99a926153e1a5f1a6895995082150ccf4a466226bd7315ab8e20fc705881586b7d61e629b96039a0ef060f0578e8de22a9aadfa53500546cdab1d9eb695f629aefeaa5cd13d1bedc82c5dd75cf86aa48c7d14b85315accede0d99b75b9e8014c575abb86a496059ec022a6333efa349ffb9fffe62a5aa3935ae87f3c46b10e39229d5d6055666b7ffee58c9ea2964d7663e38ae01961ccaef49cff6b7eb869e66aba8fba1d42d044908de6c15299763d9725975255e59407bab4c353b7c07f068f83e7371ed7027542fa5dea8c6d788a59e099e79ad3b5ad1334529a2d1f152f0d84ea8bc82748955cbf97f3b0ad65ce4a080fff624e1f4e39f15b33f9ddc4dc6993c3544df6072b16511341d5e5014833abc3a1569c0195eead5019e5b5695ccfbd950adc2c45ae6f7f3870676fc4b8904452c110953809d3081f8808e399c04be1a7444c212c277c68f5ebb769b62e7e49071af045dbc7cac60b970fef033c2e0a0d17a52cae53b6cfe39a22f600f1349351dca0d030dc8ca331172d908e28f32caf217b9813130c29e8925d924a97bbf2f2a811134be44ad0d6ea5b1ed9f1f129ba0aef0fcdbc7e0f6e2e2032c15a3211e0adad23621c8cfdd52a93f29a13a48cfc222d9b1b32696122e3dc4fe1f17a599075b334c63d6fed4ed9e8e346edac45574e4aa1ab1c14e5256ac29d0ad5b106f4700b6aa1250e1f3d455681e3bbc64b878b661cd2cc85209bdad5219279c733d1fa8e5f73fc18fae3d5baec26244ae777ba81536c9a82fd85491a504f5a9a6c9be0987eca1006aed94d551e5a8e2d650f8d3ebbbb4e8d6caad569c01c018ce6b044df3c9cf5a24aea99adcaf549d7693b12d53a769eb54725f1fb8fbaa618b4e9fec90bfac79232a92c01678b92675ae50ad5dbd1bc3688930339b8db9b3d19ec6a9080e856a69876ec012d1f986ade80335e01361c60327f69140b9b8fb507a9ff3ace60286b127372c695d54c2666cc2998546205eb9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h96c1174c9d9d4ea928125db08ea97e8132fb208239d7342deb006a5f4255bb3f4c0b0e0e9e9d257ccb1c44ff2887869ad9f0c396bbd6979fb6315a395cce0c597c6b50e85218b9df05669427dadecbb980f4cb61c40b0a58136af66a29bace29d2fabc5b1bacac00f5c7eb7fe4eb580aa651574c707ee104b42e21faa8f5693b9d65a0879c6b496e0d6f69f05409954ba30c150f4c8ded1d47c3680f2f6fe1fa0545c46198b0d4a9975dc9036aaa9378703549d6c90cb2e33a6f38da39ed4d1fe095fa8ca5604e09f5415c02bff7d7e63a7dbcc8323e319ed90f219ec0e97549aab32e007d8e407a7019a00c81ff912f22b25e4ba01d285afe66b53204e23436e1e63f9b78c3dcb66493677c421a62ae1da66bf34063a95a9a4b921e255af3af212838860d695b42b690c4e08c1d7b2b035022e2494cb364c3ca8a77be43213ed63dd7f651d4151d36fc30eaa62765091c5ebe096ed1daff62b68dfd8515bb8641c9408424573bb3e94c071edb4461dd1524b3398033a0264ddb337eca58dbbdf5cfd7915bdba3be1bfe3dbceb3b17e14225fe79635dd0ae8c968db59b796da51038f2c2f17dae8be6601e3de80d5eebeb61956f3cbf14e6cd567fa28101a05de318fe0649ba2f260922b3398f9886cce18a353f7406476ec4270906fe170b61d52d860a8510f700dee0954582708749ae7a20a6ce4d4fe21667de0d0868452a6f93a85d59fada1a4c7862b98d9cdf7c2bb2e2018bc3dc894a15b3b4bdb4a08de1a6d11edf74adcd9397762531aa597b4cd0ff7514bba591d654ca13ce11537b495fd19225d89b83553f4f1ebc05cae5709786e1ec8fa4cd85cbbf7a02b2964bfdfef69b7aadb224c60942bb76699da8a73a3608b30a0d5d1ac0240e364561a5bb28d6f32abf3858c902c59b047df3a92363d70ab6c36494a22d5bf8e658061261bc28298bacc47a1ec77545ef6848dd4d886c344d82a8f7cc7ede36e4b7281bf211bca01be7ef64f5eb694049fe2242da1386c4e6d4fed069b69e6cafcec07bb37ac0b189537ce3e15ada3374c309af9e1f871fb74df87a13a5d444579d1f7cb8ffa1b62c5575ec8f3290b1565033014b56dc14605965a356aa97175d393d5efeb7df36b4a88b57762e1dbda363b5e110cef30161abc2eb3c82e3407dc1125d1ea48ca8bad63c21b1b082c4ea5f58c411da2e11c7276cd3f916d7d3e34a87fbe5d8a8a33674d4049a5d0414616372259b2bdbb52f67a277c955494ee3ee41134c8e5f1d93947ae7c8075176725b83c0f85ed184d5b07a88cd448d967f656ac5e832dde780c797b0767812021c11334aabb907252bf24107bc7f71a98b6ba92d1298cd0798e4baa0e7764260f827885bcd99a49efbfb34b2fa62addb2beae3c6e98d91d3b6fffacba81a6750d4a9b5aa041732c5dc1260b322f141d4b3ab2a816cdd88e32f61cd7ed5dfd06f39ee9b6bfc0cce8a362229ad4acfaed226019c9a563ce3d42010e1cfcee38be8dac8b61263e856a8e01764bf8a1ef923bf26f92cdbaf9a910dbf412e792661d4d09585363a6558e78a95873f4fdad9bfb1c741d6924d91ce4fef5fcc732643a71fec140d682b644527c18721d169bf2112f954d2ba8821c3bcc5e10e46f4dbffba08f22c0a497fb3c312a57f63ac52dc0c513651b66d6992adc250eb57dff55663481d2642059423fc856fd748d3b0756e6cc64cfb2e08b7f65effa2b59325bb8db2a42f50fe24b40930af19d0d16074a0bcf0032c992909e1f32eb2a02df8edaf290f52ac6384c57bd344577c3bdbc5460c92bedfeb1d44e08ed627b368b750f963ff5d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h757bcf83177bad3e00ce53d2bf8db8d53d288cd58525bdde6ff0ab762558d32d3137f3a965405815a9dbba8eb236b67af3aa79bfc775a5b7689e13ded1cc384c418fc3ebb66f81ea38915e2feca35d94e40c4ea7c7efae3acc602f7d321592ad6a8de1b4027e08b2ce4344cef772ecf8b4b22859c247868dc8ca89fe851771d8a2b70145f660efa6176c6f12411ee0aab0531096a582490f0ec59b3a27d9d93e4091adc7de0666c33dc1c807ebd3c65a390a1ca7b882734f67ad2bdbc4e19e375d9fc65f7d440daf31850b30df43eab08275b614a19afacf3b3ea2d846a535ecb49ed6ba658326bfed320bd8ab0400c14126011ad0c1e201a76df7ac1b2993312fcd54cb95ba59c915657cc5797ecc71792fa48dbe8faf0fa4049c8b3f7f9d4b6515bc0d987d544ae9a7a8d7d793cbd3a13a50b0f6245a95c26c04a16705c4da6ca09d05039465ad98c801c4071f557b74b09dbfafc8ca01a83d6af0e11270de9099d128dae78bc34c4b8a342a2a7d510e518047d9ba683f6aab2c90a958749944bf436339dba1dbf0cddc6bccf7f1e261e00106e3e3acb094ee0ff20c67c648c5e82cc2136dd3cb391ef2dfe063263ae96afb820f5569c3baa1a7b3b8b76e6684be8856c3707cdd1acbb4d00de519c15983ed40f589d2fdc0869ce78e440848e2b4cd1a5ec6bc6aba331c56f268836de6846b547aff33f3656991586e338f6845c01a10bd21ac39ca849a1e1dd9f9b563f6a462625ddd2ac7e9b857ff548c8fafda8e5488883c8c7fe76ca8d5679b52e4357c98ce05532aff73b9144bfc9d0b796c802bcb54dd9cd87d059300c6eebf7557bc454910b361a701219882174c349e2d9943e154b1a66329395c84af8590d09fe88974baa2f9a5aad151fa1c6cce6c906d74eddad320a5df03b332f895a37626fe0ed628fce504bb047d38ac0628ddcecae95b0dfca11bc4a7c1850606359fa128e3944be571d0ecbc2af800c96af8b36b560dd1942a51bc40bc0b4685afb7410fb0d91d9d1c076f982039cab7b49daa7a8e6c6b01d1b53d43e5c02ea15c050e6ab22fe21acb931be7995e9724e3efcb685bde02887070c0376cdd67391b03315a3193de4d7a49543719951e23626d785ea61f818dea200bc195830f5af98e49858db6ca6e3c2c697c4bd6830895bd9bbd05069b1eb8c12452e241d1709e83da99a2cf958169c6716a8375587ffad66bf3d0ccddfd86d8c50817c78d7636fb5ee6795f8c1f9c7164a08c0a12087b5e21057c24fdd4a59920e5a8f993c1e0cce2e422c80b5e7bf03deb8b89f940814844b5ad52e2a20cdddaa1578b8699e3f1f69b10f3d361c095919c79ef4511edfa871a94491476226eccad6b204fdf214650dee0c827e0ac84b8e20391c1a1713c4b6944d3fd450c227635fe6dfc18641e6e8e74a8070c7b66c51f0b576e967134d9cc05b3edffcbbed937545893a3abb8f1f0cb116ddce953d6ff876c11d6cca368a5585bcf2e5052d9dbc1cabdd6b87f0c9912795d6efd378233e1fd5d47ddd9c4a8201cf7c575fa80db17993775734231997a548e1a26cc8aebaeb7ef77ab4e8f2f6e6181fadb7451ba6faa857a9451879ef7df318ad82f9751cb7c5cc7fcb8d4825294d7b8853f86ef6472ae3443c7da9aa5974dc870f3c0dc24fd2c76574f94fd4bdfab9e947085617414d5c8c6767d0810855c7235d743541dced8315a40b7dd71eb5ac4bb614402f631f4652f8cc6c09475376260460ae60cd123386fd61f382f8ace355b9928a4e6c88f9a64554612fec5abd72de1be5d06c33ad2962f721b8825f6d65e6022f7e820409c16;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hce1b25ca493a4568110e43065c46d2d85ec1494f187329d8a5a0239e0b72fbecb5e7dd4334e12eab902078aad41c30eb8f777d768d0675025680cffc5c508ac9329111935da026da4f4f17cf568c1a40a7644eacc0a7b0cf7f1a22bd91bc9aad5adce200c91b2328e3464f544089e821c4747c3aeb455fcaa4379ed35872a3a7c9f5ee0b10416a474986805987575ffb9569c0492ee63d187ce6308064fe6b975f8d2392fb426568c980b42478452301da8b5476f2b3a7779c752aeb1498a230de58c9cbd291337146b61d3b89c1fa4eeb478bd0cbdb1f6e9727e15f4f6985cc1a1ef5dcfb90f98e33e22d687990740aee8a2039efc15c4ce4596168a11f0e83c47b5057c71290173a3c3fd7d13ef2e5266860362a5645064f010534ea0884b713a4f37312f86d6819c544662f470644cd4dd3215095a4c0c02969ca8a2616056865d6203eb8e80cb7312225fa0293ad3f4ca2b4f4033a26431d6fca010306ce9d4d907e15a7d439c3b9fb8e613246423fe65743c3e013d828f2a0e435202ef40b2bb8f8b9add2305cc1476c0de4286c0ff86282759e4383a9f8eba7b616a5e8ec4c235913cacb2495c590c1126384b5a51a776639d776a420420c1854ff47e9d822bf137958acf03c5f956f61d05d90905f9332a09346ba7c43cddac62c74813794be5b52f87e4eb5176b37003efdbd574210b658c5c5af5bdf7ea866d57dd0ff2dea19cb87f04c1ee9db1d3c03f117b39610a2107f2cbcb9d8e649d91769dbfa0cce4d512ad3d35fc145d2867414c74282c176bc08f5684765e5f61abfb8371759939c542c3ea2dd59441852df41d46005be9a23163a3a68411725f561c94cae22808d2f77a221cd417c4e9308127abf6d80b236b787246fe077d4db7dfd81f1da63f33eed306fad18f1a0d4263457580dfea7e933bed8a0e328920ea85592936baed1193d3cccf150fb002ffc7e195dd33ddfc3b5ee2048b1f632701b78f299ff7a7872d1d84a3d23aa21d2a5395a69da1fa2aa58b9a47a91b79e3be24ad4a3c4a0eab90aee1985963c2ea7fa6af318b0dbbdd1d9a15536413a32a9a3dec600692e5dbb33e637f41cca39d83db8a0b02ba71366188498e76a8c8d04eb81a2d4671e28a080c8647d53b1b08ab352e81360cbc481474788c677e7ee96ff5d922deb690298cc3b6b31376dfba8456f7459075084dd1a9119963e2d754d2773abb40d813100a699f6c3132c178f25cc71c1cb21819ca37713dee888a8c5f83d055ba8994e0967e9d2bd5466b75452683dceef06ab8aaf1bf80201f2f7f8c1b7c952663761c94507cd13716760b727e202e2aeaa0935f7e383b081f84f412314fd94e200c79d3814c9e7e8076bf77309f83dca4369fc5cc7d3a3cfa32a1f52d35dbf465344f89cee3881f816aec83c2afab38e32abb1c14a8a9f36f6a970cc682dee0dfa611e943660f3ab8d5e21bfcadba8e93ca8edd32df87f4fe70f0fc8b703f79fff3a05adab20df31c7c79ec0143dce3ce5c20cae7bf9029d613aa9957780032cc69cd91e70a6b7200d45112565b41725e027a00136cbc2e070cdc574784377b80b10b2b01ce147322d69990fde5f45f12fb931dc80e95f7191462850a05933454e49824f19db08534f587beca30c073a6c98b4d8c40afea3aa7a32bb1d231cdbd6dedcbc2345ac24850ef3269c24e82ac6c4f9511f4db53c84463d9adbeb59dc84334632fefc33832621bb3083e12fd09f9dabed5339714d5cb907fdb3fe60b8f70b240ab64632dba31833097cb730e9dad8f761608517cab860005fba77cae21d1fa823350e5d64d8067a6298b5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd9c46f323ab64c14d56161e1e5c1d5e95d3ffc7d3d05588f54be9242226b7e17be2364f20457356e1112656eb39b69fffc38c4e2f827dfeff66349c24c42e0c7ca6601370aed5d6f814172c2230b72862a3aaf8d294f18303890cbbf154a366464756c131f9638c85e40155b3585a4a9b7e049aa3d7eec87432397f311a4d146c19ee1a2ddc2713619ba9a4826def22e26ebc43a13cc32045ea67af63c08077f0fb6d17e91f73183f1c102ea8f4ea8e9d572a855caa44f150193e92c1b36fc38138308a044a98732b450eb651c17232e109d43f61acf3b4ab3cd5dbc08565e695394c9516c396d49d8a565561ad894827bf3edb45e243acea06e1cc1926be5b9469be10e14c59cb1d9d0c7bdb87149f193030dd4bd3f72a78f975fe8c47a103983239048c6b42cda0d9fbbda4582fa86570887fd7d3aa270350b02a337e30722ecd3c4f9bc7c636159a58bae4b1d22f709e105c8c5e9fb02bc20942bee34809e986a53068673db41a05e92f7a339c29513f9336ddcdfc0ada4bc90a5288e8977a77da6d0a1a8512b95298532e1e404c3f2b47dee9fe1643914b9b9c827d78d0e9156b918ec82602dc0858d2380232c81a4bd3caa95a901f6919ecd12af79456ec986a4020de553d38cd79d41285fba52cca67023bf1e4ced7bbe5ce455bdbfde6f51cd1861632804fd0f748bf80d1a2f65a283cf6570966e82e97eecdb35fcb18f1ee59e860b1c55cf3cf0d6dea78e1045b9a604fb6033640a7aa24169874abfb3af59599483de61dcc89273f4ee18487b43df1f852ce193db7a99d07f2ad329848be105a375afa1209255492314904b609fa4e9fef27e294da338afc69b399a6d19c9d3625b8a11d9b4f04d5666c0d1d7b296f83102bbd4212a90a51eb9aee1358a2cb35c69a65d87177dff51fa0504cf6273c84b8a9730a3b82410753572abb1aa0716f207395881cb12889919f80d38cf4f7d832bc58ad2687f9e9b2319aa633c06443dd9a2e384ebf846de0c225fcb358d4d8be4a0b1f288631047b7298f3beb9ca21d4618a1a7ca9b88b09a70e898ce385b55bde34d3680c0a2a8be68232a460808405f8be796f71fb245ca1d21e73e8f3149577e6a525e364ea1d00dab5a05859d47aa4b20525c6ec1a42c77ffc6f9cf3fbaf64ec6f58e9a3a55e7e580559f8e049f4f4ed7ac1fc770c13fcfeaba358e948043def4636b435226f57e4bbdc99852d61acae36ea31e125e4f8f63f9539373b33d3f817abd9ae19915ab733e46f21e7f20710e7dcc7f06c10e75c0152a63fc8ae430340ef692926092cf70a08d0f6d20798684bcf792f8d53b6e105b88c7cdfe7745f9c6dbe08b23a9b2683d7a7720e6735ed6df37ad4a6c99ef15c669f39d073e4acb82e5f6488da1c3e31a953e732e7870df43694e7ea922e71dd341953c1d325b6b5f01242e25ac0f2a34e7694aeb075a17e4bb5ebed28bd6cc52656a2433bda0510c46d95cec68f6da9ab6168bf206ff61ea49957aec622723181fbe9ef3e619cd355965373f4133c907192e3dec28583aad899f6d9296045f9bf2d2996cd4b2a512b382551bd19012ae42b9a2ceeb9e34b6b0ebca4c7a18e73068017b21cf9858345d6c988e0b8768f84b5649aa16a8c874bb4a4422d73e440718c3da7507fddc2c3c1fd36693a425d5d63abf0bbba46bd30d44c77823e2ec5e6624dc6bb6b45b121e70468465658c4c968dd0f79cd39979f8ac649b1ffe8f0eb55d5152e392bdce61db8c0f513f51b2ac921ba82468d45500321712a7af6b7c005462d9f7fbb6228c221c06b4321763cda3c5327c2b89fd0e348800a0ec2e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1d43e2735f52fd9cfc25826104a47f4046f0875fe68bbbe256450c707a57b91a1a342c8b61897431d5fd92929fe2e693572c72f0f8795e818fff40963a7f395768d579570df04db77f41480c06987a720fe17a79443a2c312ed62f8f14957f691af544300c53304e73cccda1766dc0674fcb1834a7b6cf3141f9271ee0f2e7c61d94c221205abf105c6bb0117e104fe003a46f503856f398e4a94711ad4a5114fdda160f551d491d6f44a5e6d993526c75fb29ae1a6e78272447eda9accbd77063ab1be7766ccf2ec1ecf8820afa426473686b705ea71ba79539e560e94f00470ae8f146ed278a0b96f7f21e5b1a6767a1a4ca5766018d66454b0565aec9be03be4a34ee63d7e6508683ae1ddb3c13cf9cd48cd403cf7785567bdb61ae018704e91c742fb340780c8f58889fe23349faf58c3a80d337b70b0ec02f5c19534e524020c8b9b70aba2bad2b90e83c2bbba1ee05b0ea95e514d71545fbf0b4d347d91db0e605880aa0c7da4a29c0ddded0687e3849b87cad9a7441b359b92261a73770ba317fee487f0a49ccf4fed6f47e5f018ee0009b2dea5b426c1e3ef7460eacbd5b458c05c177e775e10b48eb4a9af64f8427c4bb2eb2c095ef8a3df2249f35b3cc6c06b636ef59d7d27ae06b66242ed535bab0dbe70c98541420675944b42d6eb59150a658a66db00329dc1d1bd222263dd5a21b585d8536c60e44bd7a14d3952c6ed5d9ecd6e45f6661fe0466ee2d1a3005159d6a44b5afaf4d4191e4eedaa51e361846f585d09cda26c41c10c6a79b59151c5c9594c899c02e30f67f494d9d76a7ce558c196ef2a93bf0a53ef7c504eeb32e0b9af2647ba23fd1be7d6ce7f2e4670bd3272911a30e49a8cb8c7fb128f6fc02d2c0404e6ebfc4f51d28174b7b3f713174051e37980282d976c18e5d3ee60725ad4349bc9e112a2b4da85a25dd60e7059b36960605020692053092645e7e8a13e6323853985a8f5bd79a92472a40a94c6761226a4eed191b5f619267469de92a432932ceae3ea3708f98d82e446d19b17665e407209e49c0b72e6180fd8aa6cbd2b0e28e8279373df1adbfa1bc9efe01673a6952fcdc871709eed7c3d4a06736cf595ba1c0bab63ad6546dc944541d7d200df6590473401f594c4d3633fec005157227647130a3fc475861c6577a8767b3751d4a81c5750c68dd74cdd63e38db44aa13ced43df71059f96c1af26d93c1be06943767fccdcfa3e95e6b7d98a0018f7b484eaba377cef5684f6894121eccc25e11ba5f3a98d229d45654e6c814886487ccab69a81ed88e479f52091bf24514169b9728711265c333920e8f2b66f4198833f1a22a0ba37b2388f930f2f3a1cebf239ee4583af0de9fe7e73479e6b4848cde8753b1d91dbb579a8203839dcb635facf64a71eb92250fcba2abefbb6bf3dc2955b4109169a8fcf726ff1d1ea2b7bdecc379a4f26c2927f148491736bc14bcb8920552ccbfebd6eccb95c5253bc1fd6134ed042296c9882497512c7a297bd3fef500457c64c568d54ac6570d31c41a04975cf166dc68b3cff3a3f0f203524af75e341e5c7b3121d69c16763136874e325e520253772d269479b176ddca5a3fa3b593a333be987386e5979399263630c840720aedb74888d9dd74733cbdc4c1fcc29bf0a2e066917d5a2fb96116b283c6e499ce98c0514c4963c8e922db77bb48e22bdb3c34c4a06e074e7868aed3ba3b5d9f82c3e097687a81e07fb41b507de4ed641a5f84262d809daacf7e1c4809b0297a3f8939b4e2f34ea40325652052d5eee05e29722cba6ef24431429db295dd7532150c67baaff451;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h90ea1bb2f8e13762ffdcbd110e4df9f672192b88e00b1402bf2a6654874a91a811b95772a68353f47a64d3c3d2b0a044ff564bb53b1341fdb0f636bcea8250d4fd8a06a47b896df100965ac94db8437e7de9f41047127a7d0b6e7f8c264755d08f326cab496ca42eb70153a0d7be28f9b1c0be00d0604558065cc2cdd93d0b4bc876fc22ca8e4f413c2a7c0a0d6b0ad4598e066cd6e8e4329dbef87bc9f11b166419d4486d0e5119ae9458258303ce8b82a9ee158705b48e49e2eec324babd7fb52b0ee2bd589b529f9e70114f5fd6fe2fc0f6d46db350ac402e7a19800f3d60c7e94371169d6ef69564bd8d0c604ba47c1a9cd0755963f06a4b29fbd5577453d1bc86920c5c34e1725c8aec4cdfdb340449935f345a6f55032c08b35be18e186105abb106974cd3c9fdf2e7ea024ca7fd52911241d7153c29c9cac233b19b0ea0e64bc20f5bfdc262403fe79560726ac7d9c7013aa22d54e4eff6427af9f2b5333385bd161a5a74cfb93e1bc392d8ef0b2574de7ed24a71d242937abad75a774eed464e1826c45107af9d9bfaccf9f27128d259a173526207f29b6c76ed2e6d3ea8d01de3e7958ff1ac72c9a173eaa9809cbc7533ec87fafba6cdca1cb5886ae33da29a091500dcb3b976c514cfe13fece784cb6ab2d1418a1b9aeadd3500323e7db4e87f9159ed67174fe2160145d4161a98343fdd1e374ad8fee4dd3354b848ae01a2f9fd06763824c0b96dd546dc58a9fde70ea71885ed8007945f2121c749d70e49932a57764bdf759f82b9da4c79de20954957b467706dc1a988e53d8043188d6b3d43279eede434259ac52e621a4f960d9fdfb2c9076fed678722bc1c12e7cf8e6764996680dafebd8c9b10415c82dee17237bda94feeb410e3b52f3e2653a334d4ae307c3cfb5ce4697be7eb3b600c854368173a917fe1c739281d52e6767647bd5f95d4a5cccce35f7b5f989858c6a84ef9353eb35d46f372a370893d9b9349b4f674515b7d923943936b07e6589ffec7c1ee4bd11150c2109921020fc616d3401afa157097582b2263cef50407b730f714ad0e519ec325a3175cdb663db37aa9c2be206843f9326e85c2ceca6b02bb17e5ebe691681bdc1704ed3ff5499157bd6178a7af9f53459fa28bb3060a8438858830f82420978aa0a60be2f2a21783aa0eca662e421a9d4af8d80f0d58eaf3d7f09bff059b917c88020f55a5baef9d8de1724c687bb0e50b405d6ec22d51e63724b123a7911269c685d9442135452e2e66e071183edff7d4cb5923705977d46b1fdd58440100e3e304a42eb61847d131003446a3ee06d1c6c010ac7deeeb0bdcf03d64abca7ae3312caea3b6f536c60df76f227d6959b24bd75821ee0f3a2b990cc3ddddc0a054765f870f0e75fa834942828f649e1cc7b3d70e2a19fd61f7366f4db32f899fdcec278465937326c9eaaa0bfcf7cb6ca6060ac093b6ffbfe28a313ec3903b01f40d79b5ac61b9b1f3cf68ff4b55ee38e7855cb02329743be342f79a5f4ec18dac8767e0c593c93c74376b880a61c04b297e5c8dce024492985761c37ce9abd10d49989994316c83772bf6c40b233ce64c6dd26c132c6f1a5e57405b1a4136615364bd7d1304f8ed4242ba1a4b8f3f3140a7a848e554c861aba24f87960ad0a73ee64f5ca13a53025377651cbcb9754d30af70cbf20c7b3f85f8664bf2d0de01791c226642d7db6fc7978d8acfd2cb54f8482fb34c76f42acee9fc2e365ea543415b13bf991622274203315ee69e27b76fb872c00e40d96129a664ac3d15c8e86499ca29ec9fb58fc503dc98e2a24658907bd89df7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfe66d152e795656f87f7269892c7f9bb14300ffa7fe38b7c4c5342d2068abf0093a6b2ec3ce61439e4707379c8a7681b6db57c817b208faf2c7ff18c43a25bab194e890a1bff4a719db141a15f3bc6c3a1fba838d56e6a6063d8be2577d68a11857cd44496b8a333ded2b81b52b49424500e8a1ec4559a0f28dae101761dff7ecfb9ea11a126c4ea36b7d2630f70f4e3d6aa5fbc97b7e183db2391380889f5fd066fe1505ae74bcc78a9c5fb470a35240c9a5a1f5d9db57fac91601ecd07bc05db0fbaa584529c766b16a54eda931cb3f8d05523a782c657360c09663080e7ad4bdb5779771be6a7f2ba6bb5ddc52f22d160e5e5899d80b7fc75440439cfb985a64fc7a9cee79b234d816ace8066bbb75af16dbfb363648c9ee72b7099178769c661c36bf991c612926da691f75532cf1e9bd7d0c16cd6039ead653325e9a96e07457426ec3e5e5a612434c9f78b0668dd7af93ec454414aae2ba8641a3fa596003c9960d68dfe2cfd88f39e5103c8e530524b354f7138b6a451013601e71a1c213159aa1bb914c21ef1cf76efead8dd3f59925e41441a99f1d5ee4063a56fd8d5ff19cbfc8e75665cc3e1af7f12d0c19a69f8743ff72e44fa839855e76bcb961275ef4b7c3a826af158a9a6b8e680975a1a1c489b5b2defffe3c2ddec5b7634a3da3787d7b64d4f3049dd6210afd0b6d1014c6c13debeaeda4f2cdbffd0d30c4fc412e338203d1e0548ab93fe5216d2dc282fc81b005d1f0e159fd1c6ac063805d3b0a575e5b230df811339914286798495d3868f75af1cf5fdf17b6e0fc13bca14be07eff0cd9cb33396132d9ab215a2f46476527cf311dffc7969a98ea6f55c5bf124885eb687f5f71370f9641547db500ec66a1240eb92969de98b6519f3ef90b5f3b0ff23a58f1cfcabb10c61da8d174648ec468f6b2c11b1589c86ac07d76fa5150a0b8e42c9d60f6c7177c0eba420ced6be1a8e8caa07cb025c156e06da5b7bae9963182fab5361da7ed875b2f66de0004ab0d8a260d649a2a43c5c2c1eeacf3c08c7805e832054b00c6a969714f6c4d398178822a7db1a1e1c81a6e2d7421a4cb92340d49672250effb3a0da58fcc2ea38266b685690da23154085e1cf0efc7cb2e4efc0a9edee5c91d2adecd7fd5f4df8a884c6b0f6ea39a72e8a85d433562d2afa090f04fb968f94ce5e360f5315f96d7986612cb2a23b186a1c2af33be73340f6311ac664eec2162f629161b0864c324d18d7626183f680d01d7bd4ac85cb7dcb3a8c6a93300344d5370805cbf126cb24af212093625232019818802ad4ab9caf22fc5ef0e2c1478cf20ac59f5e4dec5e160b20416846f4581dc7b4161d8c8c092d3decf702a27113b7a708303d0b5690ae26eb18c019c66882d7c7ebd9c759b7b9e39a980d419fd7caae1964a104393eeaef72fd06677b15e5fca5f2d19bff82d3a3a3ba4ceff254344a622e20989dc2bff0f4b60bd87328f43567d78264ff3a804ba7cc54385db9976379908ae58126107ceaaf223592104a189b185a308cf220ec31cd7fb711c5fb48b1625aee0cd0c5d0394f510bb1a25f1bcf8f35344aa250fa4201da27e41aefae1f78ea46069a9089ae36007cc7332f3b9c503681db647cf2ebb423ce45f7c0c160fd23781aff53b2f28a1ab911b6108ae021d7ceafbe9522a15627112c663efdf3361ae785f24dd7df8e0d76ce2f52aeba84b0c5863c77fa673dea8e934a03eb33d380360f0cb749c7f20e8808014441c468371dad1ed8399690fa2211fabbab20fd646b707f8332b6a9a1b11d22b67bc2284437a2c752136d8f0cb6bf944d71;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h391e8454f8ef78e6e7afc3e5879dffc5db806721e8288c4426a122f2db6b8b8ae4ff68975bfd0b2daea0caa15008d16c82da62d71695982ed8a9cab1c2ab099e912e65a17a6552cd728cfbdfe9e8731ec3cfb463aa2b3b68ed44c49713c511214546d264a274d795f149151b01353d7b4293424d8e98ba37b44aab3fadc86fc4aa6847d66626596223601470c130c4380ad3383e75cf3c600e61fa30e6076f26cc960a94e2c478d8795f471bf4c453fcb140f269cd5c0291a88267ee5a60c1108d2a78c325556c56a8f82d289413f66c51c74fad5918ce3148189911884319d0b07204c2c3935d6646d99d2370b575539b3fca4740080b47ab99a1ff2f5f9599365243731c01d33893b4119f4380b99cc31475fba2ca4007feaebbbaf318b0e6685cbac3a40e4064a82189b4d80827eee995ba879808efbb8ece7b47bf6fe4147b9a54044473dfc846507890591f31982c18e537d90d1dd4fb00874bbe654ff87c173688d4a204f685ade5ba065f0c084e0c3c05962ec3006e18cbe36822433e1957dbc8ec38960c5c9fdce2a60d3f7c07836dccf65d7c7ef2264eb0daa5665fa9675b85c21297b06fbadbf93c3553846983afce863631a31a0a828168230b9cdbeaad481350ecc2f0efabafa83da9413d8351a77caf5e4c28009f026314076e4981f84eae58d030542119efdfa9895073797c1bc0944cb1cfaeec9bd3e46bd449131ae6e9d6ecfb4d730b18751b8babba9470f363e37669e8b02150152f40fb446085a27aa2d1b146ab4fa2e798334daa0df33f2c1a94557e66dc123374a4bffa8e936bdf19b4ccc85a000a74222ae79371b852788ef528702ab61bff3fb81a94aca740d8a6cc79736ba0e1dfc4bf9038ba81b88a3b930a7c610930ef6c5f34fecda06c760e1ade6870b0cde986c08d40098c23341d1afbdbf9b8ed235cc3690acbebc097c7f42d117efb9f1e1469b68221254ec982768ea201a9fd900a1aa06a5391b11b59011b49ca9573decfa36731f3068e90816354791ac461610c3c6a3cde1e0b4525a571b87074a246be61abc11029b05eb64b6cdd1367ed6e40b806dfa6dd5a9fe0173d26854825ef870c426d7866206a3bf405effde1528703f4adc822df5772bd75705b32eac25c7b98724fcf3f8dd5d762375996c162e4c2a1a518cfd6119fbad9564f66dad27577fe438782010d35ca8a003504eee9cb554306ae3da5858c10027315cc34831467da30b6f79ed95e4667e4e51d6d77c1504b4a41b8b1601213a46c9b5827d9b69a27a123834b18f1f1b1bd7c21fadb53b54af2917eff0ed575a83ce3c6eadc9b2b1cc7226c6876d0570eaa06dca4aa971fc7b434a589bd931fb6c6e3905a3565a1e072c48bef5f0e2f40462b93f60977e2274f9a587b0a201534843fecef2d1cfdab3db292a26d39642e51c3c063d9877437564fe2d9e8a83b77b7ceb6a1dfd08048004000553f5c6c96d9cc9c0d49a70af2da0010b1bdb0fc3705f64d4a80498eb6c0eb98dd74e957a63b3aed473bbe13cd277e46ebec5ba04ace7a2b6db53abc98169ec5aa5113a40d9e9b958f68ad7ba79beef9febc74679941bdd7c100b663da9e16f14867034e8bf8c4e6a712d812e9b89077a2a4d51b3eb4a52012329bf0d1f5a2520d0c8f08cebca7cf791b9d375cecc38edc07e618ea913f4f4c78006d67f6844c68550fe24e409e7bbfad5e439c5e7ad4b5462de03b0bbb20e396369de4dcd001d12bda82c769df35f9bd305eb6340a43bb959c5cd0691aceb587d340a65ac6a3690a37dc4b93373f94dfd4a9a04067cce4ba4c8ce8625fea5568de8ee72c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb971d27a6398d287808b51d48ddf37076ac196ff3fccff9176ab7f1c51212f6081a4f2e648788989202777e9810893ad15c0d38a8861ede71eb49b70243b61fde3cdae4b64b2c9135f180b39c216de327654e5ccfe8fce14400c4ed3b0ea24f54b872013bc5de66e05899721e52d55ae15a80d7bdee026e74f61002a37e9d4d26c6fa601936417f963ee6af8283dcc15a928a43b1656c20bc002d609cc4883dae026692699d94078cf175dfd2d9b5815859ea1660224847cec152829eb4ff9d09fcf0a976103e15856ca16edf6081c317acf2c943e862cde54d61ec7e11aaa11304d2c9b4407bdfd08e7f280fede0362a123b5b1d4ec8a3a55dbdceca267d1a349542acd9eb7bd081fd272480ca4d5831651579b05ebdc6eed5d9428431da016b1bf486a15078381a55dc987580ea13e5543662b5657e76bb4ab5e902821ade41ab8dadd8fc91eb2ae6339687d19166d1fadf7d90dad0e14a68277c8c5574bfa9b2b714e1dff88600bba8aef2b225cfe9aaab28e5ee6bd5e11d11c9ca57ed281b0c722e939fc09e4565a8affa9dc97400229d328ea8e2645ea2108233a077a88c0a5d96ea64db31b6f9323e829c91cff0f192d29ad747a2e469b7972f5b9d24b372c0681e82b860b15e191c96c35752011c215f6ee617dc1c79db3de7363e7cfc53e47ec443d999f9b36db829769bb0610ba337d270e73a18631937f4d9d2ac7f5e6dba668e5888db008663fb6a05dace79f31672d6b05d5a8f521d54dda635e04a01132a77dd12e5a0094f2f14404f46fa17c991a467e1318f403e5f2d2a1ee691ab65f492a19d1ecca7c63ed086831509f575886225458c01367150069d5da4e1fab407e03c91ce05be6df39404f946ec2b37f0271c6f6e52ca077a5ca6833a67dc60e825afd444871894a2b9d7ed5789498c6275dbe480585cd983f461e88c3e711db5403e6e486e490ae0222878d936f19a7c5b1af5ea2a22937556020836917c68ef2b6c7f4bd45168c844266203e6cac891c29bee9eb6a18592fb8e967891fbfa99b7fdfba28519eae1c7c508e26db70236faccd3f0762e002f945a6479848420cf9ea400bf19bd0619d04fb7ecedda2a444a98dd521aad3cfecfa0a08c141587be40eb3b81885aa14367b98fd40a29d1b678b8ca41a4bfcf5b6eee06fe561809c2271fa5cdadd26cd9620cfb12910fac739f046f9f8e21af93c3fb908ea6e28ae860c24b7e80f846fad751e89e8ad85d4a53cce4fc717266a23a00c35d3c8c7dd5cd743d3d752c04668b9da54ed08cedc28fe0eea8417aae0ca958b7a42a181e4af8f406c118d1bb298d412dca0503bfe09d8328a8fd1b8bf98fbdeb5b42b426d5eb9e3f8b0ffb7baed906c0f8e429a6a79ab8644ea7e3b53f5f298e47fb37c6eec57be68e6863c8e34963a1e53cbb40c921351d9e3e15b700c47bea1770beb7b52fa29a0afdea6de88fd522b1c4942e188d8a6f510448756b8b362ac7ebb4e932f802b3cb41f69ce069dd9829e858759a83515d94f7bda7e939ca3c8b3b4e6e31c32e36289412b9ff31933e933e6261dba38b18ffe5a5b6371c97267d406aa30407764108e508a555d10f6d25c510b8ce796b1c0bcd035c75a96e4ebf43a671a0bbe5db671d3d08097f0be87476461935a6b1685d067b27b408d0a3919ad99dc7f397f841ca5f304191cb4d7ec67a06f8d74ed6c6d27e33d4108afad15febaef62c27855d6a644bb698e6e3a69536956b87760d30ba79bef56f31b5d22cfa9dd0ba0e58a4895b5a6cd3c5861bf898a44e38f8c111d2483b42d4e58b6f79a68c9c5b5de989293839dea6d2726;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hff179e7056d59622eea35dc21e3b7b552e31eed3f8da3296445570e840991356a0490c43fa48bc9af0eb039f72e4351a320c161f8358b5efe057ae04ace4d0857a02362453bf93bd75ab9819a7ace9ddbb24ec2b08b59cf8085937b99f2e37001c17778fdedfff99a8750631d02e855b8c541594b955b3cbcc8d694a028a04f8aedf7b24d77c7e0ac9a1c02c2473c096bfdffa6efe0857df812a149bd1a50b0721d838a7ef8c729b885273426d541be0d9722d845366f3bd6fe60dbd62f8d5a8a6be4e183814e04acae308fdeab1469947629f2da2da45b2a0c5acba3c717a2630ccaab2580d110f6cda510fde9aee4e18febe88a36666a28ce9b8634b2cd4ac2ac2d13655edb09f2ce47edb0a14514ef395058071ca50b611466734975e93d59684d7ebdcb1429b24ccbe46d13a2a482ce3aa8bc17dba75d483ae895f0c767d976b14c2e79deac61a938770911316affbe011383a046a025d103a74b3d16af6239c442e06ae4dabbc93b54af46a150f25a76f89563503dec424b030169741994e3c32e162db6745e07563f1c672a1cd9a054a594ea0dfe7b9dd7ca376642e1a4f7796812727acb61964c8c655bd4d9d5b821da1a3bad80fcd57f6fef41399054a57e45345bf4d5a459b2fa746f958089a4f08049d7a614cc7b46863b0c098b2f8d8974384f7ff3b70336c243906480e0ed6ec8305250e3108d8499c3da67d23bd11cd0771689031d6bd2176bfde461f286f8cda3a90bc9aca80092f1fdec5e2ec9672fc8a14830d66b31dd5629a3a10ba3c76314bdddca2e16f596bee678d5d1f76eaa726171b884c991ec21eeb9d95d8272a72d70643ef664132bd3570611f80d075c3cbf70552ad119a383b48740dc32dd962543ae03afcdc7242c86cb4fdc02c9a5e373fd52512377f749a1ac68c3c3c4ed270c40fdba85d798e649df2227f3ed0de16cf74f09bd8987dda084d467ce014cd4ba137e2b7d9817849750b35962b82847d9e66a780356e9eccfd18812becdc5f6ea98fe1645c241c27e15388c9f1f5248fd3318c015e3334a3ae7dba2904ba6657f8175d8a07e3c805e7f52892eb27a22fea986690767a7fcc7ca1d68f5f1113e8aca86b3d78c450e27586c41c4a393208759ac8d76531def1b0e89b2d356409c7da7e3efb24fcdbd3f632d00a6343358089704de80ed298e63a2f462a7c44ec0ef93593f9be2077e106d95456d8a5c3178786786d06ff9f98b6481f35325ddda64f9ca77f8d09378b7c83985a4f8ecbf0f4b6e686c79fec7e9c4f06ef915a98b30f29578b87fc09303d70ced5bb5b711580b55adeb71690d2164b6e9d2d878760d0cbde5afe5050e8a9bf12b22219acabcf12857c6d2f87fd8dd23b85bbd1cc2814c9bcf3b51142866a1da5e0e3ca42f8f6ab3ef6463a07c669556bb5a90d8e2419176281ed66b820ba63df236a857669710344550633b5ccded65c985b245177a4ef70a6f088b17cacc2b98eb98c0336e7395f440179931db78d83834ee7cca326046f18a6e1c002598bd81e1a2614bca596bf266b59a9302cdea7d234c1aadc7d18fd661915038cf5e07d92f167106cf7e5cd33bb599c62e1c35695c1d705911ccaead74b763712d338da9f51706e0c8b7ff6908e993c532cc902d2d3175d4bd80f70b051ebc10ab75c0671403ec141d07321a8b629260e9baed64ab2a78d328b3a96ea56eb215a4bdae413cdfab655e3d2c8f9baef03d66abdb4db9f49f69e7c0fe9830da26c0874c6a35a74534b64d83f2c235109230b4fa49362120180825e0ae46769dcca40e8678126714811f8a1298d5af6da46eb76b039;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h5c147428a7e4c10e0e511267daeb33286e0bbe1eed1e45dc577fb02ad1ffbc5f8ae6c070cc4207cc22b7e371850686e6e89741b8942c9af95585c18c835189320caef9fc33718f59c57faacf1c1e65ec4cb79a19646b608890d29e19b7d396364f9fbb2a13cecaa638bcf8ab850eee250c8e0257aaca031af5db50d8953efcaa30f135a0e5d2358d09ccf5cda8f9f5a7441ed376c9a067d5cddf102572a4ba54350cff98b098f45b6cc2192c4a4ee5ef0be726dc1f154d8f0390b91d522884d26312ef399a99a6baa72e614c996ec0f57b73db91ff5d7064c07a5f83e39637ceb775dac2bde8643ce3efacb3a3c534459a35b71cd19c187a3a012fbb7c7d16de2f93eeb7ba0455f1d28476d0cb1029efd6d94114f3a9b4047f2eaa0ccbb09dd99fa4d0aa5beb15ed1aaae430a493cdb5d91f5c9a2052583b4b832620c8540d7a05b4809420742266b6f47ba6730cec10c5fff2b0fd0b273e49ebfc75638e398c80bfea316e0000432d1770315f98585a60a44893f4a3ab3cc85a50b0da7dbffdd425a881d5bdc4e8d43e5ead54276d4dcf08b16cf9a0946274f1f99286e616c6153bac5503ed4155a610997c86bba016f5bd4e60d7c1b24282c4765a3204378c43955cdf98f4c05305b61617c5da47251174e60262c0538ca9e905dcd640b1e4c1a67f7f72a16885fbde5d00cc064be87f1b38626ecbe49d6dfb9abaa4d12ba875d4a02f9e1e5eec596609ee4c916f8004e73d79a9bff8b1a286f2c233e69d4c07813a0ecdd111303b2f28c0932264bf70b3852c218662f926231361b9f30f34ca6b2d51346a5d6edfde6eba31f5d491cec7a7c772420bf56d3cec48f4a21a69feb5fc21e9507cf08cdfad7f61b9f4ecb32a526407e09b8d8d1b005f6cf967496f1b5a9a30de7dce343a6648eb44897a38f1287e48319c112cd92b95d4403acd1268d5632474ebc59c23470d6aeff04e0236c6b0b35bf40589268f502552065537e806fe07eefc3833b0537ef0e79e0d078c93e4c0606bf1d04732873c01ab3ca334dd8fe0aa5d46974c8ce2b506788800e8e03b240650d0bef0ab60ad379a26e295f62f9865338cd6b0df6e8b6d12a3b6e70412ed61c71ab1deccf49c4d0ef6bf8c0bc3febcc58adbcb9edf7e51945469bf43eb0fcdbf64292734f6d22fc22b735e43e3e23705804c50ea014717cc41760edcf2512ad5c115b7b82b76d6a7f48df334fd335211b69147a6bf898dc1436d79d8591e800cc1132c81e5a4da26cd278a1407a4e156c6f505262d1200d3a1fd9888607d2fe921cb2ba142aca58b6f8bc4a7d16025a6d78f8a241a33052ab7339475aef1fe0c6bd87f9803fd508c5ec453c13983daa37096e64e9b8bfcd05a1be99316ed6a3801f170a207a5a8d39f03fcdb390c4c8df1bbaa57babf32fdbc527973f0cd5754f383e8557ea8a7d4f0e2af7d72d081745d40b2e1a812a72e835ee2f350a12ba0c8eabf20efc3035774dc958d61147cc0c14b175d473fefa42560dd8ad62219c5becac4156680c3024ba3cf0a31895e1e07c7cc2e288d1b1e3a8264a3e6708167fa77ebec539d863fd0bcee82b1cbe42f8f9df4c7c3a8988fd94b210a1f9114c3729d36e31350147311687a8d2c9a12138e18340dacf39918c9ad19e3af450f7bc3def46903a1edb9343f26bc9129d9457a0d7c8a596b444391a799127afc9dccb18fd6de979b8a7560a9afa89d0629ace7ca3d5a2c5cebc532ec9ff752615cb2c71fdb3cf30dbe9d35eec079f5ec1ea674b0965ff8d4dd92b3bf5cc3b4340e3b9cc7f64d5a7c63ed689c64b8bf1bcc77bc9ef85810e743b182;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1caba1761db077719423c7731e5e897a1cb6403dcf3bd3820910b305d61dba49be0d895f41d2c1047bd72b33efadb8b8ce31f386b7ea3e3981abd8c40dd257398881f124c165ab8b154264ca3621c7eb1bee29be922235559f30daa85bd01ead4e2e5d9b1940ddc3728dd9b8509570d7c7bfc0cf755bf7bf13a7b4590b18d446d272850e76390c8b63d5a0c5a6b2b486825e3382acc7feaca30a69ee34445e7e7fcc6b386ee1d5ec0c632f196bc89ddeda27cbd74bd940599739400da9eec58c8b9ef03dfe77666bb68660614e8727b30f8cced3b8a690113226cd9019dbbc3cd3dbc41bda9bc462e4fd6ee68b9ce93d091c294689b5f0cc63a018b728c79a4017ebcaa8478f1fa672b2679ce6f482f5141377c285f141a2ed62a97db7be0debd396e01913f3a68e8da9f7c272f4d0eccf663dd0b1fe4bc17bbae404309d33d7c505a955d84ceaa4a9099c43739ada9901622fbb9d088ac3b880c03a17eb0c868aeb027d2af3f8d3207c208e5a066406396ddc8f0d4ef5eb6f8dfe6dcd0ec01142a6c66993e64a23b38b7d40c8c6562446a9d248e7f8bb83ca6d0397c14381f13975d204d62af4ed7ddbdb0b75315f088377e2a0b990f285725afd9cab5169e18fc188e831aae2d51c4ce28d4cd948f3a88273ba7ebc4e751e844181379259d584cc50419d19941d050580e60ea4a221d387ea6f4fa78d9c319a5284337d0b6e19e952513273bf58302a725abf7d98bee9c2b5a3b424ae6af0e46bd38a2fc8c1c7fd22946ca48afe576dfe8bb2975d873d9a22b4bdfcf4c825cb4cf9d959990c4ca013727dc85542a5ac614c857ae591a588b3a7c6ea2c3203a03bd08145d53135b2800e81b116747d245af2653ae7aa04ebfd187237cd224a101c4eaf26b41b7f9fc7e020c8e2c5f647b266a9b08902a3f43b506668732b91a7bb2309b12c9764fbd2704b774e0294a1941b62f419955594d904096e3874572e299e93985bb823704d9f3dd5a19806ce35435943bb378f642162f59eec456c7e0aa9f7b7e136b8c2084dc167d171a4d86b0f5c6887957e11f9a41806468b864459a3f899159bf125cb3ae0f6ff2e712433731675f31c34faa5b7d2d9f1efed9c35b55699add93bb9881186192481bf0ff52add54ab2ac6b775533e5a79c6878f97f5346577972dfc84e39da78cf956da2cc49ca22b3e6e4dfc3a981dab7ede1625f8be771cc8d5a8f5bc5bea463f00ffa58e3f6a8a48c7c92ce2be83ed23970a610a8219324a82c9b30f9d4e295fe4edcec044334e933b41ef564d9a7567ec90d605a360580ceb07b3c2bc10488fc69a74dd85789a65a3aa02feb3e2f2e59f9a296239826ac46e2603bb487290b72428fa1a8c57e0c35149cf5fed27bf111a501900ec3aedf7e1f4476e7d3661f2edf20129bbf63b31e1f6f1f1208156317a09f7ef8012b89f2280e3399e267170bf1f9bc011945b33c49c7ad1db8042c00dce2a3421ca34091a1b53f55e404caf932f5a63858c76d10c3a3e6cd00f603895df1fb91901aed5716f327559c65a07118db747bcd2f0ee503aece7342a38e244543568f05b7605176e34e876cd37d03019ebf6509b4d56e602c15a3e66b8bbc144d70c77532ce9f11ef8b981c28ba32ff313bc540ebdcf6a3304a9dfed02f5fe2ee96ed47016a41e82b6391667644ba9dcb121bbd99ae65eaa602d2f99836220e8e2d58707eac69a05b1f5efcc9bce6485b5378cdd503a40cebe0a7b18c79284457921b4c576f18ac8805e91c2bc79affdae0beb3a29476438c2753460f12945bc30c86ce67d1c03973e6cea5fba4cb80a4f81632933fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb131c17f4cade5cbacf8c4023d89c467c1032598c70b109eff97c85975aabce6b77da2e0ed45e087979e44d1a3a52b5d2c273ae1850aaf715b9f98b406f9a6ba043405b16ba0faae4f828e24e2caaf12a9002507f3b7ee2b387f61dfcea965caf10daf28170cafae058c2d44cdd12d1750c5d3ce96b933cad0251a939890943235247cf394fb5290a8f023294430170406c1912ecdad9d1c7d89169068e105734a3b3023a9c2debbba948af128930cdbae05f84f598a5ea2130a751b6090026ea4d376e87ed2c300575b65c28fcd25478fb6c79285b0b787036af64c1fc259acb4b381d7b7defc756b5f7f82490c38e661b68c156bf1b55b19a566e0c846eb4d58d99eec69ae3f19adb18d03c11c6be90b37b5790c27ff991a9d21b8e68fc9c17543b4864d3feee2b0f78f57d493dbe275eda8cd0c9b302262e3f0b96e7e7241a7cbdd20c3bda7c9bc4af460422fc9a1450d5ec9eb7faab407577e60cd97b62fe9e8962e104f1d6d02afe99b1d89c3456902829e42480065e6036af5bd61375fa195ead8990789535ae3c37c58c681c3d1111879f1def55aa5ff4266295decae0dfb65e975c6106e5b26592641356118c01ac1b4f4792279f046abd1327f012717f41955e97a7e34e9739587eb2c7ed552762fd783a1c16869cdb5c65e4e14b0acac9da5ab57901b055e9ae28c7223457cfa59d63eec44fb7fa72fa9046da0862e7bf29ad22ac8a15088ee958a6d4ae7ed08a7056217704922a9b43aca801c965c8221c7c30516ba803173e31434f426ab12381ed87352ff2e9d2bc4056e26912f3a6f8e5ae8a21612b50d629def978b3bf257d772542ae7cba064e972106522dde750058452b5995ba817acb56a27b3a769484ded040a386ae693371cb1734928dac42ba1af6417028f6a9f161672f10b805d402a3e7ae7f0d3623d26557868a20a896d64475d8722e62065d3510a33748642c61255161307b7b873cf88065e5129697d8ba204a9744157d00b7fe395c4ecf428457041b7884adb863164c3225bd0c8ebc313b4ae8e21de3cc95346a05546290e73d6dabee749810c8a48af9d5b6e1b937e5bee5c3cef246a65cf17db850fdfda1bd704306d2351f6b33bf170f55eac63e28ad462c1edfc82941b528a6c13e8010d59dc7a9a2555f9132901c95e9ce012e6ee8277407dcb97e9907d51a2703aa541abdfd0ff3b46894d9b553c09df09b335ebe494d05b8d7003c63bcad2ab715718c6f39c563756adc0a32f7ccd7aae1cf1c618af77169cb65bb0e3f4b5fad0dfeb54afea7d5e3110452c6824346ba80559b877685879cacc31c7858c032203d856d0da975b89f9b52c1b9af65bdd906d1be2e0dd66350784fcdf84712b95a32745f09dc5894332e172bf4afb4e45db05588133ad49dd45f347f0f29649c74047ac686981577d62005798f70ea259e566cce9d5d563f9886a811f021ec3f2c81570715baee6f9219e640fcfa8985e520dbe6306fc0178c44db99f2b2791940b90f3a3026439c419178da3322e6b75c664e10a06869a43526c8dcff73d9f7b2d9f943035953c0937b4f3f05b6cc085d44cdbed3db65c2cda5320db501af9f64905b5a78dbcee9934d4cbb8ec0050f239d99f3bcbec93c4d752347b2766b0e4dbd26df6bb0ed6fb405b6d02960f0a09be04e8252e9a4da4deba0c884727abe4877fd85c38219f35bd2106b399d5146db9bbfd0c39bfff96025962629df76ec0a3e138f86a317895bffcf2ce191db39fd5671df3dc13c727c906fffb67d33f5a36384d70646fccda44ca2d18811da5f3fe2145cc6958be7760668434c1e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1200a0ab35b04a0ce381654a74d9ff282c9d863d05fa801a0b583be4390c438230e4e34ced2fee6600821eb442ad4dec456f333a5d1386910ef48a3ba9ee764dad80bee14f52117a25cb4db4e2221e4664fd0dc6a7a752d6b7ce682a96481bfb6e50028c62b47ad04eed02a4c2e709ab13a4458a432b6acafff89b46405a9cb2e1e36471b5ae4a0182d6ed8c3a87f1f16afaccdebdf8ea6ce85270b0fd0e50226ab8c46cc3987f23152bdf1661bad6a3aba812ce6f7f9512952479948fe55b021993307645e2ae55c28c2966a8e121c10b0b7c040a6dcc8858e61c5f8248507446d19e73b7a00e499d783b7454de11309269b9a206d16060eaad31de039cb9e0e096d26dc21c05dd56bf9d9b3651fd1391fd9ba45e4232dc6618476c9230a0a6251ef83f644c20df0ec870cc79e2c3c16cacf92a7ea6f3ba8f2096150c35fd226ba7ffeaf53f7f39ceef51b58a184be296c0760ed4210005d24e36b04e49bc7ff229b7c5b13fda73a0336823b5d8b7f2ef5b7a781d34122895628690c9be836d21495e5c864cca07d84bfeab8e2ecbae5fc2cc1707e6f284eb92c34bf321e132bb652a18bfc1a83ef1dd5b429de546cb772a09823a50e45e6f7888cd14a592045c3e56d34078fbf122fc87e7316e39696ee67fd459568904bacc3a37df574600f3881e3fc0cb81a647fc556ffc2735fb53d28a3ac56f5f2863ee1674e094188a0805a3eb11d066624ffda39609e0d1a28dd7076814f62a3b28428b7f40e2adc16430b2dadabef8415a0728f32445c81cc0f941513160de1f5e6c175314fd21c06a55f9af67eae8ddd135eeb9ff2f91c8db0f82d8c331a35346ef6d43039f6ec0c0fd232fdf62fb2bd290b6efb9282536f9aec5724ef394be6f1ccf3d62a4ad8479a92d6d85fa7817994439088690dda3085ea904a074463b5a71564bab8b872f9ceecd7b63e248c42521b3a122afa7e3a519a0ce4d03b1bf20a0bb945fcf25653dc70c199acda0658b89f7d45b4db4c4df026d892ba22199246ba687e040364faca078b88f6ef7a489746ac8946c4f8652089997cdfe07c9706db4d9f719dfcb0b03c6e2f5eba5b0cc04028ba6a5de5f4eec9ce9bc401d70657ab043da5056726608c8ee7e4c43e9425c2a0f29cb82aab43d8d4e13023a2c3629ed4cbce3f6619bf36f69db6ce8aa667dbcaa6b09e61d5eb68cb606a884acac118373db9f7308f769334ad6445a27e286d2a28a6a649037b6daf5deb4cba14445e532c585bd89946eb9aefeabf337001907bd3bb43f5dcaafa3ccb5a21a82f2a567fef3da5efe12430a3f36bc965f67262275490dfc33caa669ea82602fbd65a00bde38ffdbd6c48945a59274b5cc8e47989e0060b27eaf3417670f930f221ddc8e6ae37456c4ef63409fccf5b5815a8b71d422d68988cc95ff0a31124ae2a529daebd213553c52264e05142121058234462f3249dfd4d738073f199041bb56603359770d2642bc9215a6c318444d989e2a8f5fb69c8204864eba98a47dbfb6985d1b5827b830148e1ee8d452045dcdf11785755bf132cb84a4beef60163a1f1d7f84a20429b5a870145a9ed17c6dc918dbfe67bed171ef6c57b2e0716b897ae2afbb3885c5510c2b3b4472cfd74f4873e0bf220dcebdd1f65f28c0cf03fffe46dd48eacfe043c75cb8df62c9b65fcf2c197c65172802d310576fce64217e172d7b45c44770ef94e6648c975f9950a529afda3f58db708eced5527efcf4d45b24fda0d8fd540ddd8f08dce6a2647851a4b350e877fcf048edfa32c775e220eaca1c21124efa95cd35576405d5c706f5302d0cd731235a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd08280bf758c08114448f443facaa99757d4f1c837233d8ce89281639bcc42c3074707ca82b62b6a85092d905644e7497f319d00d66c9a75090f837ff312fc9190f6b86072083a7b0306b27d599b2e6afa2f3e6bc3b0768558634233fe4e77627a6fc2880aec54dec6de1c64bf41ea74f3b41907ffa4abf38492061beb6c2a7dc523643af439359cfefd5956db06a45748a00a4679cb6b1c58a4ec7831d117409156bd24c29e52382311ffddeed9d1c68cd1572540ba39d1853947e69b109dec04bb5efddddaab7a2d7b184a8227cac48c80844f2c3e7270d4ebb1d5274f9ba061476f6db585e1f9c76a2ffa0d7ed6ed611c460b49d7df995656bf75f581521bd3b7c5636452f1a70ba74ff019784f385985f615480e420f92ae703c03c9008c210cdf842acb554d7428c82779c834844a59a30910270192ceddbd0b913f8369969015a51ca0e5bbbe98fa9ac8b33a196ead9096ebcc7d653fa5ef5bd36f7bce37119859743a3a993819bce81e5c2d8b9aa2a68681f7b028ee2376d6603de56bdb4f37d07539267b81389237b65635073be46ff763b8a6e5b1798ea09db4152f241cc520781f27fa19237b090531a1c6c837725b74567bbb11fbfdf3fbb53d01a75911af351d2ff671bcc92c644072f48cfa253286f2f8efe611b112526fb346799c9e2438ccce1c3672b65da9bf8017a9965571ab44d2d87ce6ff4549fe44109b4056e038340c0a5a77deb91c6dbacd1b22eeb69d7bca7ce9469719e9ff009991687744d388cb1df7534fb7c55b809ed7def37c605d25d62d493847dd1af0b0ea88b685e57124a74d51834abe0084960362c5e163fab884bab8556c605df4a32db67db4460020ed108bdc935823d23a7ddc72873057089a9882d42b408de8027399fcd0e24b253db04650dfb678a56650165a09121061393736698cb782554350458cfe55d370d22a4e15ed74d3d657a2a32c36a60f031b7c3d259780978aeb0064081eb00b05bfb443f46d83c8b75dfb90fc9dd01a92a44e2f1cd7f4c81a5834c473dd37627fe6c9e0c3954bd74ffa6f5216149a946524e7beba3f4ed7b42fa9ffebd3f254efe129080e2f29593a9325b0b71c8dccdbedb0ffd556097cae2e5b34ad3091047053f0b6ad32c4266449b8487d61098df944dd462a91a2eb55f94fe3674e7ca2bae407f54ed112ca5787b11cfa2d7b0ef60d50cfecbe89b6269fe15cd1e49cba147694611b4bce576053a8f93c49ee4c4f5afd9d939ff338116915b21e0467996875fb928656e2267df552e0a18a1088e984c626c754f58607e031e543d7c7bd9cedd28c8339d3771e2e21eb4e2820196a823b51504e094b314d1a9b871e0e84b731308f99160a01603e2a603b7881bb4215829904783505c388daae739c995ac956d7b55f20a18aa476baef92d92f7c7b3adeb116c9992ee36a0a1092e40b0f0eaa0119b05675fc40eaf0fd63684d1f27703d5fa2334892aad35ae86485b3ef841b80258ea0416db2fb4814debcb375f60a62704a9dab2266f34f555c89d3320bc40da3b2620bbe71913a3b2db8d9181e84e65f1e4dddda879010853ecfcf91b570c6603814240f2cbcd35ca601ba17edb62f8f05e9ff98f3c6d90f22dec572a96e88d8e1a3e9114e75763edc2315648c468368c018d4ae4baad565039ceed8fb8b3165975eefbbf871e5ff02cac65d56a0425e697a46ef9be9c3050c0fc062b83ebf8fb9e84f23fd96a087870f43b78eb7923b794ea72562cea9f3cdc9ef069236602a28e565ddcaecff2dd5dfc68a2fdc43955a7a327bf8b14918ca275d2605a1ccccf2bdbb30817e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h22a9eaf5e3a01db21bab1b8267e4ecaa87109039a9efff3266d45e51d1dd0351c0a6dba60f6082606945ac62f7a2e1ff55afd9e4ee2c5ae06654b878fe69b5468cd3a5dd1ce7437a2077d2f7d6dabb7fb7c267c9cc63bb63c2066f4e5edc7a52bedb0799ffb1785662ca495898842d89bf2c7ad6661f8b0d57ad12d729a6d69121db3e8a1f5e96165868674bb98c4d9d9a15f64e43a496d285be8ce3cc7b9b10038dd43774dd1821b1531f8fe0fc9b7b42e4644832ea32339486bcc4780073d6ef69bde6d0bac6bff0d895879377b936eabbba128e00057ddbbf7602c51dcb3a1d89f67f604d5dd4d699920b35e9fa07636957177423176cba60aa1b53d27bd76b61cc09f9e0ad648af74f895de88f5f3de78f6283838c84e4b96556ca7788cbcc4e7630c14433192f4982688eb8f87b3ef529614b200e1f66d761b0bffb8f5a86dc031c1e0184e86d7d17bf2452db1a2769cb3af7253c89d658a8eb4cdc225ee20421534a6a0bf9bb46126b394eb184b7acd16fb6b95aae791e9119945de203d69cab474c8303e5fd6e2eca1f87d0409df284297069b7d99e1947ca47413f38de8ac61507b762e0b98e5b21dbb4dbffd0b48179010057aa34390889c5d22d4d7dc978a19fb8f3fad98ae5dbec8290b584c256ff1015cebaaa07853e47138fecf4a8bd8ab323b5a9f6699d58703d72da42f9e3a8c8be33404d11bc729c8d379d04bd087daa9b2ef82b30b51d8a13c4f78322faa8522d920d67d8c285008f2081e789872cebb001b19fb5c7eb96af2adc6fa001971534bd97d7689a12b0b11dffa2e54937ddf66f7bb86499458ef15f1766260df0665a920c6613324c3582158ff6e09f6b0f7ba5325d5dd1780b0eafeaffa41975fed945c24e05d11c78b93f09e8d2aca22ab593542e832eca0fd9230c3f0135720dfc48fb39f1b96edd1a6f1119c9a6995f284c2cac8db087a7bbb8025cb0b53afdef176ef94deadf18b0c1cebc1c614c2dfb1dc9fcaa6d23c3cd49cccbdcae2eee567a17ac5c938ecdb101f12ccf1ab773e75be0279805130aa636353aaea4e7865bc757e40065dacfba0c7d4f231658d38f91473b58e9567c94f0be2a75d028491aa8c7587930cb4f09bc74434531d14962bd0fac16a62b22cd4e8ef2e4e551a5afc34902f3e25ace200dac889f6090c90a1ea1a7f9c97c520bce816ed2387d9a27d65da53cac461a4104269c8c2818ccd87cbb256178a50ac7d9828b1efc16fb5dcd38afda5f0459b65055589a78e250b65e634cc5be7a36ff96ea35a88c3f45fbdc8cab8701e9558cc128d676317dd025dc0aa60f5336a106fd42c49987786c72e671a500fbb3f5102f2b89f5875570a7d61783b27642ef27bc97e2ca04b5bd41d0f907cf48cc6fe02407dab76d01b9a825d516608c406ef432d59f775b3e7ecafe0496ec8210494a5bbb8f9faf524af2334b6193b64b4f3da06c385580c60fae116a33c76c160f87d1cbfb50360cbd57dc0c0fa560faf3ee486ea017350c69abe5ab0ea1d6ecf5bba4962ec7075a897f6ecabf0ed825c082ddae69072e8a4a69e2bf794860a900206ffc93d7c75db477a990ae631f157a61545daa1aefb8c1cf0a720a3af5f1d967d71bc290fa12073b6332f959db07a13b4ca891634faa50b630c25811ffc975a2f6252d18349b56eaf50e058b68e28f58d620dd4c25da8e9327aecf7ecfeac612af0237723599950301589676ebacdae50ac1d03c8dcc63243447ad44e6efb299660808ad0cf7cf7a12353898cf7426499412e445dd62c7d297c2430ff89747b03721a95e98cf2c6d5c98cc11688aee7c3dce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfd4f9f7a3ec135732469566758f49ed9b94449d9f85b54d51ea6eb406b342760e97743ece2280e5a70811542347efa5bf1dc8f1dbaf7654291abe5a424f990d49ec6d709dd2931df09172439e6ef24b5a9d2aabe4b19b0c90b042535b5f509e43344def6877f9540291d5dfe54b43b0f84839dc10bf37fde879299d2e59b89e68a0feb901bc12fa860815073d71891c2a504d2e6390903dbb2c908686e685e325f4283ad8e1e4cbf42688eb81d97c4b01678bee661d14cc2146d5c22ca364d56cf65377eb629370a888a04712caa975f2c7450e790a1457f67a324917f1e324757758ae72ab091c2c8bc7a7ca50ee58146cd6a8a8056344cc50750c24d4afaa272e153343d7bca4c973d353ac5ef1bd9f14245485eec9e5b48f3a530da32a4012f371dd8d3454270b4ff2ae9b73f584ad1076a49b4f986fe53d87ea1c313e936d493b9108931749a3fc086eadc0cf9c950cc422cacd2b46ac52f0d95ba2e637a5cc56818a05fd1053769119de7310c26a7b56cf0bbb571bdd60b6268ac5ae88dbf06eb5e8d8faf2f1222c94a42e0ccca1a0e4056134d5b822516b14a74e09ab5cedc8e75afdb501730c2c7f5a10f700a34a5ac142eb209f7a5ff81c8bfb790654ab6bcb6d013c5f1a3401c121468fc0afc3e52c513bda4b3dbbc35c69abeaf6e652d6d14beaefe0c025899039f9b5dd8a5c218b0602a87666e8b572fd546ca9d4f95fb1f0dfea3d8fdae4e9349826d3a1ff423ddae3c556805564e1bcfc67cabc212fd0792da9e3e257c27071a6189c3648c157548487229d196b67ffa45acd0db05f61c9d786917540545c4229f52e2060185185c03e2fb6d02f96260537f9d21d721bfef2a05b9e5d510476e0907752a415478b423c4162ae5592382a8c0e627a737c0b0a3b984f535d7d0034979e4a33b657c1dfa30a99aa3ed88f620998c13af23c8fb4f79eb41c61dd78da2bbd1bce91c5c065249c4b333e366a0b214dd242fe0203cb636b38b5e2b42b23b6111a7e05cfb8c5636c3cd2d43ecdc0b0e0c79dbe86fbef094bf7997b843f3acdb7d9a6c82e316091e79f13bc75a9a2bd56b61eff21a271c2a3086660451c51de325c660cf427a22a52320e283d0347b7a595ae33ef431b65a2444a45ef80e771c490d57211b65eda9c7db7ff1737333bd6932aa293ee765a8605d226ce0a1be42e1a40b7fa4c41634bb45f6779b83730ac48ec14feeb8bdf52eb9ec029e863f598da8a81e65c26a84a1dac271c4649642a259f636a93bad6b4cf2d8fe14907a11d04198d819564c11df383ce5f7f87852bd0bf0df63ebdac19531f8787efbaf87f871093ed1844c81f1c81e5105738be4630b71f7b553b00aa749dbea68f14fdb134813a1590289676cf5cd8905da4a08b8723df5381bca8935c3efd607eea27fc038a80c2e30e1db82ee120400d217ce4956336b53d50c831cd516807bf6586e61d382474acdb97c67640f5c4947a0c693d6dfcff798ff492e3df3781a628b11e361a2abafcbdc89f2aae9e71215c32ce912bf50a5b18a227f6fceb83dcf3d1adc0646b07f17d74c14118bf089cc5772fb9a2c17a918db569b6c1aac01ce35903be7636c2897e13fd7745677a99e75914d8e6e7b2a813bd8fb8a1033d1a9d0df6c843fd3dbafe3ee8af5b31ded00f66b67193e97cb313b6ea912eb6546fae037a95b12a09eeb907e59e939549c33c62ff1a7939abcb7a1d18a9b44c73406be83a5285fe5f788616b7cd37ab293e50c49367a971b6dbaf6949d71a9a73d93c812a003b86e340fdd95a8700a0389d4f7a9e7d251905ed553d2a5205d2f4103f3de18;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc9d58a5dd609510b4dd903f8f66097a21d325d70e05b6789f0b12c3ed62392587bcc4ef24566e30f3f4deba95f338e749590abf7c3bc6acf0c9379d1c93cf9b223d0d007a69e1806760a07fe1acf6cc326bcd32eaa9afd433675572206875d57252c53978ced86665bf10557278d56b64116b319358b689a9aec94588c9eb82e5e0d949d1971b864d40879c85de374fd523c38e4230502546e9df96cc58d51d038356d8bde867755a2ece92b2e636048096e5350d73b40c5c724b3cbe777d8eac9915043008e5631545a1a8ad6fabf66ed76abf0afd19bb99efc4737edc09d3e30075eb815982f6a9e4f81512fcd4580e4abf255ceccdd39f5eeaf57c3ffa98744515231dc726507e2a8a55f49d842137683af5d5ab7802a6b4793398a52c8b5516dde03af0d4b0236ed4954e9e2e75f09e2dcc901dab359b532df6fd1cca0a862c1531def04eac70e1164f014af7f70d144f81f95fa7e03566d2f1aa672b3bc73097cb885e495f452e19327a8a485f61822e22496321124f897a4c49ffc9e34048357e7e37f6e6c1438fa34db294e3c9526838b1eac84c9881807608000619bb99ea96fc7dd6d99dea55df588974c85b9d138ffd4b53306fb43636ed25d0ab7218175c9799ef8f6ba7b3b9f105b5c4ef0ddb3df7d8aad3226965d58f1a5b60ac8f534b2798b6bae8d0a2f34377bf0c2374ab7461fd1bdeba9256b74dd7125b54ad0c6927493b8593d695ba955b215a8156849aaaf3952057ec04d703b932eea0065d5093bf8dd241a29616a9befa72eee35958408ee8904a737b5e0b5d442f830d6b0bed1868b9835d4f22b2a5745bee07b76f5fddbfa3d57845d743aa398c63aae8bc34fe19ce4e9b630b836af6a57d98e66dd242232143259774fd64776c9776d6721747fe78a9d57e6f64ef41e7c5f4a857044f79e1c102d4afbc6951741e7016eb1d7f5bead8a19e23dc3747f20106b3d6d614f604fcb8496a7c7f1a377a03eba169c3c209abb11cec02357768a11bc0fc7727f91a8669277f7f9d4e07c93c82b3c42541d48025581f4dacb72b3e4c7f5246b02032a276477aef9288445166e6fc1ed3ead88d995c70d9af93447cbbc4d64ecdc32a4f1d9073864bc20d1df764aa27d3f455055cc44fd4aa6a686225198bac2775329d2f13378877b70095aeb52470ef298cca3817a4c3ac9e262a57408fba95c259b873d3675c1fcd5d282106b119e7b419fcbfebbfda68670e0d45dacc102e36d5a664b1753b0c36f56649dfba92cf58a8eae6312bae60a1286d5923323751b690130168ac4acaab6813cd5b37f0b6c165e1693091925ff318d40e959de2787f425ed9f1a487237a7af98fc3a6f7a8350083607707fb54ea6138b91c5a519d31a906308bcad78ed3bf4e404a949038472be91c6ce65c34f36b869a7ee485940ac435205e831ca4c7f135aa8a4f42b57db45ca10102ba34d6a2a961c4b8fa2280623313a5678973f61501840e1bfe9b199bfa91a6e6924a53d215409ad50e19235bab86ed411794bbd897fca37bf9960b8483e9893af0384cb12ec6104a72fa0e843753ff5574550b194acf9c9d72dd709b946c0d1467d64e3d7e5be478d2b75f742b3f7cf8111b2957e090e2c18d50f5ddb24c73240e45ff5b10f5580b0f56bbb3236eddcfad45a4a8e53e77374fc10e0118db67c4289a842b086c7e3bc44e14b17bc75d1182290c661da79bd65005a01a15be2e4db5affe68c78b01e0a899ed61563c450fc938d788adb87fa49626a01c266b3d989d94f99fa3d46e85b46b6ba18ed89aff8dfbeacd12b891d74c973de9fb58634910516c5f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6f33871f29dcd04d29fc84c08c12db50f4ab1cefb4820f71f807f096e29d7d3e957803bca5d77a8f20c37cb932b40182c30ed2e5ec5070eca652134c391aacdf2a97290ff519dfb05e9630c3c8f3cde7828c43822d641b06eaf6a17beb1b44eb66724b7c2baeec56cdbeed29ac885dc3407714d0ea6a9dd294873a3a9941de19fb8e82b18c90565d64efcf04a1b643b8159c5ce6f0e119efa9b41d664e36f14401e430abc8e72b208081976a1c615a1dbffac2cbd2fb718724a89969c03e0a8c3a360883514da649590b2066a500eff88a5187f38d05befbe4f3db5612d4d0a21763461e694b36a71ebcce05a63faa435b01fa9d82ba0a76aeb998a4861f9e8d0a6599ab81d0a360d9ccd3b4029d2ef355ccb7778b94e435784d4d8a814e9ea92648cc5be4f16ef1c60f249ee39ddb8ec6ba964a89d8f550c971026bd3f511aa05bd5998a544aa91367b94b27352377374c7315d6f5dafe0a2383d470962009b977813ebec705b1f98ca8e17226e4bef3be6292d4d620df3fa9c1bfe8f8e560e5afd25cdb214677292a1b73bfa98afccec6d80d65880d6d360754b1223f3675fc378a042a6259540c628132be064716c5ba92750f2be43a9a860b5f4a153093b5baf48775d8e0ce4960bfc81bed29b8a30cec897ee53682adff98f7fbf68037ba931de0e352df713c6f7aa90ebc0764db4186132c4813d5ae74ea912d539d5355bed51d7bdc1109ed2057a1ed64b3ec756e9ec0b0ea1ade2da461caeee08443501705780781efdd397c05216e499a5a339610fb114ec21c0fd8acdfe020701c107a5576562bd8771b2d63a8c6466a996b98f169fa2aa7cd969991de84ed949a8612aa9f67f7bea3416fdeaa467183d7d50ba8692a54625430b46f31e64a9a9a9c90a680bf6f904b4395cf37a684a156c25b2724099458cbba131bf72b666a10070d6ce1005896209e857c0bddf508b87f546bc70bbd33d0ce14a270db371062727b1ec1ef4d6dd348d668a53c5f58d64af67574c4d532a073543fd4e5b0128856b8ed3684a4b41cc1bccefff397fec28dd438e36ad05ba44de33505ff6998a3faba28ebd61e46ed2d2067e8f0c9da0ddfe746965f70a4a611ec1681abd3586fdee53e00f588e8c26fdcac8cd5140a7bf02c82c9da7af4abf4d4cf427d1fb484c53dadef9321fb02008c57ccc9be91923b0196bf169a2a5f1204df2e78f80fa659d0c75a5044272b9f194661a9c51c5ef4a228af2eed5c9971749899c1ff7b83d12312f7381789b950b6b3a2ad823ec8c96fb2e20aa3e647690be8de55e2d3d459646a4ab3f7558777ecac279b0695b29814ca770dada4bac278f627549702075be9cf22b081bf68a72a9e69f71f823cff434406fd65af4bce9b00864d98b6ec75dc3d279f3d09c30da70ae1082070299567f69b056a6a285b4118993ca0e61e325024d16988beaaedbcfc652f802c9085e7c57b53b05e72fcb19efc9028ab51ae9aba9053ba24f096c885d43d40181fdbace0996674666c22f6a0fde5000355d09ebf20813fa7d5c25def0925ac94b072fcc570d99ef1497c87ab90d4a835296dd03af3f2c4d50e8fb12c0c7cad04e6bbc0b25d16f7f06742712441fb6d28d2912dde092ffdbf768c9cc0ae27176c6062f00e0418c4a5592431cb42b2c128557e5aad922e501ba6b80e02a2ddffa8cf809ac610115b08f5933d59d5070e4b6093991df8c68a5108f93189441ab31e2b8a21c6e054098a0bcf4677866936ef27d81386d1664268076848ef27ef34adc8dc6e335d0a732cb97c0547b41c5496adcedcf98fb3b4e5e4a1ed74fbe710f9290;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h22da546d294bd001384a25354e3b24fb320be2cd228ca75ea01ee0efe48eea4ee58ce9435d2f5d66e21627970e1bbcca3fd98d2126fe1a5f896fb6eab831a7207c68fca0cf2bf35c711de7b46eacef1352715c6749cd17cb2e297770588973a189d5839d018ab0c972d2e2270f63c4bbd9f56fc1fc0039a2c27c8aa1f1934026f92323e87f48b03dea211900b1c22aac675c026477343ee54be812a1bca92b979ea2aeb2ecd53bba96a2b773dff5d3c5584b03d3d7928df7f2e201c5aae2616df320b65f2e33dbbf8a0d7d6bcba1ede6e8fca39b88056ac395cc1384c03b6ea2a78c2da70f42f2ece0ebef1ee3256dd5d1109410cdfc8814ed9b5ce6c8841f0e1138c8f8258c27e11af4c7402dcac284788ebc533085142cb2f0ec282dd2c8ce23ad6dcd86a6dc9fd06874ea51d599b0a86bb4d885c148965539e81cfdc70141cf355a7187c1ff2f3dd2fab8f5c0551563c761d64057b20f6b66f41b3983c8f083a0f220807c7f739a62606ed6707fae79b35971bc0f6bc3074c378150e9757e5437438aa0e273bfdb272203085c2901f94a10cdb582bbcadf26c416a3ed69b2c713cf049a7be79f8d458e57a28497cd6430448681a1c3fd5a977d6e8d811f3f7ab7a1c29e0e181a28046cbb5fc959b9e8fa9317bc5183895f0ea384becc44fa82c05c6bf5454305c8c66cf4a71675db9762894ee075a8a8288c8f154bbe030f32b90a84fd0c8c39dcf2ef63b2ff5a428852439c236c16695f7dd10e95f65e66fb29775dbbe7da2672c8bb708e821964f5d2fd36f5c48ab439495b4bb91001c09cc9fa59ddc03acd4c96e8dacbc1d7247af03637d2d53cfffb53203de3a808534df3dc900cd4cfb5ce64342276c5879e3bd7bde8de60d7a4d7fe3d89a9bfcf86e7c8b3942757afbf9a6d2c2e9a49de477f74e777d13e04a20f29e12db5b41cf9f55a93d9d36e6d774191a32bf358359e63dddb1f9808ef44cecc8e4be51751d69c7c854d0497d03111058e0110bb9d5aa7a4324ba7b1c728f7aa0a31fde05bd962398080e270d3f36c500dc4f8370abaf86a6e352582374c70b66d592417767f54ca4af249befcfa5019584f01074907437d12e438c073c734e8cc49dff5c33c5f45fdd083500cd4995faa078a19264afd1b5b6de1dd8000f15252488b5a30041d37e6b345dc33f11ef8c32f4486a9885c069dac00c80cfcdb23702ce0007dbd9282e854d00acf111dde8ff27bccc50629a9cbe4f332d0c5cad73ef476b2bb9ab146fc995d9e3b3bd8c410620f2aaa12bb55e8854ccc512181d47f5af077868902d8f6536b49978746af6e15f041b5b3eb175c9b0eefca21cb9c242fad2776e13c805e13cf720088a5d59126ba1d049a336b89a37773a952d446510d984c1e42259d15d1f65ef0a9a90db68539ebfe1edb54809e09ebf2d072ab0fddfdc1d4c81f95a8806522faeb53029dd53ff1f853075422b389337365092c0cd7ba858cf094713dc052e7b43e9bb0b491d3f14dbf53b46111a7b456c1554381d130a44978de874ac5f91baa03c331c3508cf49b18227e783387a9edf91210c3e4deb709e7ba02721e7c0df31e86157b87207a17ef3fe36a3c0716fb25ec46ea02438663a92d9aa6e8414c5218e4c03aeaac0ab2f79492ea03374e70b7662ed57764ff737cd0f728f82cf0df0989a5a9964b6778f36454a5a24e3ece2451cbd42dfff08eb7b1ccf2128c4d7a64316aa635cfecb321169fcb3ca0c44a136b77d7a4199fbe0fc8a073d38c518366713942a10513510056b5df9e8233f6c652599676d2467e41cecbb181ada10c48bc258a736ea587ad;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfdf1687d9e672e11f335fafdc17e77f525cc28b031b7067346a113798ef4dc8158afcac46031c9f9e9d1944a3fade8dda13f2e04fe73b53dce82752aee5607c52ac8a14b5580f360d778092c45fafaa4e6814d6e76cce3a347f61b3ae2d55660354a5299e17c288a0aa02d620085709edeed831ce4719580bb1b53299359cbf58445ae0eb5fcd35d488c325f05c8057088e7ecf83dd4f8d2b49da3af748cfa6b99bafcb19f826685562a99946723a5a4ae81482c76041716ce60e9220b445c4185314f734dc31178aa019dad87babe302290dae0f4e3b39f29d19a6e6ea3b479122e0ea28d0b1999c0ca38f1fa65cad27fa84fafbced15e739034b9e86e7242508879be8636d822e765ffbcc7bf6f71137443771f632f9daf7f205fde002ac357337cfe1b56c8dbbac07c2b778929b12599660605d184b3e89155e821ff2e0ead47e443b3ab607fd2aeaa2191e4976f38ebee0bbe162b4fcb4f9aa4847569e0801a60144f2573993057e88ee913fe87cff65e2da717afd3542645ff3e7e91f900caacd73872e4341d934dc22ffe802448f94272df13e31bd097ab0accbdf62b17c1420b71e6b612c7b2329832d11259b99a4089be78d0339ed93e5a08b16be1323bc6b85d00de78b0aa625fb1c82f1ec0f6de8e9c1e56cda164ce49b338b6fb04c7a6871bf44f9f7a8abe8746327b812f9386dafb67767f74fd15a7d2b3d80cba660ef1f27e0bdfd5328f67b59e9d4db54ae2dce0efe1c7305fe967f590b147ef0f3972d3a1de985b9d24e1986adab6a32190717e512513da250bf831e7cf4de722ee5a9481c85d2a5b6bdeaa8d310a67d327cc1a3fe866e4d23a1f27b89a873c1554956448bc2e720e315c87c3ad1ed60effc21b3cf0e29bd35aaba1f9e0c1454366061c2e7f00035d466915c116768fde92f24d64bbe17e15e806cbd823a9084753a7de205723c4b2ea74dfdca9d4b5a61ec07da229c112a0e188fc8b1fab4263f376d00e50907ea0efbb0345e335ff1af4bd22d4f25320f276473c30823cf2b03e68b306e36e5edb431243c7b4d1659548ca65f6a9f77f75920f46cdafe29f62b3364231cef9c888a36a9dd282c9f56341d7b1f6a2cd17d038e7f7891a05eed7b3d7dd300daaf1ac571cc13789eef7a8ee3e55dddbc1e21637ad78ead7b34777f4b34204a1c8b942c3406768cd376186349c43d1c748af3a85938e313116a542addc6372181a8c688d2f51cbecb589adb9eafe151958419e7d2dbc16bb793bdf1d95b802b3bf65435abfffefb25c9b006981c8f50b67fbb2c9a3d44cce51ff93f1c346ef29b549e0adc8caa764fcc8b9b87fed9d7ae8f9a082d6cc7b578138b81b93cc3ae0a5c42853501a2b0e0ab0d985c442844ff3a9f1337bb47b59c53bfd615c43667ea871a0db3c6cf34e23bae92213a8859cd0814457a4e8b7df7e5b7c8cbf15632d4009fad096aa20f57bdb1b7e58d5dfed18fcb0c1d3060e00384cc92abce4a94f37accfaace5292b5c203282b1e0932bfdd8b207bcf1ecd7410b7a8e5e079ac75726499dc06e0bd651252cfce01dc107113aa823a4a67dd2b32eb0500959fda58c4338aee7956e2cc74fa296f93330d71ddbfbdb555d3473ceec0e77ff9eb5f0dd41128cb8f6ec0db0a827703d2515d4820a3a78cb9b5c36102811124b3764563b9f6acf4015b9c6338115d7083daa650be725488ee395cb5bb3ff14f1afa006ced3aca3674d21a2db1175a828c6e2e5dfd1e9119b467db457430f76832ce3e0da21f8f9728d50453450086b9e19110cc7be626b55b0f737310dd05223153db21765e8b1990df8fb7246;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h17e6f92dc8763e1ba29b56f1dad733652683b4e0f68fc3466676fa7fdaf0d2bf25fb7cb3dab73361c371b4c94ca9004565c8f3da19866b54eed4836dcb34a23974c79c9c9194795a1457fb4b12e5e31eb4b13a7332b4194b5088363a973c9c8fa2e9442c3eda1b67050fa5da84e9ebdcf4d0739ccefa0082ed0a43d7cc70fd00ea6ad76c24eb46c8fd23103e45b326bfaa9970e54c08999dfda12ac13b3349a171b8d6b955878dcb99207a8bb949c062893f9fd0724bed8f0c5eba159d94503fb3f55f7809ad7597b201ed0b67050fbbf599758aac5c4afc4d0431e8d0f722091fb19afd994662b9a26a7d2366475c67044b79c51b9480088628b13b255c328fa7678f87d889ff56dd6bd212034fc4e279e78cde2e93794ac666deb4db98b795b02b0c35ba11dc5a3c5f4e8a8b98f9bedda97fa7897c5983b96a7034a7c2cc0cbf689500014e10f9d86d938d66230d60ea6a6bd1eff3a93801b9279a85185f80c1a3c0b548fe47248caf0335410d28cf9d2df58a3cc5fdc4f1e2a0dfc1e854a242ffe06afb50108f34f1b8061b93d763ca69ce037b01467c696fdda78b6ff5fcc1d95ef606c316d4ad926d5bffd2edbf6d0d8f3069f6d3ec424b70e2d6bd618e37e6c8163d6f5ac13f017b4dde36aff3ecbcdd574a3f6e56b00919e3f6929e1a277af73b17944e9a1150b90c4b7bec6afbd4ae0225374ceac24b806db41f2a8285e82ff245f614881275cad7f270ad407ccf2d97fc2d0a4d7cca95a4556f9e30d3ac11091c0bbd3a91bf115f02c9967f2de09aa68afd050040c92a8faf3179c770536f37b0dfeefd95b68e5770dda267d4865dc77952dc1a444ee959070d51c90cda93cb043be1d5440e72bec6ff229e8bc01b7f40847fe476595cdaf04b7a5b225ff26768e6d7111e5d1b57906ede633348c4a20ce1b0d92f2ce1f23459a1eb035f8c3f10f5233cadedca6b4a174acc4fa9a6c09de5a23ed0eac941522cc846baf91704d5b0b9f1e1aace6af5ee34b68fdf7d47c2f11ad8d2455858169b17ef3bad32203b8b3ead1abc704b63b949b0b83a554f6fcbf9c79f6c1d684165570b9c0970f72a93c7aeb634d8d8ee4bc372b703c0b93ada7d49dbea4988fe0f88a08a76751954b9437b160101cc29c97d65cd52c54c8fef296842768b2cf36dc6b55637f93104758579d1609c410fa5e2c6abb6b4589b61e81163af3da7dc9c003cd0596b4efcb1bd5ca60f9645f5e1afcfc3dc72ea09be623f4e7953250a77ea7ae3492c306e9beb7e600376787fa739bb1b16dc80b3b570131d5028c2a7bf100b08a2c31befd9c9c4badc13ab78305769c5351e40d644496fcc06da1739f377704d1a34a51cebcd1fc1b47dd758d5bde40794a99662cda540989efaf24216a163475c4305960ac91ac5216ba669d0c49444e19a5a02f12ee778dece7b03217d6ed78d4454b6cb60dc5ba50f5a2075b5e8f408725a80258b5b094800a8064379d143f98df20cb093b7b5b7b53f53192330d2801b1a83d3187237564abcf64d999961ff7f84c01ea0d949cb3bca869ef01e51a19fce6122269c93215d99d3f5281116deb000486b8075bc3fb148177f1dbcfaa73b37d70f494fbe713ba4df96e273c45ca1c0ddc7f355bf46f95d102fdba82b69e6c73a0fbede8a6045a358eea68d987b5bcfbfc50237e51f71f12fcef400dcdfd757a0a9f6f70dc8963e21f409d78cdfdb15c5ee200bc7ff918fbaf07f96a7f0e0ff57c241b88a062fb96d6461ef83abe3dcb8105a778dc3da12bc5dd53dd516507082709e3783803e1eeae13661d730607bf7bace910e2e9c329af0731c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2c340cbce1e933b9933e85801e8e2630772aeb5c3f1b63f2765f2a6385e6a571aa37910a42c577aafa0a0d177f0d2e229e6fbc7c06f17d71e220e2c3126911161a27e3f54a0aa15252c86810d2e8707d34267bf163de85fc7117f3fe83c64a5812e05ce8fe92d7de563e7711bde0286b56bb8513790a9af799d99115bcd444d76391f2608df5d89f187f009d843647d173ea1f6f6efcc5cb6e7acf8ddf3317a6989d6a7c03168999a9fb07fcb9f0770ea657e197daf942541fab4b3865991726814a8d8030151ef4609603380c352478be27d9450e76e97f2351cabde3eb4ffd9f5a29853e92d73140866907151e2d86348ec0397e5c16dcea55a83f19d0bac6128d7a9e641d5461ef26055a09b0ef43d656472957f0aadc10d289c7a6e1c6bc3a31af6d7323661230614eabfc01cdb1f790d1ec1219415964b8c240cddf58aa03fd25cb23570090543ff3358542830e65fe7916b144e47c079e74b78489706f7e8efb58a230ec200ad8224cb2720cff3a288fd6c41a017daa5c8e84af9a4085bca58e2307fe339fb2e166b2adde2ca156c29955d1243f21ca8596ca300d3e8131f215a1f1335d52878fb0927416cb3d5947aa9a864352380c737d7a70666304f527d2df212cfab4514ef825db67bd70b269e3065cbe5a3900078a66f2c075e36ec9244a9903ccf2a2a32be1bc75ebc1acdc92103bebd66483b563359acb999a630129ccf24132906dc650c3e0a72ae9dcc67f01fc96f4cce40d26c47bde5037a811449e78918d5335e4e3ec9c808839882e86d34995fd2f4f7b9e9af22a6751d9f2c2e99ae0c78b95f2b72838d700d7e6f3dc9e986e966d8c72a86384e1e4cd14e7d24f97561285d312790f0bcf14b5f43d0b8fd5227888aa5a9d539524b75a79620f71494f8de6ff30eb5400026fa5708a78fe307a1b2b40a27593a47c6e397ddea26bd19363719003663bed5161c2f52b1037c2b992e8f7f410d81cc490847080b6c3c721f67fc3899511f296e7d0ffb16f0142f1de581684d98bd6daa4f21fd7e48562643542d1d3bd838d707b31056b162665006026d264051d1470488aa11632419d153dd245d394ee77ea83f1a70ba7adc2a3a0cfc10bd4077d246a5c7aa449adbe33bb7be1d4772602fd6fd76bd7585767952b984be750f27a34175c147927284184dc3ef1f1dd7e8ca66a64f585a34b6de96d3ed93a0650f2e56530d970e1f7b65ffc1395037f23a5046dd7f744668c292f8ed4be1f327cbe40c3d3defd115807c6e70a08a58298c58809f0bccea8ca3760ca4a3416eb6da210bc1ca95e7352654b16c328bce67801194f3660b56e7ac2406cd116a2586ec49497a25a4a145a5cfbc2e04b77c250e81b7d1a22e9ae863ade32065862e7fb1f5058e2d02685ab8a60548a63f0f2b78f2fea1f456c9805bde21a83180b9f32a243bfae7b8810bc5b0e5748f6a00da3e4d2e0cbcd0ec1d039675a1a99e57e4ad897131fd9790f605de0e6554b42baa768d10db50bf536842de386c95b85134c9dd2ac2955258b0c131f274fac0b0e649bf62d15155502a871bdde9b7ab97f59957918f3507528f302f1cb6fb1368157fb3db14bb9371a9b2489120aa973dcafa382ebca5b9500dcfc686299d1d615261e51ec6fefedb40933a93dc606ac49662d4f9d3a2e855f698740573be726988ba8b916018de645a2cef71e23645dc66d69fce5c0ae41ce4a1d764b8e7f38e965db34ae855ff506ac515ea13eafa4237f73f566e0af5a502e0958a87d9553ddb2ad45959c31288cfec5dfad2849b321e913c4e95e33884b742c5f615c2c3775b49092d090;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h569ce94169108485904d1e49ea83211aa6c655160832ff2230109a385dd0259abb73a17446820a9c68ac05c0d10af72b23c0bb66b9a63baed1c4a4c086b5dc9b4d49caa9accd10dfb8f45e7b632e1c038f4c6bc080325cf95e2067aed5496d83847b7863e655a90aa18c2fb0c64f173eb13d491aa8772a6d0f822ac9e314575be385a63e766e370ba3678e8d556dd436318c94f85694d89a12339815f5c34f8f4e7e42c3c5e1018e25b0d622d489334e699552e06ae5235c545f3961a9b60431b2b87e46493b60f0fd344123742b33cd2271d31053f78994bb191a90623b4e0854eb6401a9d4c054816c53a16383bbc11b7afeffabea56ea693827b45d8070ea2704375bc36018a25f7749ec59ab3f28d18e1b20eab7f641ad91810bf6beedec46be2a7e9bcf2698d9cbbd3aa4725bd490595f0c91a97291401f50f9fcb09689b4b2534a861f0a57ac7f4b7f750aae7b307d43272142a87f36b3cfef3e3915bcfcb6309fbb6011ca1907c9d122dad19889ae47d11719bb4f5490d9d0132f88f020f4015d964326d0d5b4319910ac0d73883642284c4268cf1dee972df373d7e7f60e56d47149abd5e0239286f42d812b1ca4d9bd6986b4e9163d8e9c59a15d91a979f3bd2181b1614ac7be577fdba5af267446118f0703f2892d391dfc04265659938a888705f1563246a5e43fd23c95b4608dd40ca3f32c8889a3cc7f498f37392d8aa8d73140948a72393904701029f0d8028a596483b78486ae035208086042be4e151f02a4e1b3196960c13c16442595a5f7a769f5a3973595f90686ff93c98a4cc4903ca6be17bbb83b117ddf264f25d8c29d88e5168feca260029b5ca54b88bb5d7b81b326f7f481cf8f7bd5164997466b065c7bbb581b5c4615d9b8ec1da04aa501e7a4c428ff860f1e8023ff1e8dfaa788a0af58d44dea0d3f1c19426fc47be85214f87733e73a24916463871a6fb670b0c7f74b995a62fef7192441fdecc0e06931dbd4df59e4811cf4a5cdbd5ac8f775b01e863a7bfff9a8f73c55359cc899f8823cb4faa67c1f4f59348faa5ac692708130eb929b2615fc528886b3c149542ac5f61672229bbc9356600dcd917b362a599638fe6c2988ebe1d2d25c37abb4e7934d116a1c1d6f823ea9766996751d145e60fe932c93c124e07af725d3825c07d64b4d60c57c30f05396c6f8e53f89ada2c83802ad0142919523976b71739c9df77b42464003d78a2ce8846d7ac2206d6843f9f1e62a381df1bfddd2b6ccef0e1e6747f870291604e7fdfe371f24d17ad5d60b58902b983d96c0ff059bce57547c054e499d12208bb7ded01ead95fabe42cc938b15c358226d9ac637c455310c50071024fc5c95acbce26efd6cca918ceaeb6f24a12346d534a5dc72835f425916f561be3b27f3634927fa9a0e340f6d2bbda621d3e68df8f86982e294d7fd4be23a8f4a10ad945215ef254cebb25e1c669790e353373e5c05ca9d23e05b017bfbf8d63c2050d319b3988c2c73cd105fa6fd01d5c4c7171a71fc9a249bf12202c891810168889f5fe321e90b5a22a4041ec1b92903cf55aeb156f611ccab5279e4c203eba4588b9a916944446bb7929284a2a475ce57ab0da61625b7db738a5b784b92e2d274af5558143dd0003ff3cbc44d0a5f2a834e57ca368b64be65c9db16a78c8b449acb5764f8f229ace6b1325a0396b5d8b29f439c3edc94be8d73cca2cf728270560ff29b8183b4caa19048015d7a676e9d06c6cde9270f5d1448d1224730ce6f1135785f30c5a79b2e38b8760c1ffeaf449e1f2a8f7ef9feb0f2bf194aa481b37974178d54ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h81b6673a35e90a78f5d3e88c7a1b880e8b892969655edc9fc65438d5b7254976d63f35bc9a42870bce0bcb597c84c82123fb443c94b1f6703a8af6599cc7d0af5885da1b3f534d63569978089f39fa8ff262a391d7b41aa3a1993517c081e00661d9d78f130c0eaad9bcab699313079b97b640156016a1226fc1995728ec777175d94f13256ea019f675cd644acf880c1c0e069c8358686bd700bc96b5338be5e1ca4ac24925e61e70dc8c60e251c14f290722cd8002b5289cf52d28b33363797ce7c0b58760761b09a00d20d6247bea3b41a1e1e49c9ab2176f212b5317477319968c0d4b4d931197517739da2f3ff251fd1505ce2f081876502cb190890e5805775edf0422d923b1c65cae744ed9656d04e5744c8baca107a4526cc5278cd6b92e2629618fa9ef37ab0d496eac2b4e8f60d8fecbbce418a2518dd3e6417a013f6eaf6504630d44248dbef61f844633fa121b352e7bbaf00bd5e69ed8668108765d9291387c938c283203fa464df38e3e9d134e96d12ca3d5b872f76b2f05a3bf3113b17198e7a9e8df7053860837f3e93289fb1c58647cd2d2bd0bd5576b36d06955092f68d84aa82b450c42ee01541b0b7902e5e9058ec81310744bd90f45b4da259872ee8f25089bd772115e5106d07ada47e13e107ac4a551cbb00b4559436e9149dd13195ca67c3d93d46735830b6cd1715f6d94f30a2f11b5c89d6d65f28d9d777eb94f8c1864f44e063072b2e42b6a51c58991be593be9c93df50ce76cba56637229c8c6255dd78c51b5b6d0f17b87af3ad1636327acccfa7d41713234409724a34efa7cda01e148a0fe6c343873a9abb67527f76246147305757c2e8abc0a7f77524bf7e32cde64b35d1f70a94edea91b1939f70e0e978b4517454d027ed598ad7a47be3edef3045d06acf633dd33f45d4e4c1b75f001f344a36ee182bef8aceea87c4bafc2bc4595348f6538d7992408b9f9857c570eb7f2bf050ca35af8da7ce15bab304818879d0e6fe1acc7d1b04ae602ecd2cc34617cf3d11a318898c1b102e9990dcfb44176494254dd2f7a41a6d96b9ddc8bf943146e69b5b83884205e82e586a90c9c79170b1d0cf36f23ac77f64c31d16e09fc9440b5313ad35e418c0d62a365f6a1f9e0d4174a67e61d6ca7ad1bf29b48e8bc5f67086712d9849efd0ec766c02a2502b541eca01c93e9ef7af53ddf12588b258aa8016ef0619734ba074e14de5b3d782b9a033a523ce0383eef9a97e5f8233e53d51a06dfb692b977fa9b30c0253e69597209868fa6eff764438e0594bcf4273b6f12e40fc6fde4373b90e97f1dc49c31ece688ccb425642f2b48891e4dfee7a65ee7321f4fc88c21d6ebc847c283d2f34b483fb91d1a50863e6f07a45d309e71ba53bd0fb645f95ee54cceaf5d11c02b09f8fede5c3151da250c59342561cecc2083d171ef51725d62c1f6e723cf00cb5c0ee13ff440455ab171185f80c4155720c31a04f0150b5ba65f0f50cf26a93089d1b4e2579127dcd14ca59ff77198c009e02f489b4496d167d8a6511b89c6026d241b2ca232bf17f937a2564263dbaa69385ff9f95c6dfbcb7d4bedcfaddbb79ee895b1d90ec541c6daa4a2ecf58099d2773685e8b9280871e01ef74e866afa361335b5f3bb9ed997ce0fe54e6fc83db735bfcd1bafcd70023fbc92f67da38732ab5be7bc1a8a70f25ef6b548ea978c464d0f9a6098a17fc1810441444cef94001d06dee3e2907db172fa7768baa89a5bbf64cc742229296f3f590948420748be3c0589065e071513ab22960c55c08e571506c73bf619ef0b630cdea93c9cedeb1097;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1f9a0ccf6a607545c9a52865ec0c66a12899ebfa204fcf6408eb3c4f70f84badcd07275a460cbeca113c7037bf528e9229520f841b24bac2bd861283e177108a7a24cd44a2750facdf0e412597711894744d7bf058ea02c396616efc45bc3358921505ba519ec54d25c5b8dd32849de6c625dcec2229541c2887c02c8d7d47d7f34b51179447bf91b794d0e1f29cb0c8fd93ca6175d33c01667cdeefd19d4d6daa2ab987afe9d96bf19191acfb913af470ee616d53f5737d18fe07e9a808af92df2c107aad99f2d3a62865912a5d55835adb0a6a2729943d685c4332611c1fa3687cebb91836b9021baa499e53df94bf7082ae91244cddba3e4e986a65f05ebb65c0a2d20cdeac596ff492a756d98b380dc339d42fa86a516e34574465c580aa338d0851bf8fc806356e74d57c41c85c5551bafae046f123e0fafe070aafaf1d4ffe0e7c7a7bc6e0f87c95f1013d925c319e781550b808ce73a66c36229b9fb4555ea57ca475c2dc98669ebb25268a024909ab66294c068f09e5b487814ffa408d3f0240d6c7a9e538d47e0b2d1b0211ef003777ce81347a801ed8f77e0c59651919ce779c15537664bba6a16739ae154037c40384eff38b8ae9f8e59800fd11b5d45f0eaf035e79eaca261ff3e5f1784f389fc570159df4a7e51b4a89230386effeffc5bdc029db646ae97e16cd5bfd51ff18c8a817ca9db6547ebec988274a853c5bb8fd45d7970292477a50a146a40627f3ab3d4cbad969e378b8dbb576bfc9da42bf548d803d724f0b61760435b0a93a882eb0a1a04eaaa6b4307eaae0e4b78b93c83e161bb9042d7fbe14583ccbe38e37520ae4f5544cf8426fd5035cd1c89404bd4a0f164258424635dce170cfb3194f1fc362ab0fbbc9a03c21684031fe7bd0dd39fbd910ec7287dd4800c2c46c54276f1ce9bc770abb1dc8f630278908165ec3ae932418d5c73699a5097e3e3f49173600f73170cb0b9a78fe28d1de90cda75113aa099183f046cd390fc63563c1acea448f8ed23f5f52b254052e3916027d202714325247055366bbc83284e615bae8cc8df6b58e3bf73d3be50b9d64fbc50ab1498c1c03e2645ef8877dda02f2b1f3557c5d6f5bcbf3a2858b8d86de8955119cf7fba9fad6811009d39232fb6885f24fc19bd277df0815dd4d602ab6b3bc918b8b2ecbc8505dabeb658b7e0f5dad91b46a46a44eb72e2016e6687cd3d0073f30ff771561cbc5d0892e20c9580843b5a1962921c3f414f5a19cc639892b9bb1074723fe670f931bba2abb5103a8030228514b36a7a5296cecc4870a31f866bd0cda7f760882cb243c80159d3f9704f2635e1235698aaa0dcf7ac253ca6e3a4ab2e62107a1c7fe5f6166c61878040dec2a73c397a60dbaae2564cc12c379a8c05043cbc36a035ccb18e33e1ae688c5569e14368f370d1fa6d40ece2e234cc2b93e85fba1844c55d7bf6c50fa0b67ccf924734b8764c8eccd61e12c39ae9f3736ab0ec633e11d02e51d4f28f008e5455c473f2248bc3214c8412d14cfd0da8ce12e4094a6d9144958ef228f1710432f5d1219a90ee0afdc839a470739d10b73ff3897662634f4916c748cd9d697008715ae860af0a73239f6d0df82a737fde823deee60dd1f1a050e325b9e2ab2ae47a72eed59f5be98a470c6ab11ac88bb3e7eaf42cf3428fd26a2162c03ad9d75b5bbb7d76ba80b2e8e08960e2445b203675f91a2fda0d4a6f60e84bd2826f6704b9a888598dd78cb045cbb60eacbb8b657b2352f85688ab6bccbb23890e5e344a2c22cf3ef6aefe0a2bbdbf2cb0ddfc5c3cb06a81da6e9e2b2316c27704e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he6de2bf72a21401ef14856c15832034e5defebd134826c089edae7de7485b15aff86f48a971b289048c0332b2c2bd889aa2e15b1700312f1755307c6837d307fcd70fc9d36c9825ac983a9d965382e78eb9d4564c7fcc516defaee980f62ac6b2088551e6a8ee329c224333c780c289ddc5216a225a795ba8b8dbb3a72bad8d80df319dc2c1494c7336ca346983854bf26d633547ab2ba2d9c90710d1d03aabe302aa8671853595592f324649051eec5e1f1595fb635958b9633efecea30ea73e83ff75d992833ae6e73c4d9aa5a11ece1fc391c45a3ec94ebfffefe57b290382ea73da84ae000b8c26473e67dcdadf8334a6fcbab9673ed2c93e3072f819db686395dfee837e0fc2507e45f60a1ec3665f4eda5ccc2f1c97347c56bca16d0606967803851b0645626ec133dcb039b58629e99c579278af6e23ae06ce3a3417f304596a5f89f83f71583b556afc3dd4e8dff16e26d88be0862180b305060a0da9a70798ed85f5ace6d3ea62f7a45bb495b016966904b102836d6fb11292d3d8de3b9e3bf66c653f2bbd9b3c8fd44b2e0566f5da43fa19d1e7f106ca189ea8df250bc6c109c523f650db2a19f6edeb9776ef49e4a6442b373ad18d0ecf16c018f43024280e88ede01a68906660fbb8d076b83df955c3b4625013189a19a29b78a5781103259cb008d967203075697db6ac9091dbaed0b07f36b37b7d083cbfeeb503743dfb510517bda6d813572b6c41344b90f27807ca54dc5b8551bead47b996b98b4ead85b79be2ad035d9583e3841f38bf078517cb1f39575e0359db407371fc5fc6a719dc178fbc45fedead0a59f4c684faf958421e722c2fe09a93477c4add6cfe6ea05e82bb1602a608b3b48852516d4e535c93e421c73a979ae1eb97ec0c9d9be8944003cdc2710103a885a45cc6d41b1408710cd6ee44de7ae478ce83c2f5a320393ce6248aa1c0b20ac1f4c853a39221bd99b09f449cfa62ebaf674af62d5c035360292dd74d76795766f5a090c5669081df3dd2d19ae4d1afb2177fb156566ea53b7d6383ba42ef1e44211e2c570828de0684a54873c7ec71f62b8f5d72af49ecf7dbc2e7909fd3928c10f4bb8829b3c437d9e93b65b7cc43009829b7d68ac3afdd35066d794ddbf6a4a57c89304c87e09d7ef28e3ebfa19822442e62a4ff9f617d1f7d1ced33c83d20033105afa4e773e7586e5a42295a74fb4fb09b8059f7ec7f898df5de24a60cac2ad62a8cbbd1040a9e80f1a3870bb7b4b4885e79159927eb75b2356b9a0bb8fafade07e781a36ab97ca095c817b7825614b3ae3cbbad3bbd1e0d2de84281ca31159b25fc505033ece1eff760c20c88899af2bdf42cffe60894c5910ea357e5753ae69aff376d6c012894b23171cdd80a1cb1d9bd13701f3fa8e32a279547654e1842c5636fca6ecb0aca9924a8f527409f5dcc4c2b7062daf37ef53a68a8eba487d0e03e387366558c58150918bbc4cf1f0a4ea662ba58b808f63b33024ecfc1dd6ba9216ee5c034c37b8ea0c191fc32392a06206d6b89fedcb844d4a9bb338094cb9a09ad9f7bd6eb02fa598d60be3310332578a8c2bfb9d63d72cf95bdc156d5deac01e7cd51a07dc77212139cfb0579e7b9bc09b5b12d0cefe3df7062e2a5ca32a173ac002df3d739b00b5a20cab166535f5a15375562c094b6ff90f8cf6f5297bd1f1763796d2a1427d0722fb3054642b0bc787af7d5a25e5a20a78c98ff8fc1a523f263c246ad04c3bbc9f7fece4ccfcbe2be1f13389642b27026ab139b7f2c76d3ef9bd17107e79832337b6118c7a67dd4e2aa8e591a422b4d79efa24b00f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7f878be4c757233bdd6bbb7e3bc9f7fa7c669c08c688841210ed20844ee0ae35407d72a87000b8ff9c29d64badc1c51c65bd3ca1a63ea4e367eaddc1713c12e2b86c36b0a4e21def4494120714cd5e5300eb88cc8f42fcfd591da764eb85f11ac7fdb5788553f978c5a51ed9ac90857df0b5c10ecdd2f9063c895a88989c3898390897f5b4ad5321817a3e32225dd4eebda7e82a75a485b33633ca212689c6bc2ce2ab53e488ef64387daf0d16bfaf4cb7dc1f66e9fc4e7d9ca861cb4479839bd9ab334feca89c8b903cc136477ff97220699aaf3aa052703c5fa1cf3f88cf65e0fc430379a18a0e3a75e9d367f034f478c7821a70b3af7cca8cec5d6dc8e818efcdd3471be5a413fcd76ced27cebb186047982cc51a3030d65ee7f388ed7168418d57e7a712d3dcb068e0d8fa7d1844f568b04b58a743e26cf3dc8958f4f6bd69635ec639f5ed6808292257ea76aaaccd5b2172e3393d603eca936a888e8f82eb9ded7d6c58ab047e7e86471b35d19cfb973ce522364ef8ccc05d43ddbe77d79b9a865ee2c121dabd7aa5339a041787cf1ef3e6c5f9ac32f261afdd8ee6298f4e07fbf0035ce3f080065031540e5654f90aeee60bd9284b135b036c7d10370c86350d6f7a53239b3ad14e7cc696ce98afab15f35f4e817def69a075f6cc89813dfc307e09c54b3d5c5e56abfc57e291f5e8e5e510a4d261e700e91d39d74c742d26b0b4f63bb9804103c55a77be4a7514bdf902e83103f32606bc4d8c506c124b6381a9ac878b794904bfe400fd5a832ec6fdf5e397f522e811fda7d3dbea35d73563158c31b32323c0f18c96b48b9d0d6c02c22449861327c1b634efb34d8bcfe7f6fde8d8feb7ad635fcd3296eb5796127651e9f60bd066ac27bdb57d85c69e65f5ff8fd034c230b7c4f4a7fd0e63292c685ab07a2f79d2e8f83a18ff8df69ae3f5f8f05440b5d85e57187e006d667b6a03423bbdc024ce95fb6900d10a5aadc6046cefdb1e890fedbc8eba7e794aeb2418df8763d634216d16b4d130748aaa6e21063940993c7c1989a8be17117464adc3350bfee9070f9ff06a75272bce3206838af92c0af7dfbac0fdac267ea9982751e979176a0079fea0fed1a1c6a509fa98fdb6b97afb4000df5c13cb50fbeeb9e3206722a450d2139d81b6518c330946bf0a7ed720dabc9179b1ae25dbfb77f3bf7a2f402daaef28ed04bb9f1273f8a5e5c619e071e10be509d0aa09df67e7200bbd4d87c67d19bed4aa1b831336079f84e2f00591f9c769897a5020d5aefa06972c6356d6f9a02e3ae807ea913c7132b4a83ac3bdeda93a53beda2009b7af8fbada4461454955e79db984b942210b304ab23bdb246360058438458a50114c6187115768d9e96190b05999fd45e21b88a1f96e51815052f047c9a0c1afee6812a4ebe12aa36d83c7e37c33b293619494b618a8e539c2934a6acac6ca367edfd83ecff1ed9857fe959858fd9bdfc1ed2e85ad67e40a3e5c9caed16a0ac42c8eb1939b4e21333145b483289bfaebb77f05bc79e112b00111b8e81302e5c6e9cc83683383282c61d8b7f696fa5e8c37845bcc18b0fb6ecceeb974db328ffc5478494e32a6e35cb229e6c0d30ae9a6982bdd536c3ab9afa75337a92ce5b13c22b978664557dc6f636dfd541b1730adb04dc8b4e0ad9a7f0a564d2deb15579111c690bed7aaef15f8eecf42f0bc2cd6c91bf551fbdbca1bcd81b9aec939270ca5154f76ddbb01a126210189226eb337cf6be4b0a4b71ab4732e43f329913c448865646bbe8e681d28be1018cd08130e33eeaa6df2996873a728732bbf273ad56b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb17466df8cb34f6ab549df05d51c558d0a6455717f757b063cddff1a20cf2cc55ec17e82e4d3c65ebcb5afb1b78ab13f97e41b23748f7015826c3b8163ad1c747f7620563de44c72acc40a3cdf0bb8445f60ff76f4b6d687fd08065265a1a9d0895aeed6e35cc6fbf3c37772b54c23c88c3f932bed1634a3b9b4010a6110f3d6691f02ad9ad1f01741fc55d893573980f7d97df3be42313c89bb9151bc75bbc67d15858866b36a4947208106e4b24c80bb2c1b73b439cecbffb3413ab16d6a9bca5caab4eec3b566906afa61f87b25deec679604aacc84c4daedb54efc821f529ce1a4f7e44f180696f1ffd9854d3f34c2d1e0a7f296f7412e7dd066a5b3d4e6d591c55962bc615e3313567ff3d52b57413fb74f66fdd30902323ab834fc10153702a1f12465a383ee1d1abcc1b4288b69cc57488f12c84c1c8a96aedc6ae244311657988221ef9a6e664b00982c86e192fefdeaedb9595be18f5f4aff009f5ae44c25397a37aaf0773707ce55bfc6f621988520d116ba6dd746ceb9b47ac859f0f6e627c722449bdd15cb7295c917a5eee78300d65b351467712a01de2f9a0afabbdd8e3437e47126c4474410a295c4d6f06e15e9ed018c6999e977f4fbba95f04ef21d8ad29d0b120476cbcc846cff3d0dae4dbe67a7005bdd38ed0ba10b96b263de6fe96fa3f25c85ac8c4fa9522e0093ef3c451b3c002e19fc3ddbbda00bc79345fc69829164adf8504405b46eb8aa5ad1cbb440bcd0cd589575150457e9297775485e4fcdd888fc3cf7db91d98211c2dff3f6c071b192141c695e0f2932ffea6c07407dca65349f808207838561cfab95253d352524bc669e42e81a8d22a9e3c3f125a47a209d28427386c9bff43abafa3fa49fb678c65bec62d6f529a9cd412ecea38601b8462945e15e9d36025acf5ff63c220e5c350c5e903c19ccbd96f1cc0e96f819100913416d11ae477ebbc1697d171d83db4eed6cb62ba47c388ddf1248289e48f26454e6468a55624047fc253ed9557c319e04b04091382730a2bdb4a6eb93ac7ea016aaa34ca8e3b7ecc58a9fe525cc9d28a23b9b1a68d13a48ad10679c0e8c5d7805114532cd064cf97872f0bbc330a60e8e64b8737841ed17c2058a2cc7d55dff9cddfb9c53bf3fdfedc0adcc57d9964de51257d90f3e6b8f867d7f3a7b41da927f1e9019340b1ab61afb6fa9b6dd09164b1cbf10f5cf038ccfd185bb587b8b5829283dee196c036865022b733378b9d657fbe8c7da478da2c860a86625f5499545a36b4b54d86ba32e4ae6bb77e7f38a2e7869e35e7617452179f22ce1c45f896aa8bab5c95f9a1866944c8efb7b65515136fae9049caac004f3c65e3eb9b23330dc8072c1d327f6035f28f190e8932bd663e3d9ef607875685d2b11c9024eaebf39e0c914f39d49c55e06d480f7282134cabf9a48167d8ccc1d5cff6d4a9daebac3a0c8ce524d2293737abac881e8d77e35ff6f0c5da4e57653bc3f7e15e1ba3b3c01e22dec37277306b9c1ae00f57f105dc876c542b4d8e9812ae56a1197124e681b45253e17264da2567a15dbe762bfb5b8b0ea9d62baf3cc51460979f1be5672bc68639637e01054f4b1598988fc9951582e89e4d04627c8e32e5de576f67ac5247448bf2f0763ae34c94dc397d4e69ca498038ba9643067d6110ccf5f2a4ccfe89cec83c08e59a1759058709233ca7374a1f6c3fd6917ba663961dee9d1c4995ef548e5713076014fc1bd8255fa70f07f9b1923daa0ce167929b661888f29d69c388aabc5b3944449a892ee8cfd2a9ba22582a057c6fdd9d1fa633a7f568cbe88f5944f0a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h97fffd07849bca4b94efa1f13a3274d719ced17e54b949489052eee656b217b27883d151bb82928ea3193b83f916d4e22382cb93c6ee142d5fe0a94270654d559a0232afd7481981591db70d91e8be1a63b57c8a152e22c58f590167eb0fb792397936c944280b71ff45a16d889934a677dafa814b556e25ecdc8a16cfea724f6d4bbce81279b6cd62d5666e9c5c75dfdc8b085c5b9b86f4343c01ab6f43c142f18b26c56d4886ac71b86678c60bfbaa8e16953f99a28fe4f327c6f672b620e76f2468875f91a484ab2b529122e19cdc85121dc853865cab0aab1777f748ec45166c1b2f672c8c05262d0dccf74d2ac9ffd31d796cd432ef77b843c5a31d95305bcea3b3e6811118b578719c4b37704126444df66f77a19a8506c9a16457128356f74c8c00caac7cde0af99c59e7fdd5d5840d3bae213aefcbac2b4897971b7883d3c2dbf1c8ada1ccfa8510f7e17e345da446e713a145e722a90d8cfc42f1e2813d10b7bcd32671269cf9a7e08aff241af45eb99fcef961368f1196337635eee4d5bf87461001f3da4ea17831c377bd04e15f2ae8fdd95d8da926660a6091c27a7e14971cb458086bb3239e038778444b62068e8c14cfffb56b77d8fa3406e0fc1e1a030cc1a88ab92cda1994f93c313a1ba64b75357f6e9549875dc8fd58950b09f0e17c10710c9fb632780b9255dd7ae9810d4dddb4d3ee7cd2b825a69b96e36b881b22115bf4faab2edbad743586693347b848c03b7d1e84c6867ad19403c2781bbf16247e0fb90865e277dbc0e2be45955124f2ecf4e3c01f966d7a43d792cd38b2a09aeaf116c91e41f2b818f1799335b9e0f16e229a50d102426fd763088ffaf2c21f6ddb418a12ed3bc4fa13aa05336394389564a175624ae3eb24481695ca2a3eb60c88f6e2ab867db1d365e3f4a66a53c3c9892af1f8abccb046f1e5bd6131a6a49f92c335635dfd44dfeed7eb205ff66b04c2d427f663531f6e8a030be3c7d2069a74e89936417af4a764768dfa73acbfe186d0ee375e4e050d1e074ae224fc865079b3f4e0dbc6e3a03f380d87523cedf9c7de534c1c221b46afb7a2aef3309b7a6813034b7e1a7c1f25c7820ece972746592b1967c5f3c783f68f6a32ebf06644fe649066b327dc470c62fcb9351dfce1200eedf3f1d7321ab01fa1760fef262ad5aa28202e7a4ae1a38d1296f15f467f914e37e4f2e1d18d2bd73bc761a4f798c557117db01596bb8986b17816240f82c7cdb74becd2370f727b84b771afc8e2166c5a8728e8b5fca8b2365c14a51ca175223f7996c7576dd246578d7a91bec305a6891aed9585000e3cdb22c085ec601795a41a5301e8bcb86e6ff9835a45a78ebc92c7936feba0fe3bcc29934bf4aee138be0b52f62fe6d16a100451ed54f4532240cb3bbb4d2b11143ccacad4f08a630a7c2a14dc8860a2b44b9ef019020be5066565e4888c6608eefdc33aafae4ab6dd880c78f5ce4db29f38ea7524e7ebab9173c8e035a8dd329d51f477e29299ed9d5fe9eaa21d44df98a0c6b5d35b3b5983833018b6b98d7fe2f0eec48d28376578c19c9ec700e85a8d6a90c89edd510633784b18f97b5953209f8af5c59be2f7e411fa4c824868d3b2ea135695277c577ab9e5717c42d2bdde01b5aee8dc11b38abe28d64c712dd8b4b2d62b6404e9190e0ac05515c6b388c6a6a6d782a0f3fd6b3ccff81bd0253ee28ce2517180f8d5b9390180d2adcce854e6b2cf9567f2f42a8039f26d1599785075227c2d5358f62f4cf6bd19c8bb2210da5f8cc997361933fcc7ead55684a41d09043c9d37af8453e8c097e89de1ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2573a7f3d78b41d087315d26ce95966e00b8801308ed57f8edfdfc6fe137352b7ee78897369a7c45d606af60983d987b416bcb8f0e8a3f61d379ffb8dd89422d4fe522c25ba2585d91ef26eb42e84edb01c303743a6372cc3fbd1b1fc328ce8bf1f012db99599a745cb4629dd6386172caac3d34c7fc1a147e6fc3747e1541d78711c9d8e121341a9d9becad2c06ecfb14de031145a26bd5d4b47640b36cc19451f0bc3611e564ba1a561883898dcac806ef35bb0cc1c627f07d911aa558c90c7327b311e6fae34f88b6d74f2f2cbeb7c418c30b1d0a752b32849903ba26c8939b54c440ed05a77eaa1c0a874b55d7876eec13f01841c0ef2910b7979e17ea66719fb4064ac43c86be69b54397180190d6729d0529f22357f831279237a1a4c724a49bad6eb0ebf6c8502c8294752269eef07ee3f2dbf079a1829cfe79f4d0f8e2d7ab64e68ef20dc0f15029c8e1f87da5d2be86cb0263ebd13f9d5ca89a6a309349e8a4fe0d097bb4e188056cd23ec7d04d7199fdf8bac9cf51faf4b8a75fe48610fe1f5b7dba753ac3905d12a4959c3314ac8b59ff4530e567dba73d86cc13bf51f0e2d3f9ca6f07dc24e030211d816fe87eff60060be3855b5f99dba1dfdd09a6f5c0c6b56e7c844194bb322c264dd824a574e8a10d89abfee314d016d1e15ee7af55a11e80a2c1ad0b9fbda55c9f9687203dbc74ea4601c4bee473a8b006810931a227e051aa4249f4e117940e26f7ee3fd713096c3017dcde3680d9d5b0a4a5e5b6db3ca4dc50a150d3d69ccede1e166f8c1d51e4d9c133dc992d4d33d8ef9201d74616be42b82451316ae2982a3c16f3ca4f3fc674767025bbd3ee1a74357a0ae9c91054ce1e3c3e009d790c9c89d0f7f88def457c25a99c0461c9ec0f078867291dc1c156eff35aa1a4220e3329225e267ce4979842602f859444b25745fb2a973c6e21fb1bc91992781513bcf74a027109bcb31802cdfae99e35f44d9624915e39581ca61977f6e01da3223f12b72e2eb8eee662c3abbfc7c4600e1fdf19888f18778e5c7e48a460409b276554c185dc6641992a0c9b82b0a2b5f694021b4919028444bb9d8d0ccc4eb14ecba1de5d023c5d6847872cee5afeb3eb01020ac3803e8297752a982f862686a3db364900ca2f54ad50abea5ecf1055378653daf246ce3610405bc76fca18a543d7a7aee73d29bcaefad752e017ab06f9b57c49e7be22403623703dedfc964fdbbd0ac1c243e1046c936ce81c329f9d5addaa5a591a20b218d7050e2692caa3a82c217bee19ce8f59760d7f6f377ed44d9aa47d1db950fd82d691e256041408744b8bae9fe95da0a3f2dc80fe8bf06faae702a2057c2e5b63803fc0bbeebb3038c0e0607c0597fbb37aeaa6fbf6868df7244ddbbed3de7cff50eaa6c585132d791a369ac9495f9df9d1247f8d6ba7b154991b3de1cfec163246430f1d6514409ee8756ec05f0a0166b0ea30256f0645a082737256666f69d6d0077712366ff79de5e79d1029bbe5b76019d4b1db385d7b52a2ba9c7fac2b204c2e3c634be2be8a220de754495fe5c38ec29c16d23e858bbaeb9e5886ad4cbd7cb7981aee1724992fd784c7adf5d20c3de02849adcd4b0dc1b7515571a2b3bbdce7fa755f949a7e58dd73787d9680b49d8c060e380192484fabacaf6e9d5eb856e89c309ddca1050e10867e904fce9e0599be90832cd169c90c97495e8a9abe910ee7abbb9b510ab75a6a94c77a7c7233d147bb7aee6859a237c65de17755d77c49969eba0481d1a41425824dccf2084467a03c0cbbbade955c10e66793cb0e83b798cfab5dbed566;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8616468c7870ff5a200461be57082a611642aef0a2231c003270562aec77e3fdee5cf0ca70de6b1630e94af7d9890c8c5da737fa25ef4825a546b1acc9b811f08a50152cdfa90dc517280dc6ad434bc0403c3ea7797dc967ed4be60bc668fa12323e3f5db6c9dd84a0c8b43fa9f986dee729cb9783c676a05d195e55a9515feb338306f2088baa51502096d7a74d34a36328fa614780339cff79bcabfef5649275acfc9119889b532a41ee7229b2e61fb36bd0d4e814ee144c7e6e698f940b5ae28ff91140918a1eaddeb3f031a5066d1da30f63a4d86a5bc5d44b88774e59365c5c18d8541b37e63c83074fc6b803fa9cea6d498566acd38ddd195e4f997f09ebed0d74ca21bdd4c99e5d2f253cf6f71f1192d4b9aed00dfc5da4c42f5da1978f282b1244460d43dd2be702a00e825c112e1d40c9b167f25933e32b46e70f588c93863d95e71b16e5fc133a161589b61069e3c2c1a5e4d3cbf39a4c6ab1f9c2889bcaad2160c18fd0d68b539005ba76fa96726024b8b0568101fc1e408f6a29570965004bb57802518cdcfc0357c7ad4528ea6a64701c073615653986e5ec57741f67344d162d68248078d5a5123861297def142d1a1fd3e2c726587f5f3a441e3e264a84bf682ac29ff342b78a4aad75a13192ec0f384b7d87fbd32ba3e8fe2ee7359bd2702ab632b7ab52e271bb17760db40ce6b00f1e57d9e8b7c4e93dace3b529bf5bdbfa52e4e60ce1f1ed912842b3fbd95fae4ff62dd40559b505ec2f7e1794fd16473966eb0634f95d9f13eb9da9a7b67b68c0f095c6f4e1594b06353caa2a24feb6fefe7f05869c8a44345b0ea0c6dc3d0fbd91a9cf6de3b5778b55b86d2a45eae19a7e70d47aecf84186e21c582db086cb2093908a7e0742e7ba8642e80b4637e0b3c992d65d9fac2e05052ff616c09afbc7b97f80ef3b3a5ce8c071c454a6c173192221fa58af400f153ca05faa85887f4133a5c7139655fbba03ea5912eaf1dfd02245e16c029e39d196b50645e2643c4a2d791145c3af6b4f9c08dba8b4a407f98be259a0d9013d26912d58c263876e203a76a6bbdc51df1fc010056a30550b478fc5f4fc06a3c110e19c1ff4246b8309f84db25b31cfe5d6cf56cc2bae149c64e4a8477dfc93ac583bb07be1137298dc95b2193c7a52fb2bc3286c85932250150cb054f8910baf82f0c518a2b1c4e87c74974721b53fdd4effbe3cedf02f11b1dee4d8db0403bfd5cca7fdc17e8aea4c9dd65b3a84c72b2272fa0bb136ba856058b7889313146bfecb33ec1b0350525836e11dc4d852be567e2e8679bca68c6ff5f841f28117ddb1a1b17e800190a6abb8a3d14ac42ae0c87cc789cf8caa2c601674298470e40d94fcfb2b94180c4ada1e21951a8493a8ec59cbf1ad15ab40270fd47cf4bb2b92255f915201350d2d32fe285059df21ba7313bf496deb35be32241a37b1bf0b761beab40fbd32830fb68589cb24923feb103e0ebf54780244b067b84292fac059bcf506ffe8f08413bc8bf78e8582223446a4f72dba722681f81408075f1953a372eb1abb686bbd99e9d0abc0ed4b7f669c4775e7c6247f1125ed6e8c297865190a2d68a0b2cb1cf295d055373325d62ffddd340aab456fb1b11155aa52f3a5d2719f5ff7f4c54abfb0d6f234530b252e12c6d469ecbe569ebc22ca6d280520cf6c13c4420aa1d5b48661c222f790cda2299df3f58452e1f940a46d23394ecd0e70d46fe31adb126775c1ffdb2c8574982e42de615ad53bd9a259debba8a84436548171b99475aaada40d819701780620e8d73d713895e7a79c7f6da6ccb8b1e74ac4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h99b37c07bff2ea1693a61b6c10c3ace3550725bef4ac94f49852502546f5b043987d8994f599aaedda4be05d8a17441d9645abdd7c4d1c4b72a1b09bc0c3c386dec4dd5842d82ba27c7241c52f3dbd2bb798696a6864256058f91be837dec32e51cd0c98dab92ed39baf462be8a9fc5cd82e61295ea9a8f648fe256243d39cbd605abcc7ac9f49947fe694a5abd5095a71b90eb30226566052e68e8bf4257380dfb561132150f51679a9cc617c7736e1aead8f594eda415565a1544275f82bdda510aa3a471703127fcbf5f8d08bde8bb8589d7c2c5e897aa2b903cbec13b54e404fc515daf5923b6fff7e97ea91f749556850ce66b48154e4374e0540b460d221c85048735c3849192ec29ff4fdc66d88ae11e9284c1d9587b4bbdbf59f4649582c6a35affcd779a484110e55ef0bc6f9efe5d63aba77bff10ab6e8d3d4ea7046eba0a1a52a2bff0cdabc472650479d95730df9dcaef3f289826b46ecd440aded3eaef0ec7af218a177f9e9507f97fb48a58ae517a86bf1cff6c053fdb6ffeb665f156585c08e4ea89553a6ed3301e439892a4832427e8481932dd2c4972a4ea2375e63113c35d1a3d3513b0d33fc7ef09801f48c51da933cbe2974d71bff996efc202a6be3433b1cfda77caea3c01cb7ad075121e0e40221c8a788144605973923fe203a75701a3b8165ae36773b636b9e19cabf6d532f907162d711e8866f518e244f97fe98ac19a37ef6a135747d7482b3a951bb4e927c3997d7cb06c8083d292f7dcc14264f8633a7328860ec590cf656d9f3511dfcd00bf8a7cdb80770403980a8f2262b31f42818017f95c9c73db5b515ff694e06dd90e56d1981c7d3c332dc91b8060026a87c07640964fb24375b8d91a2ce95976e7c113769fdad4deb54c603ccad1a1de35c7a1847d2324abf46e0aeec9b23a4ad6869dd0835b9a9b4ce35b7792e72bea97ead82108fcd951a88b43edbe08a476cfc3d31d72ab0753183557d0fc3f1f1bdb76479ef913414043c7ad4029c2aeff4b5a6814957a592417a4f2c3d7a12837553a3eed413129b6338f0912a5911695f88b114f3e330a3ba438779efa2cf4c4f5a1e41fa2b503e06bcb1ec43d38841bbaa695b23dcb0534f0b0173b8fcf944ee836a502fd1754df728b8f8a923f63cf1f4f36c48eab61dc55167a9b6d99bf409583621c7a2b4e3d21ac86a44722e5282a43db326b0ae62bd20803ae59f0ef421fd3d64d86b72ba4aec2c20ffbf117da407259bb20e803bcff86e0381ad9963ab9bb5f795f4f138e8804408fc0cbade4ce57bd4eb75087aa05a92721108004910f8cc134e4335a26f491a01b48955e868a35e47d067ca4657a09dfb54d49de42b86b1bed4df2568b65417306f4a7127cce6d0df5e0dec22a6908f82f41d00d4a33891a0aea11a692f694a9ee4055260edbd7b94faf89df6194b1558a2879da43b508f2d506cdfc7185fb1362bc880974f43f5d822564998fff40e7be85904d30512db445b0060583c74a3611a9f75aa126b5abacb2a22efb9daacdaeda4e20b88dc2bc08705d06ae5836412106a3e9d40f742b415de96cf96961dc7c5c8310e76358ae0c828f864853f4580fabd79914e018aad96d388d991e9e82c8f9f8657b8702776470545c536dd95d3f988eba856f037da615c094d6f2cc6bcc28be06de4d1bd9d079de6d8691485f800b6f4d4f9f379d16156d72c2c963fb79344ff305dd76d35fd8ed68e54f737b6d053651e671501ebd55161c8cc3c4a21e8d37f38d3f083d434c06b830f11aadffc57945f777f91757905c16afe6ae36c7066fc6bd6127b8a52e4abb1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc3660a69c9f5682d0ebbae5efc3f0a6d6a4b9663614d51ff8affb13f391c131336723b3143297967b104edaa305fc32c03ea6b85a7d755ac3682c94ca908e737d361899168c18c6e94f9552ee12c50f5e0c5def73043ff3353bb314e45c666cd72877ae878dc1fc1d98aeaf33f4c059e49ef39fa748c0e0ef4e4f28180a0fb7187359682dd5dda9309fbe612debd651846ea1bfd9adaa459ee1910d91eed4c8a4664f1b503c187ba4214a671c45dabe7b1bf5a57533053e4af6d9884291517920fa5089f7f0017ab0a8dbcd25cbe4e69e02c07613c41586502cd8186a6b4edb6953d2857fdc235da1f892bcc89526707e2691ac1bea51ee720bd05479eef7b321c3c90ac9dbc8ac0bcf6c2636a0fd0a5318d34e6a1022eb050fdea9242c4a629a7fb645a6aaa7acb12b29b1a952358fabc21fd330ebba34530217b778864c2bff95dd1f325b41f0549a5f50dccd1b5c4cbcbc1f93fdc26663d2ccbd5f26156fbefde532cfbde89d65e2375fe619badc69361ae45d9e6ee881e8cee959e3a95bd3267315f7f3cea6ab79eead2ddbee012e83e11db112d2d0facb5ed3aa40a03a14c554c2f63f491d4fa1ddba8ef867e86f2a6096d2f24790440d38e6759c44727d56103059acfb31d406e62bcb4c2c3fb83ae626f2bde0ab47e19c136810234ec9e6a462a0e54acd0bcec5b9433b53967203b2281215faf9f3e16400425a941256862fab3331e13f0cd04ce7480f0b1257dd17b62209a8641e6618421e8d1519370042845d8084f342fd60fc6d7bc6ca3da20f682397fda5ac753339ffe02a274c67434597a4039b66fe6239e5edbbbe198ed8a8439f97f804ed86cc6a70e0aea9a1f8cfbb26a83e10d511be1d94bcdfc9d2fda4badd4c9dca808b6070e032b7be50ea316b977b25828826d0421d0b7a737187bc4f1fa8d87725483daa133ddff8acf01fe3a7012617058abfd65ced37517007c12a1fe40fb4a2c0174b84830fc9fd862cc95a720321ecd280c41bcdfaefe3529b1290b3f93506906376047dca17409c6377579e982559c1df9532f13e58b8966fbbb0d8d62f1c27c838c525eb313160bf36b1f0d6bfff0e80d3e177d0a98d824867a0bb13e9120271ecdddd4c8a526ad19d25730eb7eca59f53321ce85e86dd51b019d1872a223f9b0ba6d2c326cfb91c12683490394ca19e60d9320e7c2e9ffe0a144aeb0d9615d3180556279619864a2c520a7f44de309393601f227c7a1a6713c62d7a01baefe347eeeddadf2d042acf06811d3be2f9d71c89917cb8ec932f4b3a156cffef06ce21b9cb5c9c2d7b7ac3bdf76f788a40acdda03ad0de2eaa9e8ed00be674531e33b8fbc184edc5ac401515070e6c66fca21792665dd1442799e790fde1e6ae5f722a03ff555b9a35a1ecfde90e50296cee9f3c2a9776e8c05d125943e766e1512100d989c85395c02fb42f1161c1284c85de29228b550f1778c0ebb3d10e2f4d5fc8a89eb7e934dcd4331bf8a66485dcaae2e18d4fa183ee04ca6eac4eed13cb7851ccb5d7fbabb200e4b6831a80ec5d0a66124fb0913d98e5ac31ccb8f0e986ee87f6295d03a7ca50af50654ed790741c5b974a32399333f9684f9be56c77f1095fa8d224c93309964a4996a6d78e9995b046456a5ad277c38a262cc3011ad7132052426fdfdfa781d5cec41db5d6d198fd02dfb57f7213da8307040f7b5368d76c1478e73ed5f1c0aef80ebaeae66395dbbe289abcb4067d7916b1879ca13c5c8e9205ba0953989b894b7ad1e1e616676e1e5bf4666c765153d12e3eb63ce2caf1a481e23ef0cf45083d53f68285dd729851c9180;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd829cb06d2a8b905961a2d1ef24dd52c51923d8eeb9176bf0aa85962a4391f3e878003c3754820e000ac35df0b665647044138c5fa8eef723d42e61b144f1f20437820ff264a40a3212e184a8ebdaf9e8e14939125f3c5dd4bb46549bc4b35bc5cf068e64df50ba63c5a310608e731ae1b201c4967ec199b70ed595f1b2c5cfbcb7f3e8e1b6c812b10378ebed5169e925f292c56e21904c2c504c8490f85e92c6a636649641a041c8b5654e79bca8ffba8940e39ccb933c7d3ea155cc221c364753df43293a632140aa56e3a7cc9551b8f7a839ae489b3d632cc8a055f0d7b0a0567b62e431b183d5ed0fa426a1908595129b9a2c3d6c9931dc051c4054dd38df6376056b56235121004bc8a59c39d7386c4eb120d5a1103a669558202204b7308298adab0e8b05997237866f85a7d3c0873a1d296e21d86ec796da757536e8b9d0bce6fe3fb20afa05b6ec6bb583638c109e6c77f9aa56de2a2b5edf84c7fa2d668d5f803a48abdb25caaba238014e68cf419784b38a71ee1408e9545954a114ece4742ad91f5eb3ced14d5462bad0c7b91399e272e097e81132eab6e21f6b2a824e141954b55d38d8b7bcd5fa8c20ab13ce1beb91317ceae5792e7e6cdd8f81041b6d0648d6c0c22b23960ae93bae5c137655e821acde2a56b776ecf023d8504293767dafc5154b30ade017b9270a2e705ff4ffbe31dfda7c4b724e108b1fadbcf100871962c670ca441137230a6f601874c0b39a7b1f985124d5351e8fcfc17629384fef9862bb50e1d805a98c9664c1759d0d95b4c474f69fd38d390ca113febd6186138fbad407f3aaaf629d5d5c9c43283cfb25bc4bdeab6ef5388fe0873cbcbf4c96b90ad4dfc7a2d9b8c3d5f5c17c40b8964fec5de7a629426f1babf04c79c27026a597680ba0fe0f3e2f9c570bcab54c65cc0274208aa2e5ed042b66cc2e84015cd89b08e6271b326785d65238225c3baf8f400969b140cadd09fea38b0b4bd4f136f6f91c967cf168250a69f75fe6a952e1c8f96c1020cba88f6d052e0c7b4fefaadc098db0cbde0ac11a86ca5750db4d37d7a597de09d5535028afd3b7ab9a0606fe18a66ab8ddb7f3b71b321158edf13235e82b68222bdebaf390b02974876aaf0c7500544240bb2420bb75411ba7d5d6ff3fc50f128b0d3e29d3808403cd285c121ac944212d7a4d37ef07c15167a2ad6d55642811b4e25522547521f5bc2049f9fc7d237e071f73f8c3d2bfdfe75ff6bfe5689a5775dee0d1bd878b8859ec80065890062f0403f8a203916e40d67828948300fdb0979629e2693d0bf3e88929f028c806cb71b021c819e4d3d4883455e66e6960ea356f986cd17a1498424890b92deeac5507f29e69c22cdefddf0716e06a0780ef157e17f8be9f9f6c7e2f3b958588ec60369a1c6adda3a67f66f304baa98fc805dfb193e32ae0ba029bb42ab1d6742c65ffaf9e6891dc197d81318230a366a3148d0ad84b26c7208b6f4348600dd840b8a96de59835034f3ced1f2d61523b2ccd1b2f7502bea360148a9f23ce1e45b1cf50c8e5ceb6c322bd38cd43c8a5f45c94dea392bb45461cac51ce57f3404ca0eea768bf53295f9436b191cc89ca027a9b7889a3257038ae92a9cdc7cdde6b4775d7b94700aceff6a6c55b3dfaa06ebc90f7516f9c7de79394707724173bcbd5f64cf235fe08afd8580dd20ac3e03bf5ffaf61502e0e3fdf544f6314368c6889e81939db5bc97bcd14c642f5d37c41957a2652a3c0c126a81ecc366d763e2dd3ecc84a3443f0f2f721b547bb68c333a3055792f13c170bd2bdcf94021bc0aa5e5f57b992054;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hdc280c8cc4495283b89f38e1c0c1bc07d0fbf6e49cd2049b35edeb7ccad87ec5cc756d66bd92de126953492616b4316704e3871fbe000c38aefa0784d6309e4c3bed5d87c96ea9fb6b79830903e9d61be0821040c0a7daecae25babc9ddae20d0b7a3d8bb750b1fbb902d5a69ce8db93243a60d06e2a70abd394ecb19dc37049aaa7cc16b5281744a9954cc9fda61682c0622017dabc4a2c95ec3fdf7604f31e79f7d1d090f1e6f1edb53078d2a33aec433f0b19b2d9747a180d194fc8ed252d35de47361aafaacf2ca3ab9f69964bb587aaa3a54204227cff181258dba4f21d7b30c332ca786dd01c9f6c36b893c62f42b5cf9079046423d4d155c192411123d56cbadd3dc55007fda0ce4b75116faaf864fa47fcf40d2b8515611bf3385775e4c510985ca97310ffcffd3d67f409403fe77ab7930bf16b5348c07f3ed096f293991716cfefaac0f62d865ac4ae14d8c8c1fa9ed30c7d22cba03041ff80d67c8e957348178a0c272f763dd8b46a9a616b75a4b361bcd1c146c029af273a648d7e5789020b3ba718b157ae150a6195ac0950d7f5c8cbf9d670e5e78a587a4ad11c35947031fb297858f36dcccf7245f59e76015d1c85f90dae3ded22f68375348e8a9a61b003a4b50395687c04536888a3790b0f31792cd47ed6c8382e44073eb9d129e833e5fa05e186e72bcca211d9e8d537b79a1ace8273c5c5c72744695b60ef4db4e48c7091be0feb0a9e18436b28687934eeeede72edb48ecb5664977690aff5058c85e74c554bc1e11bbfb59ba4e8fc5f1a934a77e22f7b32b450f8f6ddd52632b82b1ebe1e9a18c4a23f62aa43238ff082518c63124f8bdb50e8df0040fb356c5a2bc88a8df001ec126da1bc2780864d32b40da82065893d09f499d98476095a5873565e792cbf838a6131f07fc8032b9ff482272a9e68ebb5325f9c3f7fb8853859f4080cb7b8073ae3e139aed5f941e5e58ae9c876a77195dbc6d745e882bc51290cad188b439297cc20d5b10794a57edf86436df08ce7b328fd8810cf252bed7b15ad3f18b2507b94ecdbc2c38c968d5045c03d523e380ce48d6886ae469b395bbe0c7483ffc81a6f38f2eff2332c23d0620e0f8d401a89c86aae75d0d390335ab5d340ec38cd4364db0c57136e4fbba92115c5671e410404be95887e55c51de0466531ee70e3ebaecf1e4f0bed605122a4c6cc61ac1c2c45b57001edc7dfd580d2d5bbf36f824d2febf24ea3d6f480e1ac8f32f772b4f1bb3233e45e1d1c07d5dc663deb42d76ca97d00c3d53839439cb87efba977afa7ab21fa07cbc4af774d51c934ebc73b864340baa4b7b17f29dd2b94f63ea65bd059fd2a2a546a0e67bdffa70f47b74c50dff8b68b6dbb79b1d5ac03c50052e8d96ed1ff8bca2e7263174ec937d66b31bc15b6fed3ea1b0c6ad831be4d720be448d6c2c3dae1f7618e4b39f7236885db95bddb4fd1c7a7bf2583e12f55a1fbdc77522504a8666eaf10ba409e2fa97843550585c93eae43598616316a37be7806d4a5251948262384a3fc2e6cedceee868117fb5535558ea8f4e5cb503eca084f54b1ea18d3c0b94c0132ccfd15f9140a19f06e1dbb9baf3d60e16ac5a3efbfdee087b5b746d755a8faf2fad2d078e007ab5728ad6a96a5bcae4fc621e68de7127a7b9cacf07cbd3a55ba7101b373f07bbe456dac7962d60d69bdd6c3b6fe30708a3d6b34d273024dbb53521313130ffee7b4dce7fdb40b8c49843a34d5a9075cca4d02a1ae1428baa5cd7db35fe85b8bb38eb52954411728b1b3b46d4d34a727e6774dadd830dc8d1dab06af1d48225ac8fd4e99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h675582d34494d9b2240e9acaefb463b416415f1eafb4b34ce8fbf8ca9055acb71ac42f59183dbd10fa6ac5b98099a276649a86a004da79a56127b1f7d25368a84b44bb0543d2d7a5415d06120d864c16511f2c4941c9b583d40562c3fef3d2ede2b785b7c98ec7d703df1bebd7f781bbdc5cb26f7a22bfae15d5ff9bede160e9be50135cb32b538866b31204285e0956b6687f0e53d9f24008e2920bc2327f9e123b3cdc1cd06057edba31cb528228a86cad120d317f2927e8d179804cfeed64e53d6be1d3bd907f4327eaa779a4469d47d759830214f902010062a72dd6834fad964180cad61641107ab28519826c1c6cbebb9a95771e1513787c622f82f3c10648fc944fc41024935727a03896c95fb6df84c0f6a0fa8051fa801431771e0b373265b6361f381a567b4568294fae977167002b572846e6cccf6e520d5a6a64509958c58c44f33c56f3ea0679203d616bb20cffbcc12d16414a2d94c118aab06413a9fc24f7020f9546618ab3dfe237937ece53f15781c1d6e7a6386eb103282a79da8339bec0108915dfbdb79eb652a505230937bb58c2235490d2d3711312d56c255f902403cfcb9a082ae153a1daf2d6a1be913dfa2a500a23fe499c597f54cd4ff21b47987d14c3edfc05065436a2866979f3a26d23e3e5f0d569765eba67a9b2e4055a0c1019355a6cd895de8fc00667f5d548308e6b182223ed37d8e1c00bf00787a25c359a1623a199df79b6d77a00a62b9cd377dcc0bf03b4346c09150801019c7f0680f93013cf3e94c4da9129e2fdd366cf5ae2486d6a6f1a1b8668bd7cedec83569362e10bc4cedaaea14585c3b7e17cde98b73f55122d1d856f6f81fd53b6591defef8890f1204e63df0dd963479a660b086e3789831ec038fdb31b7fb8144ba0fa3fe609633c2b99fe45e2c3bdc863902aa8b47808e869c1b582c37416c73f4b3bd7699f713b907d65af87cae0ef57143c4eb78b912879560c04a0321dc5288142ac9601f17e1d56ababf9308ac44a8ccb6660c9fb88ca1e3f1ea1e9fbf6a1e91229a93d9380da1784f4c667f796e6c1d25fb47b2bcdf80a746b7babfc7b6cf0ef5855bce119d2576f598a791f8c6df0be61ed1a85a7dcb6edac7fe8519b3763faa8b1b16d5de2113db4ec2e9c1bca71c3fd9f9f6e162d435b80cc2219f7be2e11968eb974c4a6accefb335fd8386e1308f9a45642f67456b99013c0e47fe698e861e9d4cfad2f0ec31cee0479f04a5f713734bfd815aa3ddc21ed42d2df5c6e7771fa0d17624a8f6e05d760157e0139d1deba0ce1f8eb4f43660dc143cf96731b4982ce4b2112298f050c0b452707ed694f673968669b7c9c0d8ed9920c0ace4ceaabed242e303452191944ffeb86c9cc9eac1c356c2f94d41410bf3a633677b3ca3a5dbc68b6b6364a164dae31aae6460098c82338d3ab8d010bcece9a5de2eb1c58896a6147a9c7a6bc842ef20ef89b3bbd4b1a9e5c50387733db0aef57544a16b2a06d4e908363956358a677b832abddf62a825417ecba2f84b7b24daa76a741aa37483b626d1d1d0dd3406626fd9af519da11769be74e7b5ee323956631aa1f24ce9ce3010ff545bc99f8391f7f00440485e244fe78447103681724d6e8f55c62c6fed9f320b23d96fdab999582d6f7f65411dd29bb52626d3f798fbff4eeaa1fc0bac8ea126fa9851413bbd7654107b56500860c278a19bc88d8eb3fee0f7fe1d36423be40324bb7b18f0cbb76a7aef71beba6dd41830a00d16ec5e9d879136d1cf3f6547d95203d7b4e0c9d44ac45ad2ca1e3cb20450d787bd2d791f3dbe26982f877d1042b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h64bfc66a7009685a9716b237473ce6c8b97049e07d4012ea8e7c7327a215ac7c882961652a21f7c8dd5e242f6c4f2b81321cf63139d3ab75cb3b34a863d52ab38c9dd2841f6e9910079ee7201f216defd32dabb33c6119c7d9fe0f1ab847558388219e6da866eeabb2044c7180098ecb02addeb5320ad7c3d9310cfab12b57df83956199ae971faac40045af2e33fc472d394f95b62bba57d1d5cf537f1525071d22d5363eddbe32290a46035aeb43e927e0a70dd3533cfe15e3b4179d548b46f5e8d765002e54a2a2a922c71f8619cfc524abf613d0d0acda88d9d28863918c11e831bd0ca365acc2cf30f883fe2ba1b996e4f24e3084752b04bc13576811c76b9bf8357a1a0c1caace58736bde1c3af7d67079a7f7d7066277a5e00fde7d75d4430d74c534d9fc0e0d8e81719035caf4d3d2fee7b72b0e5b13aa299b8d14ffa8a370a7d9f4ff45921da017f09ff2873229d9140d4b63ba8625bfc3f16d2f17332aa22d671ee39f87364fbea889037b1395f06bedd9b2d39e3711176556b542d21498da7335226618c0317311348232a05a80d978200c2abece79b89316eda24177fc2520e7e170ead00c823879ffc279a68500ac861bd3436b135fc9df0354c081e1cd53e5898151f5462970a47d9c8feb0ddacde98024f538a8751e5a61665a9f4f40539e924ca210cf87bbba7bab01516c0fb3a502bc40f936b88bce722797998c3fdb1077532a36ac8c974947caa2d8234128f550f8551f4088b64d9a1852e227e25b4bd2b99d6cc0e2d61fdb2ceb15e01f58b6d50afdb4de5140c462770b4af772c5495a153728c9926a0f5aefc36191f8f9a122906cbd5c7ae4793cb993ac19bb30c2151b5e6250d346f83b0b55974e5f296b07e042f4e5d4e0a16020d919142695bed3360d3544c1f5bb7b8a0b6e322479c51305aa8137f39b773f7e56bd000885fb4f630d3a1954264f62dda5c38558109be2d53a7f0e7e5ed412c285568623447766828311445df24b0cdca21066b20e2f68f215892d52acb8dbceefb7b959efad6f0171946ec570e18fbf66d4ba63fd4943cb1f048a72d61f3ef42e83ace5ef8659f3dbf7076108477c791950e33afdd03c049b2c5b2709deb95826627be49d60e3a6bc510edc9e56ed3563a64216cababb9341160485dafd92e250f4d22a7ea47e20d30cb5f858523cbe0bdc1df3538fc83bc4c7f33649367c2361cdb04462653b86ceba0504e49320e15b6dfe6cfc4a2395a48e000713e00fa08d89f9eab794c93318e868673b16f9e18811b4073a3b2a9d1fda836fc40ad273df8ff2320fd427748cb3f81e35cd4a83178b1906ca27f950c76f7141eea6538d33e0ea41f2d286b5b083edf5664ebe568890f605e83afd5836400ffce2a9341d856b5019d819a7fcbf97adfa5e20e4ece8ce6fb72ec1f0afe61ac403b0b4efc0a10fa2f6d5373c76c3609338af8a9db7da561e68845407866a5f2c2abed355a272502b8b132fdcc71846ee58d2bf5bab55153fd4b2fb09aa0d2a8a5fa63f3cbac5edafec47857412bf89e4260251c3fb5d3e5d36f62047c81159a0d4d48c56a12719389e9e7ae0df9c787cf187b32760c6ecc80cb7c49b257ee6660fd41a0ee4d851bc5fd648eb3ef8b871ef9a9b9c4f3937ae3712c846ee1f41d313ee3b47d26028aca0076f876e70bd222019613e5ea9e393508c0752b0c96f83e101803c16391a1012a520b005dda793d2c743edd6b191db6d56e47db38dc2221e0d6a26fbcaeae97fe1db9f44947db13b18bac9eca89d745cd04aae19419d620597d8ee988a7ec154d2d61c1f8e4240bacb41681d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb56000500ba334c8b96d6583f2821b2b99d1027544f9c4af019911065a82d77bdd7698a15fdd869e2d51dd384e3872cfe114c74c641a306b149602a7f068421db609537ce9d3a9eebe93bb9bee28093feecd5cec663231131f495bf91551a26d5c09e1f29a2ecd1f6795700430ecbf132b102b25297eeee84bc602a9359b5a16c18bcb9820f3980f2d2bf6e53c960ba45933107f53999a3ac7b19444a11eb7a5e5880728f653ebf35714d1ffbb338b8c62d67f0781b739b4ec0c37aae3cbeeb09018ad59e4afb9bb9250f925c30d1ebd435922e51515cb5f4fc9f6226f85faea16fed3b14fce900de9c18115d9a85034abe23a220bd5a318d25e7bc4a4854b4052e2268c5051310889870e96d6d29933bb69d10639e7207ea47c2cbb739e9ee94d14cc471d09a706d58af370b16c215caa3de4459e9f950b1be5382ba32c4d64a9d9df5c15751a88d034021b266404ec213033e6511c37910be2401669604ea4ad92ba52d7f6dae1905f17c61eed11e4d9c196a3306c5b74c5a643df10273c19490b342276f1812da3c9f273333e4d9f07cf11c19a29d7b2bd6baf6c12edf1cbe9db02a6a92d795b2276369068236565d052656fb3c7e45775f6e725c73c376640e144a9d65142895b7247e3961134a9e835891345a0138ac755f1d90219d4987ba3e9ef17799a7f2a3c81986a85e3997ff9aec3c90ca72d83afe57639fff39a261b2949e1530a4ca6bf73a8e5bfd452c619e641c6279fce97d5c31c2c8438c9449bce62742de60a6c5e29a4302a4e20e915451312b10a913790009ad35ed54cb50fa4f32d457ca97092c9286cd5a9d8346dbb70880150ed95b657d61d3c96a15e78769cc4bcbef0d417995758a0245be50e57c1e4ff800cf868507b2c51f3197fba392153a170248bf8bfe5244657340b1781b97b9558138edcf63df8d28e3abab23a08cb1f8ed1c46e18f7853803ab88b3b908a18bf5094bd4adea9b9ec927ec0a8ec89119d132638ef7be7c7bb631adbcdd2a8d18d227a32d5c1f23b73f33ed03feecddf1988bd359382708daa815302ecc076e54ca499fdfd26783d4474e2b9659bebc81563904c86cd1ffc953134bef6f3cba3be1ba8938e5de4e8d2f7c58c255b7abbd53873865b09cd8c3370445dfb895d626fbc454421abe278dc2ec1035f0e1ad1ccb9290aeaa38c4c69fc5f15cb623187a99f494ec2da5734d51b5315990e529c3691ba21102fa8f3024a61bf5a7c07a18134f6eb3ac302b510017d9b3abc3bda8ec6ebc870470d7384e6893dedd08befea724a3640e862848945cd6c7af856c2c36162de5121142cab877299648a5f6c9b45a4f350bd0894994317df970b40417df9d2f339d3304eacf38c009732c7f3cd1e2015d4cd8636fc3e304a20f47303250799ac4196b731ee10c533eccdeff630503be18024cc400becd27be0f682baed5b950061dafe5ca7d9cb7e1b99760253b9a7f5c1668c5864cbb3f2501e03a6a17fbf057f32c85d1adfe9f0f6b17cb20ab18962d30dae0ab003d81a15b12bcd7bf4f1de497ce3dd2cdcd005c303ccc02e2b1862ee88706a67d4337ac1ac02350ff69473bcf037251d77ab8211d2d647c8fb9a477b2fd08e77c6d60a48a532297ecd33f65db157272b006d4c0a43f607f9909c7b6e9d53399bff136e035df27c5d23ce169f06e327f5f08620119b3bfc94e60b968a6dba892c6fac3d83e2cef72d6d0ac66db60539a4aa9b590cc40b890a4f8f06eaf04555769f46aab8999f3da2e37c9ebd344b186aaeb2dbf5ed32afe1e206bfce9094da74b3e30ab5225047fb4c6a0f082a3cd2ef696;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7a59f5255979307e8d06638f512a39b07e2102323d852ac2323e0a69adc937f1b9a743730fbf6d3bc134d890224702ee7e014dbe943ec620740247ec04a475003db1f46949f2bc4fba1be41d4cbede4319e216c7a9ca0e64899442dd034a6ff19f5c2f81935af5a21ee6bb175014a9d6e6783eefd7f7bdb9bb51b47058a1b10995e388fec3d6cda5310f620c27436935d01831378eea429379da21df3dd7479d381b15c8b12d35e0195e38af7a1868a2610f73eede1948dd437e2adc2f644b692f44edb9b6475b8a4bb3f333ab7739589a378faad4403510dbab3961031c6094749eb2c90fa8635b3eb5a258dae17740486e7379aa9cc602c97ba184f434e75b3f4cee9f05e74eebc8768c59ddc1023ec97500f34d075fbb5f54d778f02b4ca98c2be84a94d0ddc62a9f6cb68186263a739a7a593d5e50bee6e2c778e898f58f49579072bfcccd66cf25654adaf62225e33101b90393aab9adb36f3990ce44847c8546a0e68949a722a642fd9eb1364632b95ab610eb1f6ac278e61fb389f1f19b80fc6789e6dc482113e75206419113b1ef5b38ef93795be691015bc799041dbba9fc69bf7d3252f1367e5f7312067da5d6954c19a4f06fbdb555a4452540663c9ff02bf4726ad209afac152de9623bd6a74cccaa129873b493d458bc25a74cb7d9e71cc547ab7c63775cb0516685f5f7da3ce491a6bc014ac7512b8268f06118b141b83afddfcccb2ba7476e9c64ecee626f465f2340fcf6f08abd9639027f4450a282915c572954fd64d856a7a49c1f5f1f9da2c41c6e17c1cabd6a2a2d24aa0d81f4774580cc3c74a63d05331764734523a0c24da5b3114e923d52f4d6f699d096480bb328560ebe13e468395685dc6c110c40d8fda189fc4b8b44be6b3dfbbdc0b2f943c1059bc535ac513ac45a7dc65f2789824cc39bfdb18016e44f16ae628a146574c3e7b77e8a1b23df0f8de787fafa4df4bf3914e1e8a9fd2e1f014e4b03da9db93cf71930b2f351665ae8bb0be068cd3ed5296d60e9018f09f8355c1d87f3c03a2435b3c33637ebc2691d3797a0fd62d6a7984d3e80a3b84ee54a7daed1836cd20ecac72954ec0cc0b3ca67771ad3863711d8e5541aac80e192ef25981f71c44220d3a2371e0867c3495c7e672c3d117a8e9a097043804b0b6e0d8e6d0c60e6fd985f67da115eca01160dfc1d7d83fe2db4be14684cf477fe9e5192ba09f69a12100f59e29fa8bcf6dc10f7a88e6e6ea6367502f1395d2bdb7b9d74eeb6f11c69b87e8e50d9c6c45608b0cc859227b82a7d4426b1453afbf9fe5cb24c70a698d4ea5713047f4933590aca0eb33a4776826d1bbcb5c617e3158612654cb8ad52ada61e7c5c6c0243b24fe1df0b053518f2d3191280ff4d8daed7910ca6eb341fe8577a8291a7cbba3617be565ec8ab76f62b4cf2aed7fc2f219fa908f88edf7bf8d75fcc512675bf14f982e91217a4779a478456f88aec01c6b5b42be44caf5651bf94b27f7bb32e8d7d9b3009a3a1d2bec1dde17bcc85b03aeaee3c3a42c36c4f350af84fb8cc78253ca7453e34c8b82f7008bfe82e4e3fafb606bb2f17324362db8ee0bc10cc05630464cc589ac21ce45d741ae2c63d8ee3a603e84db4e8c298a17c62eeb87d8a9f3185a3b808e1a223a1bdd1d8dbd4febddff276f13fdba2656a947cac30d1cfc9f557896301f7291542bc65f52e492ece5c0d43606da9bebc8e9955686f2a6a34ae6ee8245e74ba103d0b2be7a1af2e0b0e8838d7d5d3d43257f6cccb6f68a1f12d02d9f7c058d97b2033d3d2e44ddb03621f7e505a36a0daa934e2a5ba1da5379040;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8d6d2b44eb2e287cf136ebb5d335c9b38cf2c82b86f14eded6d4714184987b170829ef4edc5c98fe3c6b9a0491c8d04f59694b9aac6ab25a1bfe41b120a69f42685dda9f25dac7c8d421cd74b6f073b7c8e095da989155291a95a906ce14ac532b698128c037a1d2ef8d55f227cc4aa05ab83718c19b811a90c9d10d45f2cd2138f9895c87d13db29ad559abab1cd5afd17599043e6cb5e42d813531654b4a7072581924f97da593160389c71304b338523817c56f65af8a25e7f5d0fd5544a9e166e2bc1f27309ca8dcc57d74e57a140951432cbc48328b8aede92777a1694dff019e67868b9e54006d2323ab982284dbe039496e0916b82871a64842f31fdc9567f41ae64e627cf84d42ab741b4803680608045972e7541a05bb864efba53c4f2c82f618e3eb3f77971f95b700ff8964a7da21b2574ac4f2214902b291728331ee514378dda83c9f7d031c8b8441d86b4cd51cf7bc6c1fec66718e2a8aa9b738dad78ae82e6533da47c5b9e1d3d393ee795ffffd48fc01a735681e292bde67dc73bdafb00496605042e4c58907d2689ca08dfe8ac394f9b8e4d5abb0c8cc666544e6e1c30abcb7857c8f0e4ea48034eff3afd45436ea940ee648c4fbf091ae8bc313876abb383c511ddd8acbe925ad69ab7d9d4fbe9b912d8b9389153b9ce367cede31b0615516f3cc77b8d9cfebf3ca81353eb76fe7ee04b87aaa6e6956fbceaa9988509a6bb655dcd6d3b1f6b0df4159c9d9c85ac835c4e8add7a504ac09906e9340d90a130b8e2d9564c0e9d1d66ddcc94f398dc491f15e6b753f4788f840de7360444831305795c225338f8a3aaf154297021e76a67fd6ce64dbd7a95d5f66c77656d9bba9251ac91aa64e3678c3de42b5a2d9e8baad5f08da0470f6db7c9be1f8328f3255fd1d38b564f32dc0bbc43064c0fcee18d8a4d1be3fe848443983a4fb3f4efb5897e1b4283bf4ecd57833869e7855050fab56c98ac5660adc7dc10c2230b10a7d97555bb13d185534b1ffb60a8b64a51eeb175935c19404ba4556da2f11d59bf44bea3815ce6517fffed34b8e4dfc714b0bccf3496ecda492aa5f68a91b72c1b383347f24083e33101240dc8c99fa9d4ae3a4da455f169d1e36c5bff5da36c67b56b3e660fa86404dc2f7c8c3856f3ddc75722dffb7bf9285b26367c329a7c32507ebc4afb2ce9ab2f7ff88d790b703b6ff6119b05a1f9549adac2d78825a79aae5ee0eb30b7c6567d000669fe26c5125cbdd657c86275e7615d747fd34b051500675ce9644457273e244157d64f9c398741e8d0c7b9af622e57310612af5d9f8b4ab6a002783c59cfc0ed25ba6eb6693ffa183d2ba7df37458af4d6ec1c9360631c443ae00e67a1cb6f0e9743573277201d4ec08480a04b5f8edf29913dde105920e6e1df5b18f8dbd1f035e24262060a8432f8275cecc29ef8ee9ef36d1a790f50c392460f1be98d6a8372296670251aafcfd5cb5ddb2d55ba6ce560963c90f4db8b6f18ce47d7f945f104c3f2b1d18d12c4a7bbf808e067eea56dc6a1063ef4ff90f0b3f7905e096ec8ea956589ac3ef58916dcdc00f0f377fe402b9ca5213a510dfb11a138f76eff33d8e7d75c5bcfd4d8c46cf93f0a9ff9a3bf73281d22957a4aafb47a0986d811eef2ef8900e7c3244f82d8c07493ec142831abcee1fb58101cae2f80832af8307bfe1b3ddaeae207b70c0d22c46dbfe2c9dea77509f62ae1fc0bd30c9af80c321e2cf1b2ea99202f6b1713e196fdf36857ff8504eee6712b8d62e1f8312049de00cd6e5e8e2c608cc176df697d9fb6fe506a82b37f5ae5469a6c20899e333;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4a08ad0461c0c8be1f6f48c9c1f5fcea5c4d0a2b1bf4facf12d74f94616cd84c0b251d0abd90d4b975f0ac67cb3a942cc0d22f787e7fc9bd1f820b0a5365564f3c4b60801430d9ce09b9d7115695759f2f0ddd843e24e250546b3a15543a1de624939ff2160a6d9ef0371bdbf33ae5a111cecdd46c47b3c9d330f891a0d22245e442c2bf257b95ff173e55724effc8c591955f597debcdb01972b9161bece41509ddb516632a7a7168dd1f80e75abe513fdb2016f643feb33714d8aab649ad0a69aa7f4b3e4bab6f617cf44b5b33a0e590e425577ae6f56e88f182e5dc6d7b41625c36b0c32fba4cd098d9266be75af3d70736847ce2b13f9e66df42f4ed89d43f1c6d0e202826356c0eee132023bc451a62df956b99723deb1646db09c4b187d3104a34fbb7b990ae50eb4e8633509ca63b9c05a418b8a719fa69adc8d16a6b8800638d32fc13801f8ea86aaaf37a3e25f25bb868d243b5f9075778422c131b390f49e5b6a0bbc7549001acb2597b79fa8a7a8089e1fee91535dae8ffb61beee71d4dd610ed44f6533b9568a08530738dfe0a1a6cf66ab61066dd39c6e55990b6841b0d3f33120e9541f51b0b8f3c0d349772eab12601f9b2f6e9947110c3a7378d118666d442be49bfed586979e0e37f413962ebf5404c0477b27e3474eaa550725c51ebbf8486545e3d591d9f317d4e4b8604417b922675ae0c041f17251adc9b993fc5edb3ccaaeefd4a713099c605293de65abf1d388ed2d58754515d7e1bcd790ad29d63559667556242f4d11371a2a2eae13a454bc7b161f5b174235aa46b6dbc0282fbf637e0d93f59b6c5545a0ccf74956d0c1162dd080b9ce9908586359697b10f9716458bdb32044d6ebbd2b58df38759ec186a98186ba2d7447983cce2f7fcdc6c07ef6fdb95e907b18f1b9eca7039f48e59b190f4e523de014f9940d4370130551b82a8113cb7506d60a83d0adf558e8d5920ca74672df37be9787ab2bddddb502cd5336e7c5f31ad0eba5f0ca30a722d467a4343dc96eab1b77a864993223268a56865c33d91409ffe871e71541c8ee00093d8663d5239abb33f2581513cbaf596029fce4dde01e974d31ed05acc71e4c995ab4ca749aa541523a374f7a4febd5b1e15fc02c9066c83560d29dc304fdee7a81f5a97fa5b00a3a958839f09b564560694087bceb6349b4426785ecf169f5b29643c880d8e9d280a5f01e5eb55cc4993fd4dfed7eee33c3f68cfb3d10774eecd449cbd4008618152a1f74660244a7ec3e1078b7feaf5f020bc439f2061c2baeb4f829c9d75d2e929ac7c1c1a90650c660cec754bcd3a8c5f92a9f1c4f5dbf179178e2a58b8407266fdbb5661fb9641d28eb3cd09a3331ea7ef0339b8e2fa1bc8f77fd357cf7d42e56c31f137c731d0f6dbd80c8a0725eb3a671e79258b4a773363a9963d9f884917b2bb48a9d27db3d04675c26a1e50df5a8f6cc4e67db55cde41a5faecde156107102d7316f0bf1fabf636dc21aefd247d4ecfb8cb2f6e616a55ac3c5d59f049b38113706e3f3c298284d9df955bcbd63d1348ec76a9f2abca18fdc9a400921878668dad68f6308950ca8243eac01a15e82b83f58c53e5f49b8417d8c72eb0fb708bd8f0d1aa0933c6bbcf99688f675551214cd9c8aa63005db991d62b5c434d12f4d81009b07eb9bc15bd628cd907a234e1ce0eaf341a465ad4ad4278ea4d208910b94f2cc4d8e17008ce8815e928b82b9b407ad6f5ca60e17d331d35671d2f127420db055c4023646010bee6067cb527f91a21d40be328a908f7c1df8e357628b22c03d6b2da7ae4bdb47d45fe0177;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2ed0342fbc0354bbc5bfdf9fd40ea99667bc11d62707f732c300e1b04c22cd9e66fab133a11cfb5146d5509bb478724835dd577708c79f3ac717c967738c31e814ef67b8ae7861ed3d0dae9c258dfa2c755633b130af65e90ca67a8ba7f1dfc2cb9161a34378e98b428b452c5ccd38b6325ecc1b0f7bb008a4259b870df9bee63a125b1cc5a2e41a38cc73513ec945ccb0f097bb08adb1bc0d5312329fb0a81d062436592d13946ac30eb21b34797abfc59849dcee14fec6bc489d31423c9662d22ff29dd569493a5a40c10b5f71b52ae9787cce63dbcdad3db480a3d3c0b006d063382b40163ad3ecbc228088a56962fa6f0a851b66c5f755958bedea8cdee1dbc270ebd1b5d1e1c73cf7e6546f57d6c5c46c930c8014f3a5001e1d8caef57f9f6c410d68c82df32b043dfbb30557993789bb73ea743ab130738831cc5368c379e6b4af3cde8154a81ca8f163c35ef80c78c4a6e8e0377326c2f98eaf5f7afd662833d19a71aba369da3e238cd6d4078b4e6fc8b3265840d53192ea315847e60b16a6ca700890e666b5fdf8a6450d155777f43ce22bc7de7131df61a4115f2b7090d017ad6dd30f6d6c2fd7053cbb1c28ec5ebd461cc9a8d5b91e32e0d72268071dcb9b2b88157024f1accf4c0ee36bcd9d4e51ec9f205844435898a8433561d71e1a6522a3b7de15eb9c555da8f565b9de174a5c30caabea5cc032cc682c3b035fd58c8ce68dbca3f2d366dd74d68e07814ba5a0806de32943b0488d1bf61a12f06debed55e67ebf81687cd4e3bc024bbe8b898ea9f04b3ba1d335dd8346daf58c3deb2ce3889ffe745d6c2b633f84007abd4bef838f29e069238e846edc174c19dd43391a2ab020bb803ee2742dd0cc23c6a1ff1b6e0e3aaf6893cbd7425350820f60367c81269c7d248770a0f7d22354d2e4a2f51298be31bd228c503ab036c458d3e7af6c79dfab48a32161309537da94ca34e90b624ffe645c4351c1d51d781d9813c3bbfe6b716f1dde869774833794b8199c11f0036960c0b7b40106d8c212e4b53ccc6cae1d0cb90a497501db72d3a4fe7b17062cef3211abf21e45775bcbd29acfc7d394e9d858afe3261634b274be1d122e46f256c1e5a86b2554e7c5ca02b0396b9c2478942d778cdc10835947cf73b3b3bd9f4e08ea3524ec9f53c7820b15b0a3c5df64d812e2dc41a77e0c6e4cda691eb65c7ce9d3686ce1c2701b28c4f434005bdfdb1ec78d3ca5efcc45cda64ab89de2aef7b040a29024b4b903a0bdb1ce89afc1ba0d6547340becb252e065c125a7eb79fcdaef6c99132402394639a5fad54b2344cbafa5211d49f20ddcbd97b7e48d6e1dee7f7f2190e9f72ee032a5fb073664a89cd23f3bd557ace60ed0bb038679587806c47a1fcb2bcecd5e7b6db98d52af67df8cef3e2fe80f9027fc527211df61fd4e88f544c12920a493992341d3a245601b7334cda484060e745d1ca57b79d5f943d5fdcd77369a1440f9d4e9e77b1ca8a36d908d9f0aa7567aadf05e5f3d7fe45465e769f7e53debf8695d0432197d3d3bcf480baf04d55a6725b7faec37cd5ca035405045dc8aba3c9ef59180b555d52a2ad7d2f9b389015888e06e6d63394c7f1be92b6f6cfa16e31f5a5e417fe2b08cb00afb6cc3d70af254a9f4696332482d283a64e6ad28eb59d76d57af954d102c45a242d271304a5077f91a42e098d8cb09e4fd839953d72ea5a256e47e9223d2242ffe187f557d00b80846f15bd8c0c9fedd31e3ac8d0cd164a4e5085e101262bd0a6b8081255687b90e51dd1a6563c63aa52fd9e776c05408c8e2564a412c113f7cab29dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h486a589090083cd32b8b40409a8664d6944d05292a5b456e954a3027422c607a65f4c7edafcf4f3b5796ebca55643e483ec946161ff2aed7d1f21a3d5b9a80f8a9229e83031a59b451a78b83a33f21fe265c521b2c92bd380a919982de577a21020f24f1214c3243de16ae622573b73366ca5845282397a1e3b1936ffe1d7181caf41f2f15fc92e3ada7576a2e1da76880cb9dbab45b92da4d6f90f9df6f0231a8165532520d6aa91a18a0b78c9a79215a293e9b90415354d14853f05c59ba625c03a67778ee2bedac8829de5cff53dd24124aa4aacf6808a60546731ed88466a85488410925d97310693ed8438e25e910c86e49deb1fd39a9a4ab11dcb1c6541d8af1352c88acf4c9a28468ddc5333d7993af07f9b75f9ac42def52a4c476348d06164ac975464a211ed98e9a23cc01563abe35a3b9e31db0f5fd91dfdae1b7c5b29334a4dc3a8a316db09ee8306c022def66eb2934cc38fe91102408ad1fda633f85b3cf7518ad352e4fce6bf4f31c87cae92034c1c850ccf83b14f259ffe0228abf8cac0106aecd6f28bb96ad5d682e4e8ed41862ce605c39e3bf8dd24782a70cf8233121b1f7704af839042db39b5063e220bea2b233764ccf524497944c44c48513f689c8753a5adc94e9896f0b51b3120d626214da6d9c12fddd32741fdd48a4f873e7991cc305840ed165860d6e5b2a777f164c5a94cda85f87802a8d96313a4ea570b0546cf507b8fc4e0d7e9ca7a42a3f099d59e6c424c14b829a192d7660e3206b8d3f2961dff0b8c6066dedb121b8e841dfea693392e899c05cea138407daf5ff1ae37011c5ce4f4caf9cac2d1be46695bef4e973e34122237298783299b779513e9c090d8adf62edc121b7982d9b9ed18e0ecd30f05e43c1648832b287662309bb59ffb8c540e96d3c6b3d81cb79b7371ef492ff700a2b8362f2681e729884edae6a4912c798ea1486976125d211883bf7bc136162dc55b2f1324d875369b908d0cba040c19053a00586d2241e9566277be049ebdf5f5a4a47bf21baba7e81326140d87f4e6b663121f8c83fa68b8307e31d8216d9f944a1d363a07d13e2d415c7fcc3d8296cf8c1f227a0ff464827f3857a5cf2fb87599e981220875ed8c96c9a57844b8562dc9a91e39cca21da66a4972b942e9c6c7e218ef4c8e1af40f765d82219d1a76ee51741ced0ff5cd19c0f72f9d3f9a8d6e8ec0dcdcd73b4cc8448da8f523d89f36a2f46b1c330f8bf952d18b159d9fd317d22b5e10eee92fd5e99386846d80f5b81f0153690bb59cf42ba983729e05fdc48d9fc1a28e96458ec2fa75688dd2c739ffbfe71d9803b68e8d6c2604920c5359e75b51707f5afeff282977bbab951c3e89fb1f053d3a84b760029558ccb318d3d17e3f88a1390877b401863006db65f8d9c5aaf717b55fcf1d0ce40b92cae67cd6b2b4ac7424f70d5147d4d653d95d589707d57808aaf27587c2fd7ab728c5b8483614fb3d7af7402bd3db5018d6b2faa46637ec33e701024c72bcb11ce58749f7b512e576f20a92256d3aa6c29b9d49e986134129f127f1e2f390368f4757d0d17a4a29bb65774657363d926e4a77ae776aeacfa9ab6f26709cf31097c034205f7ad16119bebeda32d188ed1fbe0d1beb7001f52dbbc45901ddaf06e13bc3843f29c0210237fad2fde02e4a0044dbdd0c7886b9009962bfb2e0b4e28e16f28f40d8ccf9b389e37ae43dc21d3766ee24e1691f61d3f0597d60d3bebbbd293606424655304d52489712d4607702024523e2a317c959066b9b38e7898f642f555dd89c56f797ae5b6e5cf0f76a35c332e29afc8a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8b47b92bea439e6a5f9fe01972a98e22b46195d2d40836b5d5c09c95366dc88305217bfe809e163dca45a8a83be6eba0a6cb351a098f79d0648b7bb0a11ead5547d1eccb5cfd9e7c19b64a22e2faf0318adcb15058b79add73b4cf27bd088252d242c097d23740e92560087a30233a23293f2a0807322c7ecb3cebaaae03eeccbef4f80e53e1bbf2db9d5a59bc0abfd77137528af08e8e3b4a3bd2580c0947d5419af73d1fe26437a6d24fdaea02150f3911e0fc0fb217deea18c46c91fd9d303109221f5879b286438d9ac39de22fdde365b25c874cef9c482d197907d6e1fcb8a09cd85cc2972ad38e21648bfdf91f6a9a3ded8986e5e2ea0653d2ff43cf529da3e0b9898652252edeb6db54d8eef8c867cde5c473b5bcde4cd1b1e3e36826123558617312001f2152a2aaaac6a97e69064183926e901933f4d045cfe0e3f4564eb2319a8121da39ea14994d9b48cb96725e370dfa40730657c80ede58adf8a6ce364df4dc9c6f3b5b42074477a2076984700fa7ab22c5b475deba46dcf8ee6e542d43671930f03b3cb744a26a694ddb4149051529a793a879200ffa50d22c2f6e7685299fb311ac39ca1b4d338c5e743a70bd107f96dfe13bef0617639335dfadfd4667e12ee51c225d931a8902c5eae2106a2454125fc9ab8cc98110f3d9629f45ef078b0a29c54f876734cebc4da8f8b8059595e15c1d488359c71ee8addfc96419fff660c94142b8114caffa536a614a2cc545f8d649f8f160adc8f773c315bfefc1f5bc37f6abad2f54db6ddbef044c8f774c4ec5cb0f6f5b8b07a63c685ce0eda08378d7c3652858f7e433bccc829a994675044f253fa1df30488d4745260d6fcefd10bb6309cfc31ccdc8a91016fb179f7df30587beef6580ee3165bb2ee11a8e5f6aaca4858b6816552f0684321c4fd1f643b0a9c116c26d95fb1da4cb1eafbd09a3f4ba65f8eeaaed363bf1841054204bbfa64575e8a08240dbffaa625f1f547af5e9ed22a1ab39e4454143a73b7ce1e4cd978f320fe6521f31d7a027083b60013adac315c237ed19d38b3af8fa01d62f31b3d8f0a871f1a5298341e5ed72925c674b0609f531dad77e888f366e91a8c7ab93dc214dae0c59c8ca2a34ac6360029bcd72668d588a0317dfe5841567a16c70148ff5bf10f07410ac57710d6283a50eccb77f1ab775d3c4539a1639db5af86fc475f5a439be3097893641fbd7f07d521c22d909a44ca2addd0fd202b8a175df0e64d6ddab44d5f7dcddb58b00140521295a70dfa0789d740bffca532edf130ba1138a68739e12b751c405c151fd1050433fe62ee5a753c45e8debf130d4bc23f852e2ab2623273890224b91ebf453564a288b7a4c690971655006274705cc6e5661bb0ad9c6f582ad314f0e84b623c1148f465be8f9dd6af00b7ba67462ebbeaa53351f98d248fec11d1602475c22c578bf47fc561297ca84775eda587e306ed49334363fc4c938ba3bcb0b0df81317cbccac061a25820e902da6df537732f31773b80589fcdac2ae743372cf148158a26e608aa3ac4706bb8f03ebd8d149672e5397d6c856d2ea173ad578a27daff6407683268b157f415f8eaac9494e193fe7df9a85fe17ea72bafa61bfd4104d17cb48051a9552c45ac4e0198984812e4c896056020f27da4817c02c5cda709d262f0c6f0d7add48d448fd6df147dc59023e36713ef8496ef0f7c3f28e177c8c424dbed3cf12e43a1e89f332299199462c87f3dcd98cb58b612190d5c9ce5b2590dfa885576eff100c652109fa4756fc3fc488c9d5076bb9b2c0831360cdab34a96bab0c954c0d88a01c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he124ae2a5a0fe99b82407de414c38748812107cf9959d8e6d4da911b76bcbf406df65f473ef6ff44de6f0f4c498e102649871b423363e2332a1a6a088793d4f44a1998a2fda410066b1e7f87f0891c27065e2cf9f52a3c006168c480287a3a1416f8a02bde2065d9a0e239ba0c12a0c05f640ef27be5fe8d27e76679512cddfb9307d2e0914d0adc541ba579b411e2a08455149f91052bc0a74f19601bd60bf99cc3cbe8785fd1fea68e5b2807a02194da9965820556df43d68a83ad35cfd288f1ee6b9f6e0dd86da92a56cff264fb52e02d42e47d0140c4853a4d586cd3a5f6880b4739515b6efd1ed3ebdadcca1cde14cc933f8161a00974bd32ccc074c06d45316c3bab9c0c5490d964862d54a2ce031dd03197d5ac9d1eca607cc6e14ca7d228c4f4cde462d44e16fe940d2d01ca5462317a3401cf2d1597e2c868bc9b5ce5693e8b056cc26cb629e95dfd215cb8d9eaff242dfcfb5eca5919131e5c827eb5ec4911acd4cf911dadcd181b2226da0cef81c907dc09139dfbdc7ae879021de464ec7915c60fa58f3c01c718ecf89b01e0b0bcafd1ee383360fddd1b06b9e490978730e0301d61af5d5918374ad6f29ebbfdcc026eddf1ad08fe235afcf5a5cb0a18811883fa0c5554bd286d3a426960978117051c6caec178261fa6f81a780405001de5395b80701a3e1d3a06b07678df59d8378c0bb34409cdd7402f8a2c5a9e71851e472039ed02864b7bd5a60b20dccc046e80fce228f93d696e7fd602fea86c3df06b9da890d2b50d954cd830828bc59923fc1b69a6706abff8ef5924b1de6174f8314026b79affd55bd63551626a9da5c5a29b7c94462330779834d33b4efbe48efcdc6096c800c30fe18d4c66214ae55161283433f2d520248f6b8d94908ed6f1d580a1e04787476d394127294088e6865f4113219f232344d6c2b15f3196e94df006ca04322c037323848d7617fc82cd2f9d76ba85a9e70efe06e9d4b6c45052018057481f633c29d5dda6ba20534cec4988db54878bdb132bce73926b258dff1f4f33499e1bc2177ad05d02662fbea88133a696b30e89830b41a2df6a155f462c325a6d917caf1fe5a2e48a9d795c3f131d6e1a9f08be89c1fb334b7d92e8d0cd4239885e30b5eadab3ef87206f7d637d53c7dad3adcee18a3f72fb01a20c28a0b23d1107d57f2c0ce8e20e65d8ed8e71118fdda14ae764045807e936a6081a2c25853a7109510b8854674ac045dfb2cdb1a1e5a887a758b25b55ce6a0dd63e26eeaf98258ca50516fd1fe340278cf9c981087f789a7b148f375fa1678ebf35e1eee08d3623dcac56b6fcb6028f7a74fc8f4fb545cab6560512df72646493d72eff782d6c38c06d105e077a0c607c192c6e00b636f13c2a1fb13376021414cff6ba2af426f01900aa6ef17b81408ed959aa41cd6242110a7fdc09f77e4806a3ff32e4950a29bd5fc13a52217cbfa88c36f0bb2b1b37d41e78c8a8144b14e4df2aa8e87177822d3f6517eebfcd728539cd83a0063d992b007665441d7eb1d37360b7534221724dca46f48fa35fa8378af06b7788fca937154da368ea31121f0dd6e3bad8576e9c2130b83934d71815d7bcff0c0235e690a46371ab688b23046411596a396665981242e0a2ec4af23c297f8874b9c5ff91a1ea306c3dadaf3b14c7231c1f0c6d170d2c1774efc1ecbb4471eb6c9b6c39f82d106445bfdca609a5ad0453f1703c0923c0c14e450ab0584960b72d6d4e0977902f5b002b8793465a9fb7e1ebb115556a8cc8213997e8ea3dcb6280975fddcbf70087e237042dca5d30cfc7007a087e28bd19c9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h47bc8adcd09b996f8c1a31c6e897f9465a93c90d50efc15af20fd169afd2dc212fad97c2cb22d38323ac0537af9cfd01c39372f1af097620c6788559abcd2e5ff838a41947cd512e4dc5fc84b1e0d0b4c5712bd4e7c765ec8a8c5683529ea622df68e161088dd0dd6aa90452ed20ace036c7a31f19071d3fee0ce826d07fe8c24f35ee19be402774e9cb0a229a585de3c1ba59360fd67fef10a37d36fff0db0e39cb6a91788b493c2f23f81dba4de84af1da2b76d0df953b7f89c34084a5c700bb5e6e039c218bbc9cf30cdcf713c8ff109d9281eb90f37daea0888652bb4f586f8d5a599cb1b52d872fe5a0536aeebc7f664e13c385c23e1bc0e1e7bd3fbbfaad97934450aebeff48ec879697ed8f9f38b76af9052c612a88dc34cdf632dc2d8ad92ce00292c804737f84e7733d37c6db61d84e39ec23ebeb240188309b5413207aabdacef98d79f1e1ca6121db6b881240ef4b7a1ef095aa435f1749f4b5f6d1b958b5e7c2bc1fe1a6c57a2f8c15bd692260a8f0a3425da9110a0e42dc6d0a0c6e5573b254f6211d9a911c20b732a9e32d626602340d683e53190422777f5c1d16ecc7a9a9d6a6602b1174a424d895ec5ec8dfe4d25444823d71955a8ddbd77277f62a655c7cb74fa8660b91d1d7bbdd10ac75ee07ef044210d3f8a046dc780b316181c4b0ff28ab5347c522e7751f96cb0bfe649f56251caa81856e9c5f5de6511390d678e3283bba24dbf70eb8e71edb1062080b2e8d85515721b21f0d85aa7526c6c9d27ed0b7c799e63aada6ea6fb9064a8dcae4076928d82f93d56a9fd04b6ba5986b61bcbe1c68a9948b8ef5dd38b7e741aea822adf556a1e3af1676ed3270abf2ebe3c44cdfbf4832111efa8ebcc314174d29b18ad06fcf291498caecc2c4eb09759cd43ef8d89bd18a2f6ef2a031d60a1405372df0191df35e30c01eb8449bd0ffe980201e9cb3d2883cbc3359bb20e94b6d05aba7da2afc46b29a3ecc9ded45b855e19a0efa2956b743edc4f55de2707e6eeb0d0b277e531f89843dbdd4eacf2f6bec2188011c60b88b1f1eb61680f1b399b37fc253bc57e4c6b845691dc2fa50eb7d55dae1a378092ea00db56fba34f412146b927516c65f4a536f34037af7130c369418798820beed6242ed37659e5ded2be94ab7d860aa403c5ed573a47135744ebef233a10e8eb3f53beb805a93583454de397c63f5ed044cc52db9224ce6175fa77bf1e32a059a9ab8151b9dbbcfb16cf77997c004f64fc1b8d5e3e06ba3b37aed6ad8de985a767c521f037f26fa6dcf6de81ad29c875755ad15a10369fe2b9336a183f3b1606596fd03adadd27b67371f7da22a5ed57bb77a7f9ec8737a1c2638b984070a67a0d8332427a412c9eb5eaf677d327bd888195b30365ca0418926f194119a86b9f38fce038ed4e8599897ee550a851ae1c6d3f338540a875efa07ac8e25fd2408f2c70d9c70d5c6dc495012e8841b32c2d49de20ecd32856abd6f39e906d9f6a0b6fe18f895ae905e694a20fdd7bde853436312c0c71c774ba57bf649948c6a0b0a7388440101af91cdc8aefd1c47591e48c01d19a69e26a75f2c76ccf759eddd42becd77a3d5c9bffedc39d6f20a7cabd86756ead7d366cb7077556d7bababa08000b47ac61a3484df0a7595a024390ad5221a9b5f428e013844ad6f2a68088566fcdeb9508050463f14b46b54e17ab9bd065a55d14e14d1d819396127937dd97270ef2463cc3ac5c200a08d40c9a01f764937840c445e0adbbae92c028f8f35bb7e9369bb4d7837526f3a5bd3b367887c9beae3c895d4f5057ab080512fb8a6e4f5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7711844d54e5c6e66f66f53f262bc6cfc2fab452a1636b5ccc80d43932ee6322152c634127936f138039bef121c5179e89b8448b55215dc809c6a467b855c4a8ea9b7c45e1d8ebf56f6c2117bd8ba052870a6d2a60d2c3ea9313abf353532b4b3d074173180515232b87503400247807b4225da109a37be1c3279edaed4ccccd2e8f1b8399875f969c82ee86c1b2ff274c64aa69f9558772486ef571b29b24b73aad98bf530d3cda68b0ef2a83ca052eba199795ef7fb39f0911191e3e2075984992a287b6a162c4c41d1fe814333e82f1e610908068d60d0f6c74cb36d43c0e62b4a491ceed50cac66682370c5745bc0a2f98449a3d8261654cc3f6a8143d52ce178c6f62c8561104a06d44e76a53256fd4d1d544bfdd992d82562f23e9e8d9e3fe5b3eca3e1d02b19af7167bbdd80d437fe03c02c83e98c8381739a8745315c5a0c3c7f3f436aec3061242bbc5fc741d6134ea6fa7b51e2881de3fb3c25b12db627fd88bf6499c7d9a4608a5fbf360f3940bab2792e5a6e69817483e73417e797f35b2742ebbe1773da04282b5b059b873e19e0825e37fd5278d8ae8b4da4dc64a6d5b21cac4201dc4ac3e21fbb2c49096edb46ad2d32ad800ae5a1bfc6a038ba36751532fe7b7b7c7dda637a2020cdd2f40d3e4c593faa5e60c426d5767d4d15efb3ae92ce7ea50d1200e17f28cc9dcb8a38a198ff50d10905274df5094abe3e6853b5769a033b8a9d656b95df0c56c5ccd3ad6a30fa79db0c3e0c52bc6251f4d5d7e9f6f371e85c875ee9127a63a521da89c5734b89d45b9f6020f24a49efee656040d7a9f62654f08dde52059b3bfa07aa09f9866c5e1d3e9467675aeec8335c3eed010c3162e58af8a3182b77e13fe8745d1316af9704f5240ee614f48af6c629fa08f79f3883c8b4fbc80b5dd8a0144791b849096f967591f543957441ba587065e440d7f781efdc37791e851b12de76bbbd6e0c98537ce53168cdb4ec3dccdfac812ee74386c04b3d69050223f89363888d6b228d69fe4d767520dbc696333fdce2468f7d4db3ba8a665044fb0414151c256953d142cd85cd03aa43161690c1ccd9584386d1b98004b8c8611672d55d1593dbe22a31b21eeee833290a1942cbc604aa97e4197d55235e9d91d53ae1c81bbc4eab0bd2e0d35951838f145ae228d89cd742aed2ee68c9f31e0989d226ff6a30a2c0b522cbfd8e7077f374d2677ea91d8f02b378bdcad94d7d1847c99193e1fb2e6adc1402f1c7f3ee0e439292808498d3776619c68a89672504c129a7057f96b2aab88044ccf28396edf9fb0087565699c27a232158a2dfea95032249d7de5a8aad76cb9eed9989ccc3766623af6612df7cfbf717a340e36680c8e93e5f7819790a265ddfdbf43130eb7da8d76c82bcb5593ae78bde21f0c16b64bd951ba83a52295e409c57b4118f6fb2d69996a48fc5afa9da27f3e70bdf45327ca0e0b0d38a80c97888b0ea54bc195ed52ec33b1fac7f07cfdae72e6006579890d1ba0f16a9c243c7a2785af246d4a2faa5b5b855e34fabf003623a5cdac11347bda490e0f35af3fca3270b63bacc16c03f160b02420d34a858cc141278bf0b9e369789da92e7e866ea5c8dc5283018e7afe4cf761378d739dae4be263ae465e4088cda3fc31148d8b57749ca41690c33fbf444eb023c21ca43c58afc3892cd76dadbaed85babb5f2e37cf8833d1834b0027a9b77b35cf274bd9041493afba52772169df1488882a7b554ddbed483e91ef7efb765c3c12420c0ac74009f7e0bc5ac3c3fb50674b9e341a4ff79705a18fc37ee1b7a21e78e69136e34487798d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h48b2192af84f7478f2ecbf075c05b886d20331a11234a55ab6fd65f717b986c2a6f9958e7e7916eb27768cdef7f463558154ed22240efd15be3cedff270cca09b2c2554000600335010040d2fc6021e476f54a08bb49efa90b5248e2c09fcf46a68c3eb329be6b9e9b151747f19fde373f543e78016849ccd23afe8fb9f16b49a967087ad6a22738b2b7fc6c97bdd8ca6ad0c188d5a51841ebd0609c6bc8d73464166d239e42eee4f049db6e65cd132849fb40631d7a92531e46ed1a482df6d5cc96d4107fc902f861c1e221be42614f2dea03b721105e142159f08e8f5537718880e36a4889d54e2833b8edff1b15cbcadb54fdf7a64e53cbf629da3d1b7ea3d09539decc69d10721743e8af34f0b3ed55bb685f00984b3035f30b9efdfc69784cbd9cb516bd42dbeb207219971a15d043a48f5e021835127b53493c4b0c716c781a4b01b8765158f132a5e2ff3acfa713264efe97e99c2815f36b7fa25ea393f99b5df2f01dc7cabb90e77044b8b4f1c83f440501b4b70dee7250184c1fc71c725405800e6fa8079dbc66467ef8030180275a399d0a32339b7cdb798365269c8e29673803251700d4924b05e0f578677eb62d4626dd64c2f6b5af15164808f4dddda24d3fae71c5845fc43109ae1eadaf1b9c32717ac78a853c65c43a7599875fad2e998b38c4e1632fdef50a3519d01d37993953e289f143affd952f0eab679f6e37ac338b785e44493ebb92856ad295eea0d81a7d1c4b4d69acce1deedc359345d48abbfc166a62ecec8b798822863020fc984cbae522479b5412a961e3ba014cf9e7bdc625421c3d5064f7ba88bbd7f7f74ddaeeba802aa3371fd9cef3950ca5f319100c1a673956bf06ecc02366856a9ff0ca0281fc998e16509c8e1a194e7012b95ae92d8b0d8c04092029985412f0aba2acef37dc73d72d56d50c2bcbcae8997e9f21ee8ac0a25558afa8cd2c25d38fca85b4a695e9e84c0064b9be7d9b3122b9a4fa875e98d4da2c59012ae9f4c9749c15d0f1e7b67031bc471877ef9eafddabd601291f18ed38d2d7d5c5b5cbe7314fd8171b52c243bd78921d07b84331f476615ba77772e81b0e22e1a6cfa5e7e306dd78faaf8702b30dc0940824c2a083ceef8187ef815dde2973ced3999c66650f2a482a11bb8d0b83da327a6fa66f94db8a4f33c021ec72c360814e77a643b40a7e8fa1bc201f210f20bba526ea7a273e198fda3afb2963790f1d5ec5d3e5144b65148e858307a7adf5a6fa1576734440e01128b6ad1238df83f70f58b80d8d6547f23bbdcc8e201bf7d251e1c2e249c23a0b4949aed3d3baa687bbcd9a951e1d63a0f665e931ef88c586da5351adb1f6fa9931bfd7284b64f7e6fe05ad8bb4f20141ee8a2819655afc390f3e30fc399c72d1f5c31135e493794f568124d51985071cac8828a9b3f17ec5d30de87e58dfe84634291151a0627d01e1cb559fd43127ea7d2437bde7e39ec7bfc776937049651a9cb6b2dfd3f0fa4f38fffdb7540317c133dd87887f4f7d093a19560497ad9b28236870adb683ea725ba57bfa2be248f297d0a8032af00a0c9f442f32b8f408f00355cf4338dd87cde98a7ec1d5e24d8a598ebd490e81e7055a5da2c4862d3cd38b12d077a1ceed35655763901ef39af98f42934f3aa71cb2fedfa20bd3a23075f4119ad4342adde07ae8332ecdfc223f4442970cdec1fee65ff69d3fad3135fc5eebbe9d6f4c9d0f9efc9bafb5b808aa8ec2f112a95b540980b229c9b6d2b5b626b9c6efa4558499295cbb481436c7994a59292098c7895c2d4fac79bb87fa525ee7111ac1563bda2a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h1e72041e0c67eaa60f21a580e5d390db8fa2fcb0ec5f2e5282f4b982e9cdb1bb7fc89aa508aec51408987897746db76e78bbae641939647c53cbcf84a65eb871e957fc9a44c3e3d6c0b80463ae8e0cc7b08b9656e3aee06aa944281c181b87497f92f54cb6feb7c52ba1de764a58ed80b87cbbd63f1af5504ad908f707286dd923aa17d3b356563db55ece92d9cd1ab72058987fba21b7a61c7770063bf6e8dc6f76e0d8237edf85e4f6c5f4977631c355acd608469ffbd5b5f8b705da96c8db6af5d5e706d739f464ef6ef1ba3a88aca8c60e53df9948eeb82a29cdff001612d1db57ebe295281ede7d99fc10c59572174f6435f103a9af38f54f6d6d6ed3cfc3045344cde15517200fe2a58d8534beb56b1b398270b59bf54eee76cdcd21b692432bc4ebc36889a13d7dff86e33a133a9078ede501c3973e05cb252ec27476212304aab40c14a6bae4c79352d73b1e8a8c90c21b3d25016a9f2102848bc025ddf67301d3ac8f29f80919299b9429a1888d15b5da47b49264bd02a4c8c0456a4cd57ceb8e8967a00bc0132e3e46934907a44065e6329bb8b2bc745bfccc60c0e72495a9bb9284a7bf43d4f2478f08830975917e5bb59e0565564b254b6caf8fa1f11f1a8b3e72f5dec70bb5795b9971a515510436fc94471c54877760ac1e8d3a978bd43c83b7b403647985d6e3e26fe1d1a01ed1743788ce3daad134746d1939bdb78281c1c098e1944ccca161be841c90ea9902ed0f7f49559a6a7c370f0ba7889b1be4ca8539ea8eb31313f02d2a2a119243595f559ba770903223574b01f0b63513bccacbeb68beee84a02317ad56f9a9bbb9c9c23230065eea8245e0a2a42adf820ee269a9733f6c6ec26288c9f2a3c2ebaa6b52fa7744b50878bcdef5dfaca012568bd435133794dedefb67cab03e389f2f31d9927a63558ad545af9b58d55ced747aea49e72ea4b7fe1613de9142534339a875e04e0832913f51c616c323b271d6a2482bea596ed7f33ffcde35ac70676ec0b23b62b567779ac7d79f32b46cbda18b947566740fa624e12a71a24f7895ac5dce7fdc41313345d4a8f821e7c81285082e6a120639a2a82569632fac2175dbffdc0e7d24bae86eaffeadb041a4f0a91499e8208a4fbf20497c4eff23623db53ccfbece402023a1ad56aba27bf625405c634ea6f3115a25b48b11a720df38e8271ec68ddbc866b3eadaf2c98f834dc90bac336b62e95587d27c6963993bccbf807d2290aaeb78d40a931bf887cc459b88044a631da7065c3b0b115b26fd5a9956c2d473d4b3752f1edb4796a6d5a7525ba17382ce27a76e4f63431a18e0b45fea64916af3c52e73b89d05f6ed71e4004a3748294422a9489fefc7d431d12027acd8b87ef4b3c4add71adcaf65d4296897aaac6d9226e8bdb9fce7bcd5ada35b82e5116b04a03fe3b6a67cd23b2f2edc35a1567a9a99cd396c54acbae9783d4653c666efaee31c5bfc6f1637816dc0d318acbf3e7c92c7b8d3a436a056491679e9df014f39eec8f4dd6ff2a076ed45e2d3f0ee124cbc07ada2b0195d2cf9bcc82802cab65613530ceb831954232824426684580661a971c1e0d02d37c4b854d840dfe2810d35acd9e8e43d7af28ba34ac5d3609fe6df9ba64cb2251d91ce4a9c25c7d999be700aed5a2c558521a054f4cf9adaec5dc1c4bc800bb9a81864e0e239d1c15a40b44971846addcee7e41712746a72e345f0b31d0d09c3e9413b6fd99256e06a214016ae3734b39f6ad3df4bbf76eac8aa752c32070c36431d722f23445a244a304525ad14f49a3eeb573d2a2d1f09155b7a10fbcbfcb7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h58f80958977f02dc6ded7829e15b94ce65d35665c105c133d78351ce2292dad3d259e395f08daec5ecf17a0a73e6fa6d03fbda0158bf540e830cd5482a223c2ea612667096c32325e523601214773af547b9fd2c7f81932073c235057547d98a8acab6e8808ec433e1fd3883e905b8801f10776c9f2bd2bb688241b5f9dfbd5db502b5447fc7d9437e6ece58fc52df3588b04754a72c9ceb86406929f7a8a1ef6977cd01640ec68e4668b8a89281e69f7e748ce899f21a99db63b95d05367eaf0c82de33e3e0a1d7d425874c603ddbcff721ac96fc96fff86740419f94f3376ee45db90309c1f4e1087406eafa905df1018bcb6aa47343da493402e6eb5eedb25d3e6d563fad0eb94297be4c5f803d7e59a3027e200bf5e12548725615b57135cddb56aa44a3cc62d480f23ca74b7b9fab491ec92c761a5eacf57f2365cc4687f3f682931feefb2f0a8ff7142f471ddc4f0dd8d54e07b383b105157bc9e744e8d198761e37e4c818ebe6dd3afef0bb4007175646ee6266b3d453d30f809c7b2f91267c5ff870d7570dacd213831af1295d30a22c551b37f6bea67d4df91d210fb16cfd43517733efc7b1fc96552c8e802d60641f76f908950b20853b42a9eed2bca012915a027a4feaf85003a67489787f168e58f146c3d3647fc3ac744ab16ab3c85e719f8d329da5be17fe352e87a22040904716c28c2b6913206f54cdb7e9a1def1a42a4726abd936d5c32514207cffe6ba7301c5c7b2e1fb346f9445c867cc9b83621c75481fd5a73c3aab67d0968cf81fe8a015933349bfa1dcbad8407385eefd488caa77b0073463cd652949e3579bf642cb05c1a45dfe736bc9f2bb384fe94bd8dfcaa3fe3c812368c42ed1778124ab4fef0693f6ac0b054fa9cc1a41ef5b2c3be2e24a9102c9f86206f46a302011797bd50c6525bfec15008e82a22da2ea598b480d51b079fc6c6ff84ddef046a491e3b150796edb4b635c1f43a7e68b2b640bc481dae6a8be8e979c4e0156b601f6f75a5215d21d02e24303594f89c019737f1fba7055789d739b24abcaa0a8e72bba7a01e5ee3de05ff744c4300f3120b17b33095689e8a1cd6d8b8b937117f7aea43e33c0f891ac7d35b8d3189d039c213a8fec3acaceaf425097da7554f8d867b47e66dc6e8cc551329840c6e7721eff8246f1593bee6345772b071c5fb2e402acb25f08f0e9cabc4cc817ffa7180fe6ade127eaa94fe02b41efcfc715345e36cb9d8137c3da066a36bbea09aadd20d79c1a71978b30ea9213e20d3d8d52ab3837772f63482b7cf6c395a0c42e7bc3b7aad0dccb5e65ea13aace68f67348bbdb2cff7cdd1f2d34bacb1629620ca00dbe68825c145bb42486a1c42bb8475e93f37efd42c8d562951c19784d25d54b1d159761b76436572dc2e161af6c699cb2d72935018d1882c4c33124fcc0889993103130a8caa8b82f43c47abc7d49b75d1f73df0d86ad3fcbd8b884959f4b10c9554390d651bf4e1547257bb77428e01c57b1fe9ea7e6806cc5ca08dc51b14620d342ada5ee5ee64b5303c758558c2b5ba39f0d4ed538117e9acbb1b8ec8dd29ceefcad1b4902da52eb2b701fc4d84f208d7052ae02954bdb127fb71536f077da82dbd97e54dfa04a8f039ada0cf1195ad849d4ccc08a780ffd161877f86f01ea93bdc0a191eab89c964706fd5893b8b657d310a374c2f947df3140275d3b2ee9d19c390801cd98f0a6305ab7820eb91a80b18671b442808017eaec2b74818bd4b84fc61fb0dc73a1a30a54d8c479fe1ddb8737497e12b243d8ee62a6c5ddf6a6bc51eaf40289c8f9cac766676acc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hdf0c55cfc55ea68e7e3a43f9fd1da98cbe68c37b76c0f78c0e87dda5599c083b74a143d6c933ec172f380ef27b2afb4d1db1010a741bb2e40af6df6cf0a2d4c0fb7909a1b17ecad086a4723173580c85a2e2f20acd3f668611267e4b61f62f0b122a46e48d6dacd77f571cb89a3d45a192a29d3b57199819e8d8eee9d2847c4791d06a3e793ab8d7a90d1504e22a7e667320ddf59ecb308d48e0f8a5997d852a3ad6e6f5971db8175aa3970ad30ddd34544f2ed54fbc19816eb8873eb4b0ae16a2955c060724b3f2f43691ea1808712bb8f9927b1006d3f735d2a3e40027f384365b06fdf1c9cdde2c1779bfc2abcde7ff38f1a3d5051cfdcedf41375010da0de933dc32ccea9f96bca53dfab0418ebd6a047a3b931405793acb1e1ce3b7db524c588e3fa72255a0bb62480d33f6765ee62fa8d8a4cc15eb0b96d065926f8b9291f593942df5ab3235cb94c6462bf7705e8b571aada7d410d3145f6558172a97cb399e84672e69ae31727d6a7fc8dd0c11798c143319e139316772f308ff7aecf7ec878e4f408648345e580a40fbef9e5ef2b7fb5f504688b46839b070c5f4f673f1490accb3c244e34d9b007fbe145088ebf901597adddf4da28e52d9cc554c9eae0fcdd42cc8272981b9f0d9d212fbbaafd5d659758a00b3c2a6c70c32ce521b55ace36c481878668f06b2e67f685ee155527dbc497157cd091762c6d6b577eea18d3fa51ab132a712938892a6367e628421f62ddcaa01bf710f21fa89403213fc9f5eee5204b0cafe97516592721ac6d2e88e8199c5f4f11ebc1d2d0960de2e8d73ccbcc85614e5ae3d10fb9c11bb8f7de9676c0fa9b4034fe603b049781443b18accedb02d9b7ed7834536ef24bf9919840cfeb09c091f9420543c7aaa7e8ade91b74ead0f3020fe0ce9d4dedc02a74e9c0227ab26f2860a60d3b3a515bf64a3b297dd6291f4f01e1a84ccb2b219c6e37119556739b3b55a4b146554e61ca457e19c5e652973d5121c8048068b6de0fc320fe6c4b72525861f9c351f2fe9cbd382806e37c6d5e76415aa8fd89908300638902677f7eaeb2b79dc46b1e6300e2f124fa7f636ccbfff9cd162c49b8ac24156ac7bf521d9922e2719869ad856fafbc28d97d70d0f238bea8c5b1993a79c4cac8e6f8a23b0d736a3b07106b665b4aafd663de5a50f7982544706e78a68b20f3ea6493fde0a1300cf4590abbf2eef18ac9d9442ae8d3fcb0a7105b02be3f76a32d39f352c8df61fe42497e3d952a29b35e314e2f6d813cb0dbf7e8bdeb401b5a0bc4b64952b01e0e41055e10161991232151629cdb1c54a6897cb5a5e4a6788bba28e72a08e6886a555927dae3ef0848abc1b1774f1e3a51aaa2e8403b5b607a7ccd357fa5de23824cf8e7f1b68b4c77ad3e5346846276bcfe11c6324939bec7decec638e87027cacfbe615fdc1764800d3edd366ce21ba3cd7b7b4b6f7120bf74a69901c46453152519a42011ad7a7598284d4dee3e1c5c1a1f6a0a8837ab5d0133a0dbb15244f22d5029355d803dd6831b20273ce5eed31d34159140cb8ee826753692e4286a248da7b7fcb707a6a30cda0126c94e728adfb4f76ee0596b4e1e1a96de1c333225234fe5581c19ca7b39ee575b3aec1c4a61b9df7e22d137859d6842a915bcd4ca1d671725893d8603afe8e2a748cea8c1f47a536eb0cc23ee4ad4dd6c68147150195ac4820f09bd3e3c53519fbb86c249f96661d5846db5c21a5e0f162f6578316d41cdfd7673c602706d7df5e3cf8d4d17d5f97a8e90a2c97da17c5d5764ff6c4564ab267a322c588cb1735d10020c919b8d02a08f6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2262a09c0bedae53f983f639e02855b8f5fea21324434e152466fc4b1b4eb3572ecacf04ec3fe3a6ea9d5ec2cfd21d4f9b1366d4c405f9d7e0a16048c676c0b44af0e9a511e4fe7d9b378c45d9ed40f2346d4fb6ef365c61aa91207521b84bdbad00d5f0dc28e17f77692b2e6d530822af92617c2110dc36258b0365317d2201b821088bbc5b0c45bcebcd4ecdb5ae225a5707e2b92d9f6c14ec8df86ef975a451c6dc714c7b88720f8b529f0cb387778c782dff419bb27cfe6765b234088a1a5b9507c19c7fa1f66b9695f3b7e3b569d6221f751cab417f08cd6ea92d6eacd3fe6380f14e5feb6c5ea20b7532f905957a3a78f1e307b70cf50aba838d19edc6299754794a1735bbc498e10497961305d715f9856670da5f23ab0f5db210ce879a8fcde22a627be3cf4481468e6200aea7955c2fb24ebbcd57f2c5a0d9cc42f882519ec463f132121ca76be3069ea2e0c2b260886ead1d35c79b1cd8b3ade9a92bebf7b89e47874010275b9ef36aef64751cf265b7712dc5e320cdba6b7367174aeb57134c8dcd37e3658d7614969da788315d9e71c9f6b57e3d2f0181f53a0dfa34c5a0b1580426f8b90b0263782956a5b274a8a104696a685a03fbc478391538c797ca75137d3ae79318122ec045e92494fedd960f866d7072a0d31efe408b1527a247fdc051cda8106c1c0c93c3e20183eca950c0ae4a5e8febd748371e0ae0cddd4f7e106e60cc17569384b2b15ecdfe6bccbb42244242614083a2f5327d8f6dff0f9f8823446268b165f3afe711f6e028b4f3c01ff792f26a807c36e6f27ef5b2acf371d43f18ca7902eb23d2d1d31c8301e1fb09d1c4e85bdd197ce05a5fd5470baf0f1f7d3032e5d5b96ff5e447572567ef7cd29b7f6ee9ed0ba9ea5434b7da1c9de0c5c427971ccc576fa608b40530b4d4f05e55e8860a713a3b75955d5f52066c33c67c358d64e2daabc4d3ac970bd02e8def56ea9fd627da1f56069b0ca43d2e4104d73c5d02e6785493eec0ac5009e8e382c42d5eb8ca1f65cd820fd3031785a9d2dd9ec0632f2cd27d7ac1ea270e5c99bb6c61e25b29bb978073d0509eb9414ef91df593adc9df76f5e743c6b7d50bcf1d954d13c410452f10b684e9c4c56c99b9fe4ea5260eef2ad7ac0da41a48657cc24a6453b00b2ee6d5489e39c0b6e46c34f19cdcf736de7f31ee6d4dd795bb489e67505292752ad924663914beeaa38e2077f5d6f7206f8979b61dbc598bc63d72bd8f11e87d98400b3a093d07c82f0c1977a012196b877cd134b2fe97a84b28c10f677194303021ca6ae1d6097f840d444e7b9a768b17e0a793915151e4423d3d3d730021c3792b23bc98b55e13d148914e4358de35d0feb29a9e32a17d5531eed2bc9c5b2912a6b23abd8e1e43829495ffa7dd3ea920d0e41a514d92f35fefdc52bf57a8de424c23ef98ec3af7365f9fae6a82232ca43355ded65115b83eda7bda0eb64ae878d49697dbcf71ad689de752b1653633bf527988305bb5976233fd008765e92aea5bda1ec506da3981898ed011c9cb6ef9942a46a54813ed78872e6848253ca2e20ce29bf291d8dcdcd4d682a3dd5258de2485f7175d9ac9a8e0d15bcc10fedeb8bc48d4cd28ba70ff7dc94980f4606de17343f0baf4d0fa368859951f617b8bf2780804edba40d0e788895aab648b0469d893305867d1fc83a78ac9dbb3a78962dc32bac0999958edbb1492813143498a050fc24bd3fec05a61e728a05ed6e451942aeb5fac6b30583af7aa385396d95818d97bf669fb4a7e48fd94020c3a229d030a225fac49109b7781dd43a455b4566eb6a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7abb069f3e705cc84f8f7344ab954e0d5b628f0ae4b4b6c3e7eb47bf13b256ac656f3f3047fe3c3d0ce929ecc9279cccf677563d3668a3836d1c642ba97548482cfa5819091768f691b8afd8c14626b7af252b7ac215f9ec9468bcd0049f278ca06bcad54a3e2abc167e06679cd04b1a93a8571540d87ad8277523b18812c4542fbfb90840c7ac482455be87b84f1284aa3b90fda15b50d50c1f71dda606ec6711568030456eb29515e472cc16c92581ab55c85dd8be46c78a99e9591101ecada8be2f7c52ff0443db9dca8401c125a63934a17de0d991e7f20123e414f677f5a4407f19851eaf3b1f8a80de85ad3fc8ecdc215e3224b88adc463671c60af0bb4736d167d37b967afa23d72ccfe1f388667084d5372f0aaa3aab4c4ec7d01715428dceb2842d8d6b95ef50efe3f15472dcd8ca8e144e751242afaa242cb3b81b7b3b76ad22e39860307ec2e6b9581c66956f9e4828361dc373bfd07fdd1a7efb7d571727084689155094db5046219c9e45162634cc64715ca22c5f50074bfc610fe870a7d740bba7972104f914a15ccf990f7c5e0795d6dc5f8ee2e5ff2caa4be253c84771fe1b473190f4ce9216c3968b135fd4601da6ccd9b6126ce178f4d780484b4acef12ecce5e2be9d45318c7571ccafad9352e9278228fe692ff5edad624e8a8403caa0260cf8415fa898453c7746ed5b9447fc07d2415f3e2b3dfcd67d5e3f77516bb7e628810547ab757472aec4e28c368cb1a2d868ef2e1596cfffa882a300fc23214967b1d0849f5f972ee16f440f9f63dfe9e46bf1f8455e6017dca56c50de2a0454a74bdb591e6727cf5812007025f0bffdbaa6f728f2cdda2ead9966792aee2bdd65002460a2306192e004b2f93315c28c7f87d82cad6a89fdbcfd04edcb7af0891a82faefa6eeea74b06ff587606e9848fcbce15d7bdf414b6f8fc02c966e408979789e27a06fd2e28fb8dc2ccefcc48cb8762a1fe9fed902ffacec4672218ad83bf32a680cf5919563acd35a7b685f4fbc35a97cb2347d66b6f5b5fb102579f5a2afffa2a14f065d8c99d40dd253814d8b0788d73f5b078ebe4c58c7d2ab95ce0c1cc06e3edcf0e2d52b5fe25492854ea5ad4b3a439711c3869306102f772d2868db7cccea6a6c16220837201741239ed317c595193d0b1a77716f1360b1c211da82319761b4b6e3782d107a80bdb8028ed6594223c98f07c2cb42dde5fe94b95d0f113bbe5824f91fb23b1d8335a7bdc0d8d74f2d737407488a5871f859c76432bf083eb79be530b1ff6a0826b206f05a7b7a2f6095e54c745e73f6db5714e697d89d4867613a3822a6c30a20b7d9e15a1b2cdbb28624b845d981a8bb2bae42137eaa517e5891975f346780f680617e4e84a08dca96f24f55c9c7630c577c2b0a1362e6c52b51221bbd0300a80686a8e0e3859ef4c21c8373c6ea1c62ac01981b8c869139b6d7cc972a1b6f2e8f07865e58d9b224cfb2b61991d53f1b4a5bbd17d20955d76fbf5269e831e30cc330a2d188369547478e76e8293726bee1f69fdd71428ac72bf61de1f39b2469d938ad0b6bba3ca684e716c5d48e9963aaff2b275615cba3998cc06dcd0307c13c9dfe112d0b7578a2d69fdd203d0ff6c47e243b38b19c0825bb3713195fa8a7ae5e4b847394cf305c61f3ccb9ba886e1b45aaf515e216b3bb43c3a354df4aae60f0fdea19bfd218c445bc63e088236907e44923056c268317209720508a50bc2b57c64a8b33d9de43028e8074d59da4d58e466242a7f71c937c429871a56daba27e1a5d207c7d2fa3433ea9f0958a343e79e6c3db192e2ca4fb47;
        #1
        $finish();
    end
endmodule
