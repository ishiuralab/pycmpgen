module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [24:0] src26;
    reg [23:0] src27;
    reg [22:0] src28;
    reg [21:0] src29;
    reg [20:0] src30;
    reg [19:0] src31;
    reg [18:0] src32;
    reg [17:0] src33;
    reg [16:0] src34;
    reg [15:0] src35;
    reg [14:0] src36;
    reg [13:0] src37;
    reg [12:0] src38;
    reg [11:0] src39;
    reg [10:0] src40;
    reg [9:0] src41;
    reg [8:0] src42;
    reg [7:0] src43;
    reg [6:0] src44;
    reg [5:0] src45;
    reg [4:0] src46;
    reg [3:0] src47;
    reg [2:0] src48;
    reg [1:0] src49;
    reg [0:0] src50;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [51:0] srcsum;
    wire [51:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3])<<47) + ((src48[0] + src48[1] + src48[2])<<48) + ((src49[0] + src49[1])<<49) + ((src50[0])<<50);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1762fe89fcde51b7f49190818dc7ddaccfb879f6a7390052f3788b9f278170433adc6a5c2bad600c9a9929b8e2b1ab2ca233ac537c0b3d95ca89ac731b47d968f85bd90768f35df7091357ca953e929f996cb4251;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6adcba6dcfbcfee6c4ac2a1637802d443f14428dbccd1805d768977ef34401bc001cd64082714b5aabc0f1b1e0bdc6de111149ccac41541bed10387cd22f8b80882dc4f05a1a60f5f240814d7df4cc477b42e45cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa0c4a99bf9e3f37b5f8c8845d5c42e8c921e5113b755dc4172d223b53d113b53f0a73da6b6311adc0bf50d0d79bde913529fa708c0b0534aaeb5aa329f5757db884418249bd9d24681894e050f2613906984a07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcac244072868b4cf14e66883ff0f2f8ac3bef0f598d76940e08d33ca737a641c3d4e16ed8f66860b7ca1089354c6edaf1f35edfc68c9bdd7a3d39b5bf4fc3675f3bb55f0a3a86c0c23d9b27c563e7bc3ccf3dea47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed0d8a1f804bd7207bbefa4ebafc61003710785e1126b76ffc7b24f2bfecb991cc5229ed0f0726b2d98cbad16620f4e0d750ba79660d685d9853c1c93d8f04700ca67e3f95e033402a183b072ed46b1b5b0e758fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90d8448b50308c33a42e847912ae015343071084352b73f0cb7da344b62893aa3460f62d36a5024eb6206552a17f129321fdf2ed3d79d2b3b7d71319b698903d2b12d59858a6b0fbb15b1fb456ddd5c472cf5ff86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff0e37aac4fbcc86f662f04b0632b56b2299d270dd6ed611374b30d6d6e2415d16c59805ebe9b546c76987b377936e2727dd3ea8adb7366e88cd2c86f18ee91f8dcd5e3277447716d1213f43e6b159375bb6d1512;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8aa5fab44e16d5e4b6ab93ed6bb94350b297ee54957e1681779e1abe2a5758f857e3a550e754150d959bc4f5d51db933ae9e6eb4e5771a5dba4b1e56290c35b9137ffe37cd65e09d14d3541e287d0659743eab40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha66578a40d15e86d3afbd7a00a8bdef0a1ede37033e0405159dcb7ddb246f66dccd8ccdd52c3529e2bb65c0665019929d4ae3b8ee47d3de85c7df0c3a8683d52d488c29da7701d82d3596047355a42fdb1e7dc009;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38b84dac4a7f98d5b51ea8e1155e148a1ee334e844564e8dcd1be1c4db6cf7df86c6c024789d90c3cdd9e95e09582f98c935cc96e37330a8f56dd1c5ab783cf4292e1ec7665bbc292d351a6b837f0493368e011b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f36aa78eefdf7c80a7a19f7be13358cfa426f67f639c759b34543cd567d2bd78ce1377a8e41aab2f0c9a5d93e8e1feef2d1acb470de4f650330ac5c034a88c8b99b4b2b61cf8355b22e3cc6a07e7389a7c96281;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacbe26c68b54f9e8dd958005f1da1b328b0089044343cc5ac4f437123b59405f9c10db7323ef5c98d45358ab93b552758c3d4da25d6b435f73708197793f35a6fcaf4a1485b6f58c18cbcaa26d09fbc34ae7fa99e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a046282a4d892e739e7c8938584bf0a77fb97659445995839b215672056f9ab796d4a404ded80408e513fb116336fdb0a5fe97da728540556f7f40962b61448ef2148be641c556e4f14c3519b78f48dcf6effd06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c9b96f13fe0c617e3497511ea9b386fff747902e950fda1f2fd7f2cd1c25c0bbc3d9470c7e8c0b0abd7e0f88bd8df5146af8b612b18ab99d41840524cfcab9361e9d2415634d62da290895f92dc8dd9b8230092c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h435584ed1d2d82ba895952f9b05364ec9038922819a136ab9ead1a0a3a128fadd8c8ff963bb241044f17134671e8ad4919a5d9364832d00e382547c5f81d52763e6be839de9334f5a8e8c1b3299571e86ad261b50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9fb12bd5a9e96614e429a4379eafadbfd3a118b3a2f52f5979cd815259fce24b6d412d3cd6c24801264afd4da81df80c82db18b25f9bd7d48bfc9d54cc6de47e5f968a74a29980bbf13e76d05072f44b86a10a88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ba6f78154b19fc4430523ea71ed3118c6e3f92a80cdc1273a45ca5d948b4162f76a09cdd8080e36e1f5148cd106ade22d7f197b053a72d81293580a5b85de74f8dac607bcc463f18f1327f32c9dbeef233f1b63b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb31cf713dd328f8227219d0885ab378645cecb6f9c64034b5bdc452dadaaa31545d4405435889ec526d7d731248050e7a7ea6bcb2af7597a42510913dae7b4ef268328a6d887011786ca109fcba284f6b1ee46dae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9296c711ca88527203bbf535a961d0bc7d6a6ff9b1887e2c00baf4a8cfb86a183536fe42972af5b59f88af486897b483b1608e03002ce2460b73ac0d8f40c2ca4bf634a0c90449aec3c12699b10b00010901438f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb44b501076d6fd2759c43b3a790023c9a86cbab6f4e33144279af8b55cdf76973d792c19b244a23fe60ed742e4e44d49167c635820becb7f1a2b8df915700b27b2aedbd13d14432c46d46c36c878bb5b72f13c317;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41bd9101dae8ec2aef3aeaa05773812459dcfd940a18217a4005a81352db7e909dcf5a198e8e2e761496c7268b5fe7760560cb437616e08a107cb855a19b8b4d8ddbc1e89ebb9686caf173b6b9f61ef9ef2734456;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e3294d7b6ffd1ec57a0fe649698b32ab8cbd4ebee2ecb879612051738de3561cb4354fc449c2944e9fbda12b0dc51ecd812ac7cad09a57c3b54adb315f39df2089f9b4931e5e39887e71baa72324d87f894d08fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcde50f57f5eabba7bb6e480f051e328eec806a277517602b2063292aea0fd02b6bc9e8404c5498654cf1ea5ace350e596fb954c5ebb00a2143ac13341e62dd75fd3685feabb766457b81ddec685f02698fe09d0c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3496dd5c463f536dd625fdf8778bca0fdde75aafb466d226a029e141a6c38cbe31d2517ec43757b65f7e4cddc9a41f803936c9ef45939304a57928adb5954532d0805c574d0db003d06cce3854e4263c992921ee8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he253e338f5446b0a0e24df28a7374d4084aa9a105d5f56e6b981faf5d9093e70a4d1ef32e201436a85647a8312c9508792373cbb12a5af02da2e242ed9e35d21522c4dcfa1dbc0bc036fc991806abbbd70c8a9efb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f0a80704fe2f38e80eecd11913f677441d4e1825410083b2bcd299fd3532aaa2324ff0c83dea0c3626c57f489f6326adb0af2036e960d5a9ef121120a09858b981c05462c6caccc695f9f7715d31d4850f72b47c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h806a5aaf8b9e65ddbf296ad0ddb31dbf1e0d1aafe777c455591cef0881f421303bf55297e33f9b817e5f768d348ece989d3ae6207bd777e40600e6a908f373764ff9c8d9d130aa499e45b90860276e1eb3fd3b35e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8092c6e84e741df8ac9da2579adacd573c9f5ceb3635385b38aaea841ffab985a94fe0d67cec92335662505c4c748df89b22389ae9c2f93681b9e18848798f1bf347da6eee86b6bcdb73ccdae525553f6155a97e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67fa9973021a0f4345196d1fb757931d35da1d6a6677bf667823940c3147d2ffbaf3a57e8f6ba895fa20593457bea1bfdeb2c78c4acc4cca8734f9ec3f563fda3b4d66200a9ba6a5b8fbb4de5b3be3dc6bb622544;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2055209148cec3cceeb9e7ca08f2a31c25278fdedce0ffb30ce7ad8622e582020f709c2bc55ad2dace03a860b475ead1bb361b3807356b5ac92cdd710ca4557f3c97e8647360e4e256897e71f078a0193396b42e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9024856ba2ea22c668a7b18e058be4a1e7d0e1bd6ecf81b9502bb74cd4dd4ba20352297aa59a4a6a3d7c138bc73047136560db60a8a05d13ccb09d0b51762850c84690711ddbd2b0381259a98c518cecce4e6dd4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafbec8761fe4c9fc14ec2a227022af8c6ed3110f0521f5a1f52f726e555038a323806878f54e23ee7c84d053890b0618ade825cf393e603049976dabca2741876e06a38e910358b01a0c24de0ff6c60ae1894cea9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9a832d971245be7f22c8e10aa4c3737e3bc51663af8171761f267ce64d30ce399154eb114f130be179739cc838af7a5da5b2442cf7928ab7d6cd413b144145534796e237dbf937c89fa9097ac62242d4e3039206;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5bdf1fb013005b257f362666b796ec1c0c68f277377bd7cf72cb8eb9f061471f477346b6d5f2270fe0db7e85f3159e108311eadcdd741480e8d66bc7015942ff1dee890a33cc71109278dc15f6392683440b742d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h455e679792699278739bc76c7f27d3571948459b79689e76f6e78edabab7a013af6a78185830d26dbce083df52fb1c9435938a0164a64c8ecac2929cd15e8c96f5c8ad0994160b107aa6019f5fbc994c8b10f0418;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hece60102734b2e0da0e3bb52c77a2e7024a95f3e4dcf73c202c6bc711410880c46cedec23498294f6556a075766f1fbde60fd24e6a7ae0fe1b1a45cb5836ca7bd1a7125c578c5add8580cd55c14578b5370a2fcac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfa2df95157f52051eeba464e5927b187f37509be1a3f7f75a15d1804a96c1ff53cdd8e5b8d4f4d950ed8e77d917e1c4e75e55c9d7fdab890aa1c017a378fa68ab62e3662cd301b00f367a54a4e75c745472df7b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h209fcabf6662c31215f79a7d7a21538850bfa71cf0a08af589f12688bc1338f5c81abcd76150002ccba524e1ee68ee22e172cca2c151050dc5976b05895b44054bf84d44f4f84d6c4d4d68a6855eb70e656eac023;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf56645de863e1eaedef416cbf2e9b2f8e227542ca120cdc5e3105c878a88b9c12a350aafdc534bb072937dbf7c2bff61faee3221611aadc45b8dbb80ea24c67914161ab5e760760f31edaae97b9ce220ea8391477;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haea7d4e5bf29eb46f50809b17ed6bccd0d16e15bd074261d71226dcd77e8bec551752ea73b51c138a149d9dc7d74ef224ba29a2f2715fbaa961b05ed46c92d07601f08ff21f2692ff520b18142b4823f54ca03b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5902a76d1520460c48d4a72a3334eaedc7a63b60f9ead131be11b958a2d80a377615dbc349a55c3625f9cd4d9deb44073b237e240c9f0ade64cd4a4c94253cc72fdb28a8b86c130396c7fe7f2eeee258d45fc46cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h132845aff2073b629b5e4bb09ae527460fb7fcbf6f69ae239bdc3f5a12624b4d8a7c32e9413f671df90c8fa1c8d6fc02e8abb6641b6f7fa588f70d7d8050beaad4935ab198019c511386b96decb5076abe3f606d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf420a3263f7543ec006a4a3305bfe4ccac661c4fa30f1c91eeb22968089d3332d352e1dabc633594fdabba9a47e47d3a0046e0d0d3e113498d1d16a0f569de8bc6cd73fda6293928b78e5f2ad695968b78ffef32d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5400db57deca852e001f2a3ae07e244f881040638fa40adf197fff8b1245fe5332a7c652c95793cf8c1c60306af077eae2eaa77e6daa4755482e46959035735e19db620253b8619462e50021f7a533159ecfa20fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h333665446f4efb82e17c3d7e01a87ab312640d295be7941b19af5c91151086b282ecf40aa1e4afa2e609b80b8e3a898c59a8f76075ff159da62280be0b1e694e5d9917a16dbd8b39f1e0cb4ad1f7b09a79b274588;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e673a5fa422cfa125bb3d85b047937e1f7445552392a63d7c5de8d0dfa6121c7d68514c9e1c5c3a9a4ea78922a3b226cb5d11c8d35957faf9f9a4039ad66b40cf0ea5b984364d066a12d8aa2c17043bf7045a4c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb618594a4f3c06900eda6652ca5b5948ef544a46a08d2b76458da344ee0721d15e04c2c59841c9ed33df997d0cc6af951c88f9d71760a21c9b4c55eb9e6f441db5ba736f335fd85696567713c756aed51c73d73c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cd7279a57f28de9c9c5be0b42016a86b0708bbe216c774f06b4c9adfa3f8d4d3eb9cf6ee48cebcc2a28fae5df72c85310e6d79e1f0b7be3aa1a739996978308e78a60502f6a3d66b3febf7eec5344d02527c1c38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h734b602db716908b46c0c2c00434bf4b60acca1a295cb99321271881e69fde6b7529907cd8ca86a0c6a6a3b629a88b426f5a412caf4c7e12a2e89f4121eee9cc7dc879e1078a4565e160a214a524ab8b3d7e24c8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf3ce535a162e2c979521f170697c9aca4500a5a82725284fda46481c227ff057fda134817bce6d8e1cca904accbcc8346042644fba670cf21808d15ce7e3efb0548c92028e7b8c2a2400637b5acf89597a0d513f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd68925ed0ce2f1bf4b0837913757f3655f4dacdb38b5d54426cc3d9e35d6b153fe4eb076a14ac1a738d378203d7f3ca84815d485cc2c4df064d52ad978bd09eb81c004e62e35d773c7326168a52517de1dbae4777;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h927e9939ea8b37a375386629aa201eb34892228b42b3e79598be226d55ca79eee34817031854db2beb165fb5c2b59777ab78988003c1cc55a38a9223346daec2cb4a2330c6988591eb540037b85a1055207fe372d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9d3fa835f744bd276215e5de0c24321bdb9a631dcfb69065412c4d2679199241530d93e7e284a377aaaf1107229678b8fa0a9ca1229eefb9a4a07b09a6000b62e80c825fa20c7b1d0625a929e2b8bf44163c493f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4751c369794015f3f19c7cfbb62aa684682c4a824beb93813eef9a27299d7cb902d9af71b075c34e50fe67cfede42fac16ba558ff47e0cbf2ba4fc851aefbcdcf9cd16abb439ddc6d76f978c11b8c76a23a369a68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51e3dbfc9d5db5db1e18783796bcc143f834409331e9d6215e1a8639413fd0b294cc57239d2a11311fab0697fd27bf8f251b7098c913e60c74b4e66c56d15d9824cbcdb8bb2e5c9cddd864911ef26dd7a6d450b76;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f295f2ed577d0de33a979f6d6b447d86545686195d0c861b7b426bc0d8f3f6d2acf533298e7e41ddb3c4a603684fe7ee98d0a714bf2a2893f25c729fe584205e0149ebe80d404cb56ee801ad7caa7fc1375244d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bfc0a6f35c7ff6073d2e06444571aa3bfd1c5f7a8e5d7ca7c456ed7a5c77e6bd6196cc97de9cb3b5d4a48750c1acbd26797f832eed973380b9f2ba6d5ce0e08afbd17bdc3cb3ea9f5ee7c7544b2beff91a49ce89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a016d68cdb53edbd8cd04d84be1fd485d2e1d4d157a57e694f5cf1a71163fc2f9bf000fd161d121b14e7a605afc427b18e523e9887950c906111b242569a3d5c936204df2aa146f8aef5877697a35bf43bfdf405;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b6c2aa3cdd3ec510fe360e5017f6802451baf4c3f07bef059ac43c2c1b7c0a856b3d7b2ce1163606c97d23139625de3435287904c2831aa4d71624dde813924b540f73dc64e6b8ba4e3a027e121eaa5e5f923c7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h610441688893f0580df7c15e75ebe4258a70897a8c73c5729896fc02e33b6bd2ac103ca4350306d1ae0a2877ee5327daed7b8b8f802788c633b02719c86ba0567dfee62443fa7973150941795cefd2c920d91ed27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e303d70861bfc8cf310532a61611cfa26ca04a245b838635591f4db29c6c0f3cf517cbd901dcb09cc630c6bf6e7ec8bcd6fde12cb5f1595ed55ff94c9271b5551e19c88b544596489c119b004dd0e31d337d22f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8cadb02acd39592ab694fe30cea208f3bc0e9a5ca2fa039df1942cdd6e2c454910a687e4d49438018a61def5c34de4a77496e182dca65ff1047d9975ca07a775d4e269dbb3c47c41292cea205565e76c6cf7a846;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he25a0076b91af83f07de5167cc0c2ae4ee26f4cd6669581988856d15daf0cf8a077dee558afc9cb190e7e540cf7ea1bb94dbed07c9043c7203bc2cae6b7d44e43323412ff4b545da67bfbc511da73d5f4dfd19fab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce45c5c652a5d20b8bfb51bd7fa913da12c483123fe85798184ec2afc768f6aff5e92d83302caf51b1ef0596d072db20305bd8a5443b4b289d245761777a5b1da63aef95753618927a7c170f95d9778654e7b6540;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16f3027c27883781dded7d41f6f6f06aee1d94f5ccaeb649ae42294737c1f7b34c9a8b0928f540bcaf6f6615d68f6dcc9eaeb5e2a3064e2238c4c0bceaf70262c4abe4a775dabf570cccd695743a354f487ec041e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3601799ccf13aa03d950692a7e1083686760d95dc26ee084f2d7fdf3bb470308a4b8c443e8e273688e4da6819e3c339b00136bb736a54a58d15880099bd47abbad898f545244caded196185c2cff0249470cae339;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32cfd449e1e8534d6520c0508672d9d4a818bef76f7b6196f8b251098240a771920ca2b6a3ed87c0e52978b38f9da3cb9bf79a00ded5bb06f915d3acd8a7d368eefea0af5f624d42399a705606126ebf6ed48bc76;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1b473e682b3c220a3d81031d028acaac854886b1e6ff8d01be3228b5badb5a61f864ef8a002be5a9f8fa7aa71a66881b85851e75dd4591b4c43797b8415669b77efb7884f94e6b4402e9ef7c6e3f8431ce1ab2f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd157c798eb5bc96be6bb47956ddd1ebed8dfac29c2b396d5631c182c5f52d3abc220da44d4827eb7c29d883c0e3c22c60bc221149df4bccbfeba832849709cbf125ad1f627d400b14bba373cfb2db7a2cdd7f6a2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32d995b18ae7fc1c552be3e9a0bdc230f26ab4554ef53b316f71c48ae06a0a9eccc766f8d81f38c9255b1f260610bb73aa3d0386da980fd6db998b2632f10642f01e8373e725b54bf88a9686be10a0d05c8e46c9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he41b119481e6c62068d830de66c9303dca82b3d6a3094f89d8d81778256f4118c84fc8d290df8f1de9095e7ba4f5156eb262171a742e5fb06171aeaa754c81061510a39e32aa6bdee8ac263084025b9d7d47f24de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b31f8c6b459cd42bbd28c9bdeb562c5a94d7027e54177bc43497b41f47dc8601a5a9773935f1e88b8f69b011236fdb57bbbc6ab4765199281537a190c107703705ab1cbc02f797aa49cca3eed9ec210a5ba5691;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b435454883190b8df69be371477257809de845df652a73a24069090cb199cb285054504ceb3e0b19498b44fce6a9fedd85b4331eb10e4aa2e5c04d209fa9d68d433a8079399eec9989bb8895310d6e1ea08a8053;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61f3f091b9966575623ff5dc802f9566a612cc363880eca005478b54d3821b98107fcede8843085537b05f2e95c42f2a6d829530f4add88254ee93551a78f996117930aac9cefe3db8dad04b22371877e54caf82b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h200c8dd18a81790493449337174db2c3a59670a361659a88f3afeae2cb286b1573e5e25e343f6124f1cda5c856db2f5f5ee9cce65f7332d7d4b77dac1175ec5cb304acb1240c384f817044e69545d2eff5a7eb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7ec5f5a2b9df9d9afd2e4df57fe6b959a4bc26ee89ab55d6f0ebd89d8e6fc0b080899c5626cef752a21503b6b2d830b573c2e0a54f9b7f22319eeda5ec9faf9b086e53034381b3208ce3a20d0722f641dc969847;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba7e80a8cb4601cd6d31d38ed03d7ec2b0b8ce675e810f877ef0c35f3004bc680fd269275aef97df98aed4e754e9d0d6b851b3fe6238a9435c8273d2dc2c0b233f949a77dc18dbe86993a1a4bab208a9a3379ea2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a4d4a8649e0d1850ef5f270e88304a9d6e843c99cb6cb07283f8d6a341e760991a06496461dc0ec850e90e5672c1c60267eb5093f17e0cdcaad1c8aaaf9813862d1717764f013902c40beab85a526514facd554;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde4e0c6a3a577bd898106ec09c9a05c01402103f7c68e38fa8fb3ada03a98e99e67f412d82d336ad6d7b06b8f7306035154c7c1212f192d1f461d11a04a785b31866f72b93c90ccb1431563763c9f7680253a213f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ecca9a585577e25f5652ab8166453d32790d3eec96b8e81358247fa507c1c80931e8e409be1f27f009f72163479076f3c34ff26d543d534f23ad539381eef31edf1fa0faafb192dbceee46ebaf8ee92694c832b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b6095f8c69f2ece42dc0bbbc6bbeeb3e346449a62a7b3c07384b052e613070fdee1b6f8709f08803e6a70ecef93afd482d03366226d47a5839bf03f95b483a2c8e4bb4d8a6b47b8308b68ca40acbeb01b1156c1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he49eb800306e790e4e40861b9ab275ec022867128d04148a5e7d12de92190acb3e8d2cfcc79603df505d5b634a2aaa929829d774ee55f9570e8e61eb87f681684662ff4a40eb3729bbd292998f9b9d2896e3fdb79;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed8fa4257c59791c173b2b0ae8bc475c8aeb11234da13f575d80706d5e93a7a32cf84c2abf37826925920bd5b844ab975810553f470396560db52990d5f6eacc0c7e7d126edd40b2acd1c39c7d774b68bc59ea378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5f107938f0ff69e2461fc6ba77a648ae395375efee00849968e8b29760629eacb3b6479c1954b49fddfc877c6bb64b3e07967e648b4bcff80495e261a554a136305daab28542394c1e73271affc9f8cd39da7e2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2c1d2b643f6c4f114a8bce72103ae68a4df21d2a72d904daccb3be99d1254bb034b706e5e4221f57876b08f0197de1c7920b735cbca560e3e5a4149448bd6fab3c21c6fc0a83867f96fdb22c57192170f3075ec9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdec376753a724f6112ee25e3cc39c5b3423c4ecfccd2b1a5e9638f8ca9cd18b697984496bca7e615a60a1d9a21ca1d649943c5a24b44a67d7f37b08cb4a6c0633e0f3b7ef9d8ab10eb9d8dc02f2383c3ed657686c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9098e84869b3969dfe3a5a7693b2951bd4741eef2ccf5a579b0bc074c1754beb24c6369fbe1482b44b2ab67a8014a3a8d3b04295676ad3e58080697c243af78416bfa112bb839d3c0cd482d2d2dfc5f4b51e7c31;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57e234ffbf5cb0b764fa0a38ae5b37c2b8b59d352ec7b8c4c2f3667cf5e0db5ca8d753c7e0a86b9c7d0c0dfefe1a2b50b232f90896ab732878827750d9d9f40767155a3193adbc4dff3ebf2611100b414f15d5cef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd98bb57d6e1a109bc327ea3751879a74bdbd3aa6a0731d5ff119cf39c5acc8c34c11b2597e7259b43adf60def376c3586c64e217af13d42309e3e1cc0403f2f9d7340f819274d7b98e2387231a2c7578d5b157fc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b89f91e2013c91284b26129ba1c8b939290ef25d42f407a3cf700930a760aaba7f6c7ef97a8835d4278c0c8506b148dc7483c8629d112a42ba6b02129d380b02d9b42aa386ca63bd88724a7eded5460f56faf606;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0c6ef96bfad28752efe658add54eabb73beda7dd81058c2ee53cf7cccf08beb51fc9bcb4d8dc6529e8ce5cc2d9f0661795e035ef01e81f60c291928ab0428803e5da7c8968e4d19826d5fb00978549e97c8eb4b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haca2bdf1c78f159b32f5473ccdc3efdbea8e82f38e2691333ca51a1df5224c9d707d7c621c779161a302a3866d26ecf34ccd0d337d37e79a6e9c2d434de1ce693c45e0738a516002e53e035660cfce0cb221d8a4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd3c7857d46f75312c9e1df738ddd2d2afce8693a2fbb3a4b373b109640fad4cc8d3ab93350ffc6339d8e48818a55aff2fb303a1490c335f6561fedbc23ea91c9dff67d898dd7e2dc6ef26ea948c470519b5f1b4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb27cf0d57ce768636e8486c3e0d15bf5d7c7c4cd77fb50b4f8b4f68b0c6f8c59cc0bbf0fef0b7e639ae530f9928be462fa02acea7c123cab35cc7a4287876f6e9dcb65e65da59ef92b7f844113b8905b0c875cf0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4539015fcab934b8aefc4b605352d8a858c82e265c90d85292b03edb7fa740c321c4425d1c8ca2774d3934302a1b8a1f05187c18eb37de2b0a5b2b66e7567dc1163585602842699ecb42baf3e8f6414910d2cbca2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd8df9bf5824abb3f5d2e3b51d14ca54be6d7ff1ba9ecd84152330c801dd6510f3b9c9d2eb26e0616befd1481ea297bd549d43d53ac3ad94b4b297280515f87971e98bbeaa87a2354b73a93551aab9c451741e33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb5379b361b6e5b5c0556768194b07b165d6286c2bb511562070402d942ff8172f4988a5ab5860174e925ee34cbeb0e49e777f2fd1e97671d623a13a5b12723454114144d230b9e42a0caf9dbbf832f0bf21223f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h655ba6a16c032dd7e25fb1e6c0d4dea18a2e016add5c5f012d8881f9da5377c644b522497884bd0881c9b5764c342f38151ed5977620431013f06eb53d12935c5fcc886ac984486edd02a7e6a6cacfc0e2b9dafbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha073e9b9cc7adc4769466274b9f993df3f21fc65727df1097b666cb1a93e45559ae708d09abd370a4c206672aea4999962cbf4b06dfd5af0eee1bf25f583f6968f12806855e608d4329beb2507d48d3896d281ccc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe2523925e2f12315f512d3cac3f7bf7a6d50feaabe50e989cee4c27e4f6a73f0d3d7df3c93ef1edd010640da795ae239178b4e588c3af9ce86548762defc80a29a852146e7314fd783caca2384faa533cb552b2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45cbc13a792d66d70eedb831b3c142def2957c672e4d3bb8ef6e3c7f5c29a10ee5661f6847cefc2c6014aea81966516de9edbe9ef99b16b394c4549e26a1d35ae77cfc35d3a0e47e77d26559e0d8fc9f645194c13;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22a97530e7656c7eaa0faab58fa181edc27bdcb562aa2396764e609eed6d1ae526788703652cfbaf0c149093572488da07f7b661c3d4ed7fd7f4058cd06c36e4e950f5fc18e1ce5b14e02202e514186537c88ac8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22e27214b0f7384eb8d7fca68e37f343974e62309debcfd77f82806c09455270430b0548e94b14995b9e0d2ced7329bfabcb6c4f451840d4b8258126245a9c8e9c4868513e2de5017143d54b572f80dc292454d0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h580a39df0c6013a4d4f4fd4f1388902baee98b5536c0ee10b0a81881187038b14ea3f9787c289358adec4adadaa5dbe19ac4e339579d9042ce9027e224298eff4f04c7ec3b9977af0414c1cfa57a45b3ed1ef76c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h805b1be1133aacb33d158b5d81d3d727f6926e9cedad0c2bb4d4cc0b0ec01393d189365d2ea00c03ea86f0e0e5665209c57bb9a3530279070340787b41165c5e196d53412ba313877f2051ef107f857e84877903b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h266702e000363822acee26f3dfcbb015d9fe1ab5951ee5878b7dd05524cefedad2a4065b7ff18e9d7ea51b7ffc57c8bc286b67bcfe78075b67ab185e8d16c406f0d90f4f522c239e6febffa8fc4e9ad8156d64dfe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c02d8534fc94d44ba9afe9d73c770d01f6e749e768bb88f58e43021bcc8ec8263c0e1fdd4129767490f376334c46e56fc5d8a33566549fcce7009513c623911a8c1dee3006cf1e3229531c81f9df3a34f388f564;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h575890afc45d66955779e30cc16ebf48bc688c59024e202f71a45c3f25bf2e46d8ed86e4d76f933ffab0276d0174671d573f848f67d0b2f242c35659185c6876f5127ca0754649a3e562997bd4e91dc3ed953f389;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb135e6688d839776ff04f89e949dddc94b029e1214cbe6a1d96d15becc9482e4614ab656366bb83d1cb3a6f4ff9e07132de03f0e2065a8a8b020437ca262b5638c686202c32ccba1dd55c4f914feab6a1255b34c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49884a62b92d78e3c91f27eb3da4a6cf865399b547a98b20864344b9d2d211befa145dffe4d5424c2843c44ae330181be59611a8e0642e76b4a58fa248c03c107735879d8a44dae84743f6720b2ff1a37fc31441b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5c7c01c66077ad679615d728568c63210c9f67e7ecf36022a9cbf14bdff000dd57688b867e3e088b928c71a67d2068b528136d01c38bdcd1761267f33204736672162679d85a8015e2b2fe1efff65efeaf810eb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d96e6682836be548032965f0874dc6fa96de23bef181f2be70a39f19ca2117ecb2f296f137d8c240509026329de35cec66e796d990c38c6a875310cc6f3f372169ce34891fe592827d4f9b4cb10a5763f0bee8ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha43ab6990fcca88c094c14a48754c16cf558cb014c5259d85cf1bdeea03673ada026ce45c13d7b7da604919b4e30a8fc29789fb0f597270f2f1d95769653429a3e2590fa231d5adb7ad3de4dcde39395e6414c834;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cf8079f490d603dba78f00b22dc9a1221c4816d501926e8c6b2255bf8002a927cba6bd07d08395e7ad08c626bc206cf1c80ed270e47a2e919b38581643fc94b05693e6580b10277b1a30f0b39593bbf9d3b8d939;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he06c4566893e26dd20a004394162adf088fa7d83f70aabcc7ce1c92bd2d2c41ad38d7d1637c8897f5c33e76f186c4b292b0776370d588f5bb6a7062858ad391a3856597c4118a36c6a3b7d1dabb0819efb74cafcf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a8bd194e853fb10b45bb86fa85a5f39892f78e8c8ad6deaacae1bd056f8e2b0e65ace27ecd52880a7d8f55e6283ba56805dc29a4cc8f9dc8cd4f6768d304ce47d40a79eaab89976be114c4230b57a6e92f05ada5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5732c8edebb9a235250bfe3231106354fc8fd3e0f4389487ad1702d79c09d8220c124ee2a7e9679dc303c2b0c0dadee69c4a994f44a4541d3c64f781fc4bad66bc2ef5ccf779e9c32196dc3c3dbeac191dedd18ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb56140c9cdc73944758c6ddc4002c7b2e5b3db7de9b08c5573136500b41f1882d470a0b12a9b6fd41b835b65eb9763f82bef87eaab235c831daef420938337c43286b9d97b5d233d248184bf5414492c70bf7d1f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd6af9cc54f2d05e76b129b2c58a6a163510acac6c8a990784a749be12b584c3c30330c0b0b072870b0076347064c9b2de201ca43e7b17fb932a80a1a7e40cdcfbff872fa45f78ddb14f287bf5e516f1cca3bd082;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f2c911b141ffd6ebe66ca6e3a95d971bb3fe39ed8525a9bb0bdb9aaf2af399ff74c56104b313ada2321df66f6ca426f08919beb2dceda5ee94fb537cb4e54845121f0b63954a15fe7bad13f4f84d21cda36266e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a2f5a54dc70beadf3a187fe862187ab528ed948f6f9084956219aa190c08ec448b29bafff0ac2f5bfac23b2f97cd8a78ab6722ae5be2ef972ebadadf199292b02988d581527db3fcbff80bc99e447e6350f9899;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60c5f4a6d15e430c48ee40148938bd3a68d7e94f661094f6a4038c926a612d41a3904fa9c49d149b7355d4db1d68bdb40ce79a35c50522f5903d059e1b24b58c3ab95d986c35faeea0aff5667ade4caa06860625e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fcfc00b6b70288bf1be68a2f2d81d37f6cf98a771f0846a1534f7cfb21db257c4c549df3eed137be050a07adb99f9fec2da51ec7cc40a6e23ca43d914754f3686b907d26d5e5cf062a8454c88abd4b8a34d8b1ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87913fed78556074ea985e18530c56852710147279b0ebdbc66ce51bf3c3579b4b303fac6fcab10b0e19f730a70a78ba6ae7e6400692967d3d09301d8de85de4a4bc4d1d93918b3093b518c2b62f203b529bed7ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h657d174b279ef2ed7a93e086a1fa9173834bde6540767ceee3b39d9f5f6598544d7f58f47cb1e418d64a1712325ad5ce77ae32af78acdd86334e8aec2ac4ccc75f9bfab8fe577563371ec6fbf4c86511a938b441f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5595c301bc6763dcd674c01e41016fbc3db55d9c6c332024266096a97c41b639eaa4ef72c2e167a21a4c6968071c87a2d4025513beb6af3acc6c1d96bcddd1d586fdd64c24ed7f24dc451c7fc1b0140d340affc25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd25dc4bd6ab8f5d2594767e23ca1781d86795c18bc2d5fcebff9883ad06103f51567585e6cee8260563f4a452256bcc15ca3c5ef9d5b603def5a26474fe83b5b915553a247b08d8e5a32d3001058775a649f9ea46;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h142576cc24fbb45459e0507f2f121fb68fb9dde6f11b62fa0f2fde21f4f44cd9ebfbfc351f78776c67d866f6cee76f38f6e66f900ad42847ca21d80c4dac7ba6a0f745779b4c39ff6774825b1989be91f2534ac69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3178b9ee77402b987c4a657d03c573417554ba2e665ba617004521129f19a087048d06c250ee1a77a0b2b526b5115af7e4564fc832299d10b50a82c288f1b191661374be6ce9c246aef80383647380a69e0eb13e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c87c152338d60f8ab4ff99f65facffca38b4bc49a5b2a0bbc0eb4246e04fdb7f8e3619f93b9563472f682291a4d831138cc5d147ea2ff81e66c388d83a9b601ff05d4ccb99592f63760a688533f0543f91275653;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34abe70c6c1979267f1fd42c380518d51b27cfa3e3b66d809af9a99f31e9299e22702b6ed0c6f06e73586d5f66112795691ba9e9004e1709acf06c749fe484912d9f316fb36e9d5e2dedff826217581a6614a6040;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51d9c862f4a4980eff5453eb70e9aab5042079399ceae9bbe6ad081100008d50dc236f710e44cae12ad4b5ea2fbc24408eebdef0e12478f345fb444cc15f71fa24a18e75660f8aebdc4ac89538a9bb48ae6ed304c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h662f7735294da25482fab173046b8b40e18150cd056825886ad5c281c8de808f7da368f81f5b3c73dd78a11c0bcaf425f48a5d817acdae42589f3a1e8fa9d77d1f4be9486f7d2331feda45a80adce9d59248e6eb8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff5cc83738c59ff7bf8467cbc031fca5de198e5aad6aecf2df49e05afaee2520140095ff51a0ae6ef0f84bdb95a450c563c790714b50cd2ed7021cc1ea370029196b71864596976508ae3e73cb88471ceb35bce30;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddf81cfc3d6a160f2240f9980ecaf8b934a57c54127a1037f0a0279bafcb332c7e53ad99fee681f7e13d63ad7a9d1c11fad8182462244572869dba4b02e732a3e74211011bae153895e4d0589d51df6ecbb26bf7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbab5d044acc485b4e0c1aab99ac3d414066158bad5fcfef96df27c65da82c3a4f10dc494466d61fab41e416962face4e4bf5b95c3efd0477baf51fce8ddea0a9745744969484eca0d06f66537bd30410936355665;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb44b2a2a0687be0c1d4e20d1487e9d0e23e23c532a3aa96b73db720f06612dabf55802cb8686afbdfaa1612372cddc5d0def6fad9823629e4875601f7efc14e311636a03d4f848cf5d5b81769c3cc67986ad682df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7430ec06262141f6a040686e3238f3e02816300fd32a22a1361e69fefb132b5cd112c56f5e0845d75226d827b30f5b58362d4536909aa178f1fbc95e9966c219c8317234d13b30629b4b9dc76ea933e1efdf0247;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f5d41cc964f175d41a37627b7369b11a23ec14d36d37ff5e2f4ecd46c51701fe225a4945b3c116aa4e86ff573dc3098059d71b1ab268ecb2f93907119888a6291529232eded36becab621f730ed4d33a95137e37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha45796d556a3419d907403d5b709ac42caf5d84f98f02b948b8fe515024ffbe741176673cd3d6d1f52a5fcae6deb2187ed1e857a6f04eab6a78333f431f4651235e4c33c6528af75add7ef8c1cc39cfcd259239e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69d21a7002f23762ffedd64651db4e3ca834ade84810b7c28a1a5984afc4a10e9d3139c843856ca4e16ae97edc042abbe83481bcb9a76e586195a7a8d871875ea244244f97c5abb9fc8ac1a720c46acbb7b445adb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d40be78a147c113392ee9209af67426c50856c2de0576fc117734dfc9d0a2543178cc50d36023628ad93c9cf92a18a5714276d01d3e45552d834a7b1f4e4ef18d7d9eac6244c24739a30795bc4f5cd32353b29e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2dff27574bc332ea5bc814d08b2a24e6bd750e837b58ad8a7ca871197d86301576d79b2881667a05f821825067b7cc4f6b0bfb0ddb45d7eb36e4d3763fd85ed779f46cb94135e8972e2d4e3cd9f3560cb622c93bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40d1b0955c2e30f925920a6fc510378feb4fbebf85d4e88ca1952f3d56a7a2676c95d7f7f5852b7394a5c4c1d2c61112fc4c18821458a1d7530303b4ddfc9dadc88567b5fe02b79960d4159d8337ac369204527a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12ff37cfe41ad25ba0dd8c400d15f5fe3de57acdea591aadd2941046a26f414b96e9b4c084f9e87bdd39081b408cd3f99b10f679a9bdc3ef7468a4e649a4e7b5bc0e12bc5c6af5ee996d907d9ae2ea75b01b7fac0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb198964ef2aaa02d20d7e1f3905209b5fb13509e0d31a11e524004fc07264fb937b5fc79bc2182d9a9832ed3a175a917346802925a5c8318af6c5a1e0cc9df55021b66687d7180174de70876c4f772389a4dedb14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc3ac5d4da96ba81e2fb4e27116a6d570ba6613209037debe058df46cbabd8568dfe6ff03f7e3bb5262c82f5ba136e46930913a1f5cc05a314bc65629fc6fd88f6acac2b6458351fd016b6fcfac0e66356cc10d2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6315aa02c826a41c2b2705d8d2d52100e25985a185dc271a9f09cff6e2f49d7c6eb04dbcc859ef46da46c4194dbda6a85645a6a45cd6396a17ab1c2b166959ef86008de6259b15a39638b38237fb45f1453c124d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1d3eda86691dfa8df41828189a89284637545979b81632083d95d6fa013c4ef0e6f2d17fbc69670abecb2445e2eb34f0713c7390c4c4dced2e25d8f73231fbd89966538e5c376c7e811ef3d7d8f576c51d7b3c03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f4de8e78c8d7e7a84631d93de00db13d538f07f3977c367b84f4cc039cf484ce7ceee67984db72b2486037c3085d0fe92be7041db39104c8ebe0dbe096883237b308ccfa3567dd907082295005d7b0fdea5a0b74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0e0baa1344f3647bb57da3a29bb530762c1ea0ad5235f4076bdcff731cfdbeb47f323019bf763990418df23dc6e87b4f83d03afe4a5c1596762b3ff4350eb434fb6f42b2a87b0b0306f2f070e6c89ae12e17a4f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cc59a1513f1bfeedc4097792ea1238b38042b2d01c360941fb7baef6980306981e42881492c5173e7be78285a9c63daf0e471eb3a9988fc7f1d53081bd7609bc1ff68b48f3738a22ef8e5a3a3200abdb0853da69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9779e68dd890c0f9c77ff9cccd41371241598f621978236686164e2aac2ff8418c5a57154ac62f2d3b523dd2dcd9b8d7529f3ee61b8bd30e3bcb6755809bc16b9c042fbc5acd48668cb9c6c455b27c267283f4f87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23d640c1087b06e3586c41c547d51ef4c3a07834194df598d4de9eb64c7318d9793a6ab421f4e64c0f0114f5bc46a2f1fdbbaeec90ce12c17b98aa8d5ab3ae34fe245ebb214f765520b7e98e4e26c719366b9421c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7805ca7a558d772265983b6c2ed0791590540da5c24f583693a3182b63553888b469336892ed96e283a1d82e22cddabe12e6b4ef294702e751367327fd6296992ebec10832c7f66c8f5e0dd69ea1a9b4a6fdd9733;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he36ed86c038b69d56d5777a411473bb85211620e2cfceb69daf8a95b9a4119a72e9cced950f4d6fa9f12075593388aa2d78ae08db54308b5b561cc9f8dcd742ede0791c6cfee7bb027203d939b2e3f568baab4f8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78241a0e1f743523108472c0e8fe0e13b09a016bc78e9a2ae5e0b01a6c88cf372cbdcee8c98b2f053306685d2c52f922a2e3d9f60f27e31528a5d122c75eda187039b7b91c7da46a40dd511f936eb973da6b3c9c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35194f6eba90965922af7a295f58c195a2456f5de9100b6b7351d28ed2477f64f3fa5947177093b5f6a455eae1172cfb8aecb43d0e7bef691a2f6f2c305b2bccbdbbe275b5638a20c57e3092ff3f2a94dd69c8033;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2dac66488924a74e9db583be1b504d70663e87e726a9431552e3e13d280bea1217645b4e7efc0a5516ac908bf582ae821e446885e6614652474737873d0d047856250024c47eff5b9169d22f150f31cc15badb5f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2ce4512e47ba23e362d2e560736092d577d195aa194e163feca4f1332449a084688ed810f17ce0899998a599a652d7d7aec53adabb3e24ace4dda7945dd6c2ccc569a3934dea5ee100547a44555befb631153430;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e1f9b1cab311a0165d764bdb95315b72c9790320e8532177060a6123b8487179a67500cf7e1d3b0adf8af3fd2d73cc5abca09d6f3abaee5387e3f052f0176e7cd532c1e750ceb87babd273a5e1e3372f24b35900;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80af46622ca88ca4c845ff7c5868b31f7241f24eb6cb1b90657137c35def4e22be4730af79a8598298f16ed15fc36b0b2954aac0cbb750efd0d52be9158df67cd599898bef9caca420e2e1fd1d40b85540a2409e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55c922e1fb95807ffbda523d933b8da97f3b87ad8185c148676fd3293fbe111b799e5156eb32cee4ce2788d90367fd0d2d2fbffb093fef66663c8fc42542e56d363873099667ab54a64abb56017da4b43d1318b54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed90136c41d06f8786c239d9ddac7aab5bac573f04db5cc694c4c0aca8b914ca5e89f292adc6f9ccd8ae554420a7fc6c9c7a4382450219c3bf2c0af992d01d694615b3a8a24aa4bd075d83dc66819a9e25daf90c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6d8027cc14ae82cb197f796d3e302132b4470588d492a0aa83a0032fac7640ee9925db8e9d912fd99b6ceb24efb45d359c4596ebfb1ddb63388a1128b2459147f2faf803a52ff91b42f2affbff24ee86556a9e33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb534a8f8a36f0fcfb36b39b9d65106f268d1d99c4849ae22c75a5fb380aa0427b2c9225099686f27d4a6047deea517951936581ca4813082a75f2058312f48f7c9090c7e3c86b25c1798fe0ed3dc74dc202051f06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha723d457e9dadf3acd98d24c2f2fc852b1648b10e7d6bf4796056d66159f8721a7e9c1f7a6cfd06e2601a79c00c2dd64e79f08edc3158b85cff6cde5e05cef49ad7f40cf4402cad52dc513bc5f06ac470034d51d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f7e88dae6f1d20449a63d6e7f570cce0a56f74c07bea5c9bf3219f5a35eea2c7ca5ae714541f2cf5aedfa8eb3089191f2cd5b9155fc53e9d181c4da225edc50e33a14b590cc78589c88fc39026a40582f39e2208;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81eb6f0b3efe040b0921abb3080b5685e518fc1e3502a0f3ef6c67ac7f22f5e789e772ee895efa63ab42bb858d269b85d68c2e5bb7ccda14f9c12e7b2ed919b5418b2b683861ea818b486224254d888d6a69b6721;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1bb06e77e0df732d34849ad27a4a7c526344274e18f0d8bf154c3306f21cbfd4cc3d04797aed0ccdbb609a85527c33feffdc9a8d918fb4408588302cd30a9c99e9933e20e77f0d152b23da6672f8990f7d342db2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h627623489e903277e5deb1172cfb303b893c8c043d07653078daa148dfd69d85370a016ad1a1997e4305e388dc49ee468b3e9501e40e0dc917ab43bdd1a1a701f96784cc1602832c6e65e0f83faffbed48b53415d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb98b3f89dab00f1bff27208acbefff6a285b5726273ecb53da1c1d2f28a6d333add42a866b85c42a99d73c0ec2c30d86908af8983506ae48b8b4697e493a26d92d1503b0003467e2aeeb4c242266d1e23cdf46a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d49956d29532a502e70dfd92d4560801a49ef2356c10cde8f962637d45ea1abb415a10b71f3b5b44d88688561e85cee9700618df99ae08e8caaac32edfbc21372baa73dc874f03007cbaf7f9f40a6cb1f83a2b1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2779a8c9266317e130333600b80dceb4e37dda001dd6d603bc54425f7bb6a224671159cf88a3b94da89d742769d08aa9593b73d0a9fc2d7ec64e5040c3159fe14af094477f27e1d3b085c06873f5bc912d5564799;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a9ac906481e7e1285cc1b55f7523064a3dd4f54623edc55b5d107720eff901438d8c1305d0b47d7e6eb2f6ce6e3d919402d5a06733dd8af579cc23a9a33a7452c978f8ca058b8235bbaa493c830a6cbe8aca12e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c06908565b034b3bef2c774dd245893d042eeb2c17989fbd6a18f86d88ea20d25173c39ad21644d8d82e6946e49f502b3b9fcce4968736dda3b65b453610e7c5567e664ced3377e4f719f321c203b32cb78005f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc05d365d4682ebc5c53a902edb8d11b92e56ad70c70c4d408e37daef087b1bd29dc287262c494d69cbbd653eee26a61f148707e0e31cc83502f99c5fc5d61b17aaf61a2fe63528b0a47b3e04aa650146ebe6a86f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee607db49562804770cb2328314a3350bfcb13dd0cc8a2a55e32f1e2f483338835f6b9d76ae3ecb7e1e74e1d0d9deec0e67e441845f773b747612c9e9db4ab828e6dd7af01cb9028abaade32587907ee687c62611;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67589ac55208db3c11075dd240f3dd0cb6c1b15530ebfbaa9ee858775881531f1512b99a4d1c559bb26783790b49e1a46a2d2a230d071ca8610916334bd50f2dcceb28f5a4e224837b9c092bcdce38710c8b2c7f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf90cd5b21005dee71f9c5cba737ff10910a67ff341f310b37d70ac35a5d1053398a1ec49e96ab8657b15fda37e3cbf6b6443bd55a54ddc489e2554e03bca862863f0bb24accd88cf31eb9a3e8e7420587920bdd1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53ecbcfafee1c298568bf616f97c65af0b0aba43772d3c5435a3480eed3c55ac95af91371731f642322fba720e1ce16e84b96892ab0dce8d4454d6dbb590e76e9927a09443482619067fd3cefc5f221ee43507f1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4f392b649c82383f39516b081b6a85a6ec929e75a73776fe2bced201dce9396e7192931d27863fc98a324707c40512c01883c382a0573dca40f499ec3f50ef0f799995a06e3273c075f1f06cf0b4f39e68631844;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac11a2cea69414df3a53ee76aba20d535aaf3bf24db08142e45c963a8f6cc615caad2a982aebe2404e12781cb8fcf80406fc23d487afb6edc90457c730e14cd9b74bfa7bc35043a8d707f4e1c581cde6a0dbff136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha702dc509f2b7cb99309552bc0fb19c61c299a9d755e6858c1088daa7e227ed80f01d36433fc0bb5153135b3a1499cffeb1c3d9f33c7b4972f38868a086caba56cebe38407f567225dc128cae3a9d54318a8f085f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc16afa065f28e274dafae62ae8cd1010280182fc08d09f1b961920d17906e19118c874575b8d2c1966a45b4113ab9ddd3a76845f4d957a5906b18f7dc64016d1bb86c6bd4af7288dd0fe0d7dbe77835fe93a37de5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed308653ebbaca08d01ee53fceed22362aa9dfa26cf6fc8c9609f9b0d9df741f8d967de74eb17bffc005313f587471f8b2307211f728bf3215d75ada488d497cdeb129131d6773efc7c97cea1eb03fb891c92cc7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he84592d7e4f0cc52f5019a84772d219531e6755a76b0e8e334695f7767024e3d537995c8ad09dee549b8203a90d33339c3c04c1ca7d29230b596b8865273927ba396f674d2d1c46fcba3d76808bfe6d2af53974d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5b769675bfd62aa24e08c18b6e7876720a497598a812952346bec5c265d5c23b3b28f760ea96504455aeb908f4fb85b2705ed7ed5c6d25a2712067340ec424ab909e8b3e6dde3524e3c4fbaabc43353b816e1758;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3b0d108e77f08ea148c2aa6c212d488dd3da50f27bbf642ec19fdf82b9cbbaca243e072807d7276210b1623976a478ae12a61e5e28ab2e6ea4d83b0f9e6f19c8410bd08850953a091400a9d3f71fd7168990ed45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3190720c33b476609c096532d98d44793e95f6fa0ac366af703cd157ab71f230dd8b438885f9265bedc779d9c9deb2efa7a77adee402de9f0e3bf4a58a489d1aec01e2396116f2da1ffb587afbdf7fb3acd6159f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25d07b0b3d1ce137ca750196fa49b27766ee0a9811de6d788857966d8a95d35636ad8a7a2ad76e8dae0961c763e1cde1c8cebb7adf9b8cc3a2f6b1c49afe4c51d04a1e23720e6cbeeaa6bbf62b95644248b30b218;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecd1cb6ce864ee1fd51bfa0acb23f61d7fcc8978b2b6686700277a2586a8f48a53c993754abe0a59c66f4c1a4214ad8b7526ba0d2dec7668f55448e4e7f7c28a96f7f89350f4d794adeb566b729101e558ddf9e8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b209bd931959e1cd3869d1adc47690dfcb842684d4f0d602c08e400939b2ad08557d47159888e4440ec45cb3123dcb9a0d59649341d88bcfa4d1e689a21243321fb46aa44fbf7ade51e195fc853d9f427b4343e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0ad0db970dd1ef2ccddeb2a8b73445d1891b6c818a115a6cf92b212fb86d7a61c2f3a3e8ed07b6d3ef6e2729a69ca0b869b98e6817e62c3e6d8089dd81be65894d901fb27052f6f43186eb0416a393ec2eac05b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e3fe75c44be93638ae18e2707b117ff5adefd794b1d5a50da421e1111b8e4910ffee3547ed6ae069d095e4390d5c4bbb2ad33afe191927e4eadec1e0c93b0b5509b7a7688efed5b1acb58e3c233fc207f99db999;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6907164a5224af4ed000944dca1f0d6507c561fe21045ffced483a80b0eff2e8dfd85303e608a7243117c583978b8be83a67fcb2519c83ed86b9d367c78c42c31e0e3b188fe1de726a812571f0a4ecff5710eb0cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85dffe00a80ed4f33699031fdd3cc63291a70a1127cf68535958f00bbb9ef22a45b58e08b5380b722d366979ae2da449b50f3b9324ea76b377cc0d5eb65eb1b4ce3da6382bbad51b5b91506dc2e8b53dee4ad36e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55972dc21705a3b50aeb52abf855e857e5f77b37b8eafeea3b37ed3f4f774ecbaeec6319be89b82ec90eaa3c13daaa8d01798af20789f9fc6e99adc1958cc190bdcfcfb247277742f945adbbe5f3ce6a86f784e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab10d854a25aef255a623cc503660ccf66fc51113988c772db5345f90fcd82f26a3b8569c4fb475ec4ded152dc22214db6aa9042efb9caf43aa6598e5fb98fbad2d04cd8c891edec7c77bd69ef6a9db8f21759fc4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h987b5d92b50448ca36f92751c4c28b02107a8b5560dc218a1ca019a3ca5f1e684c5c3bf49bdecce44739fa020cbceaf0e8844d520b2500203749e454b79d8cd795cf9b4c34326375f920ecbc89a9eab9ee751139d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3560790555069804ea7a98ec54bc7d64516a62c65da3d72b86ce30c4441980fd97ccfeecc79beead4b7b281c119c79e8a9cfbc5de6af4a31ff6af350a69d43d5b22ee3e8f862eac39404b032bfe9d5217f474bee7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h520eafc9782078794818c64825ccd20f2f5623a4285a4548d55d4e6b69e18943f2faa6ede81ddf6adaf91b6ada9432af2075cb6a751db7ccc16ac0137acaba355bbc0c6249201bb8c8701ee83fd15f2d89052196;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha02780abb6fa23af15cf4cdb3e9f10187f1407c115b84f7936eca386d510179e6cd012d8e3fa077d3b6d9bf5e64365873b75fba57b191c434b2c027cbc50ab78311c09eea7a2d07b4d93da4a73814aa043b18a67f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h343f76daf0170e7ed03e114ddfee818b4333aec47c5b5679d5b6f8073bb9be56f999082f7dbe0c1db5cba007af9db9978cc9b51485dff201d3bb1b62c982d41a451d483244412be7c678de56b05fc8ab7c22baf60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13437438b3962a92d4b97ee4dd1f920e29e0dd38218a47306d4ae9472c6c5a4984a75a43b30a4e240970bf91e2bc4775887ffad1a98db4cdde591771217a8f9bf1b0ef0d3cac237848c2cc7de00e2cfcfa7a78488;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56c0e80113e5912aaafb1f4039892f9b3ada105de53b5d0020ddac4edfdf1fc4796bd1d2527ee6c129ca08ddec0de3ee6a38df804c350dae7b1aa9d8ade9117e668e891fa46ade5b94710d41e491283dae4ec9b7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h458b4850865b010be5ddf786ef7aead947af121d179a473acc4d15fded6036fa6468dc9496376b4ee57dcd12c40234f2020fc9ebf6703fb428bb8b2eea39adbe4f2ef09753a86b21de4b0bea69140e7e6e8a71c2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29bc2cc7fbc4f8cd7bd724390b9d145945f66460472ef7aa6686219eb3f21201ffbe8c86aec3197141aea82bf1185e41deb897f2a5a61cd6d66757e8761f44786b0aebcbc52c4406836755e40f1560ed1512b70f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4ca7d0ff8fdec02e166ca9b04aae6d4d012c890a0f69c9b63ff2cab4dbd7e0ac0b497c5e0235fc9c8b3c943edaccc7da260178e5831ce348c16319556618928b64043cc360a002c3278baab45a0d5d99ab546ad7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80a96051f1e2c67f5e2b149132122fb6d167e382fa610a0f774a17ecf6831c39155e5bc7ab336cbbb3c471aff09f710b83fbf96bb2d16eac78995de136ede8e86082e81f364bfdada92ea16d0706cbbed3a40775e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d56784743f060eb373b4cf513aa4bb8d25afe8f75eccb82c802fee4f801287be2e00963bc10730e6d1ed3b42b4421beff1db94821d288722979ecdb7e75c243fd13ddef71bc85dd88f18a33c09c01e81fe6cb670;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13c50983c9d25b05f07a5fbc0abd425f10197011ed0b9baa2bb59dddf16d619bcb353b1a23bc0d4ffc44e51e42c0f3e0cda95bb8f2765003a7059045da0f8f96f2222831d4ca85fad2fa05edfade53ed7c1294fbc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h194f1605d4b3780e7a70c00f703d6c29f6f121975f24a3bd82849dd19b3aa328287a4bdd79de685cdcc93f5bf463048a3fbe290ec2c5f280548fdd1da8bc61ad096b54091f37148b3823d24f1f0afdb57e381ef8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h702f5788d17db20b5d209fcb3dc85fb34776c018dcb3621220a16b5446796c8320eaa394f872e1082cd7d20b1c7edb0b1c1fb425950894ee42667461f857643a72c0782cd6b2261947cbcbd824b300feb7df7f882;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83962202b21c1d9c3fb751f5a3391154d94802284c8427aec27bb03a328bac966a6f81b9535727220666224b50886aeb758368f405835ca0732f27fff7536d0da7966b2b22619daa2f87eb1caf8c138266280d3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d91789b6679a9040f5449fcc9ce69dd2691a10e07f2a19d23c70506a4d56f39ff418c4cdc81c0758cbb687e3bd9a9cef2d5f027aa7fc4678a9e5f72ce289408ea8e6108df2839a671f8a296769de77c65e5efca3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h270cfdf46911371059f97d4ee1c4b0c28c2ca559e5cc32d0611d51e69c44a094c7751ef1aad9315179dc01eb1f10c58d58d8c10c5a8a1ccbc6cfc0f967450dbc9f4057b8170209f757b2b6ca2e4652a7f65e8d5fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd31f6cac82d5a6efb858f176f96b155005b127ab021887de806a6ebd581964da74ef2027b239dcca0e0eba803a124a30338222b6d5ade4f542d5193b9ba24925f55fb49603531153f3c3b2c95241978d320836872;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he70545a5ce52404291014dbc525da77b1964a7bc67fef3e042117fe3ef0bd0d36b193d07caa79f125c5ca590051900959283b0fb59f2b3f10793cff03d7cf39446e6d9e3aa28c32bd0dd8d7da1af5b20cbaccab12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77a6f7d6d76cd9f6c1911570a9eb29b0d204408953c18c6e4c68a79269ea2a25d0a6512547081b1325047bf12f183032ee23cbda60b4e9ff9bf4d500cd237316a3ed1abadaf697c580a417de0700cb13481541e34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34407895396e7cfebef9a56366dadd21a38b002f1d48e355442a0f4d328418987ba91127e5abd25ccee82b1ac771ee59016210df3068e9ce902ff0a42532e83bcae325c2b78416a5b3095021f4740c3e366f1f9e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88b45899794d413a5653c6287483545efe3b1285ad3accab3d3b0229657b297ec9028aae6d40bd3cb911496d782764654cb5615fafacf8b0cee0758d4aafa6a8131874c2b716184dba51a82a3fc44da85983f6d85;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2436a10ee7763ea148b539faa1b1741dbf707356545031c1db1cfd26d6e41c231c8c3dbf8384a8090dae2c3436909938af7b818cc3bdd0275f8d45330c631d67f42ccacb74d14d9450223a6381e5bd99afcd7aed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e33c976f2ec34de14a53541401e6c69b5a01200854f6148fbd4cb4969b131684bdf02795566b07399311ec166ecde2a3eb09a6978d9747e825739c8c450314578a5265b8ec05f8c27486a42214f36b9db66ca83c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37f2984cc1af3fcf35406e75c64eee660f5f2feb50d3c8d2ab698507b2b8cc57ab349d48b03638de2642ebf615bc0a5fa8be582880f1f569f1c7e9db86b04a466a87a6e6b7c03c6e81f316cbc211f0e9bc3d947ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bbc0573cc430bc8e31a1fef3ebbf99f47f181aa281aa2c724dd08901bf443e3991ca98be0b3a94fefe03010ae3ad6ace936988fc2a44eb5d1a78cce4edc1d2edaefaa2adf355cc6697038a2ae4a156317352aee1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha67a109424214dd4a4de658f6600cfa8cffe9eb8d86023916765ab2bd72d87c5ca8f54e60d1c5f18f4cba1c2b9a1af5a4767b6d00e4e2d589159483636c7a105f0cb1ce206c07ee8a206ec1a7f063212ab78dea3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfff4729adefd9288e3c02d522e3d9e2ea2a699c4b546c8034d9d8605a2a1f9f0077e8c631a5f447ff759de510b8d83143b4cd5c13065d9dbdaec031a757234096192660503543d68af3f9f09665de6e02f2065d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47a7a5ee3aa0a32b8d36dae48b081793fd52d16d5ad085e67abbb9f1189ff2cd10d14a263c2c88f66c99829122a413eca72ae5781148efc9e49c51da6fc908934b4df7b77d2b133a97219657ec0ced69f73879587;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18ff318edf78655e7cece6619317e5d699cfe6da2556615f2a47217692807de19c26decfff7ab9062c4f28622f6979fda8c8ad043f6b52878527fb1846f3d6a79b1a7db6ce622ce93f9b9c570809c3d89abd652c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba27f16608aab7fa2b1a0178ecefa93151e49f945432130e695f557b62912af2af3f015f803d2f4b75d45a1c55c3dcb42806f8474bcb97e7e33ca311d01cffb16d669ac7415b005ce36c84da47ca2871135c0004c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf410ce4c31f59b85bb75db44d6969506c647177edc7889133eade049f700a4b01d4e14222d191060ae91a39b6837ce38a5431ac9cf2339f00ff890d139d33252737460ff8db468f68bb4f0a8c1d4b1e2c52322c3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71f8dd0348779d1363e9541c5f13af4f2c24782891712eb3185664c105db563274be089e55d381e4fd217bb25376261388059c740b45781b28335721c9bfbeb8898e5f1255e366497eb5f80399084cb3bb725a4a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a9196bc293854ea3c72a6ca00232ad6eeeccce9cd649d67c21c4d61f063dab6543e722a569893dd9b2700534002e5828a3dd763b4729ac4a0b68bdb50bc0f9e30397d89cad35828f322d3c7fca76e24d9a724ae5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1016d80db6f7613f284f84c29df710512e411ef3a605a00018ca75ad606f055bd9dac39d1359bccc96d1c5df4ee2a74dcaefac0a733a94a123d180fe6a171cfa180eb2400d2167d5c2c67606b595ff04a15ed2e19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h818fcd6ec6e8227d0c372883f97309aa0ecbed6a71e2b411844ec18446fa3390730c4d957da1f511191eb338dca501f1e4b3f1e9d9729bec0e2d246ecd34b853c91ae30ecf8e4da4e05face181f8175f4efcda8c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadcdf49b12e0953dd70fb8f4d482939438da383e337c87a7fa75032b535261e1eb033a5fcdbe76b0933d86889eeaa5ca3e1aa2245d4c3d259c7c1f3d9958ea0cfdb20c51f3fe6ae19361ce93398c82696441abe24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h468481e4524fa7a83d41f34f653cddf07f2f93a21e88e0ae9b352239789e6c55e0d18e4080264764173068d3349eeaaf22e1b17de8afab232cd5bade7f52edaaf335e20a3115d822dea7f5e0a64c34debe00580a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c6085995efd9223dfcf0d71ac4a34f54583aff4962ef60d31c5435ce388c75064cec548a21bffa45cc3a1009c1eb3c28a4f8e88f95550235f72159f2020b8674ba336222bf54951b8ecc84fda0d3ec5ef72aa702;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6a69716abe6cf8e930814261f851d1bc57f762736fe80331421aba346be4a20789093407d8b9177e39e2b623cd696a0cc6fde5fed90a4d1283ee85ff012c35387bd21629d61956289fa285f910f7bc0b12e01a78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbeb7ae5955ccb8bfae73a7a9bf16ad4f3a9bb6c22d489b62f394426a14c76cc4e2dbb9394e996165b9a8e5680576f3340ca56e4b18514b5cc7a971b05248703789996f7516b121432980d13de986eda6ee5e06a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51eb3b3a1317fed310e2f9c5d2879c97d895d4480f1af4141afc44adcc334e10b39d26c76e5a49f58ac33814b963c7f3c03f98d351796dd48548386de83bef22b0dbac8fc6b5caa70ad6d8a336c84ee14e7aade3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf153082a7a5bdc44744cf0ad172eb6922fe9aa82b4d6cdea0ca68bcbdfcaf0952f53aeb16b02fe62592a4408e6f39fb5d09fe13d264e9b24a913b0e4e1fba6297b764109b3de1d7963ed2fef986e5e3ad5a893b36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba2684863d850baaeed015df986b8411c0c612e8b36288373792f04d80e5bc0e4e8b8f91db3b813fd96a088408fbb9f91b776138a8db85e4bcf243180c21d9495df2b804dabd087755ce63a2d5bfb20fa88b9b6df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd08047f01e93c77b3110611109f447b8ba1603c640204c76feb262d4f882189971333a1332cf32d2e38f382813e37f21eb2c3cb8c0f01d58bba43026f914a2bdf7b06810c593cd18f47196ec257c5472564af21d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd30a500c0d8d84af65452233ab68b55610f95f2480f0304be0dfd32ad4ba762651db5763f6b1e297e807dfde0cf840d4d20552e4896078a8542c70e089a373b069d1fdce2ebf0b6dd7efc1144efa30554f4116ca7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4ef5bbcc8881de3c59a65cf0e60af51403aaf4931af8afdb5ef6d9423edba08e606411dcfa572a837fccd78177a04b4ab08f3f08682607c5c050a43bc02d125f27fc8338ffc33c80689e996f06b7b54d20a0bf98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfb9862a9272877c2d5f783413892346698c6c46916384d6f9439e6546447d1e398902327f04f95e1800f43cb9af101ff16887cd08f4e7c0b98d7da2a4621196a0612722a46a8774c8108fd41199c3ad2baaca778;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f293710d92818f4da6cc940796a52dd325a819b33653f9e193f13792a51217bb1abd9a58c9d40843a70d5e9aabc4ee22bdf68d5fc9c5877a732b92766a3d65a3266c25dd7fe6169a97922dd825a456eb4f0f452a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7b60e40c17b47e21d47a27bdddcd61ef90ef1eefbaf261a20beaf1f75629c666103503dc144b30ad714b0cb3e04e9c51554a77f51fcd6020cd9dbe9d9aef0f43ef45a6c4389a559fecef5c5252bef1780a457e29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e00604366907ec29e02e11682e5c46d3f7724c420cd88c710982a9e218d2eac22d71c847d7bbaf1af11c6481ef90483efbec23cd981b86e51fb064e3e8fc512cc9ea005737dbe0f099e75912a08fd29d72100eea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcc5cab267b8406915bed9c96d49d09da44f7adfed42c7c1f6b862598b723d171a3bbd93ac3cbd6b6d0275c80983bc0d40c7c008dffb5a1095892626e7bf474300482f3bee0f3732051d0151124d0177adf7f266c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b7022bda81e39145d7952642a565eed445eac1558281175c25ef9f432490545f80ecfcf02a31ac6083a00b68060208db8ee2be0a95d8589e1c2348d6bc0f76e189f440406f135db96ef3cc32d93707ad2c6ec74c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cca76c79d38dc04b420858b7b3288c84aa131b1e733de207201554bdc58fe61d0b641abe5ccde66869496b88faef25603de322cbe56e1da118f5103fce1e629f5e545e0823862235ea10786334bac7b08dcdcba3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heac9e0bfb07d72626d6c20555a2f694989e6fa091d45abe05ecdc2b8bf0bb3e17de35d1b56af929dab7a3443445ee33ed17773df021183c038a9655e9629c5de23ffa095ec6e5ba92e050c4e2b6b8843d16b8fe51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66f0db857491f527a1fb9a59a75e7df4412187c1af22b8fd0cc34a5fcaf25950d28f6eb89d7a3cd49c98341c47c7011e71208348aba832c57dfe70f3f5e7905a6ebd6b0e39deeb4731208d0b7583e1473f14a9049;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44cf01a5aa35a6a0794d56f705018d0db7c424d269df396cb4614dfc429eadf5c6a3473133837202e9ffd2c235ef5f84d6028665bb3a9f69c53e9c3255cfd92f201b600181891df08fef82109fa4c48fc90d806b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h725c984f34c8fa286f32075e60cac8125968d87130536251efd729822bbb290ba3497d97105741816dccdd8f979a961a7735756d3f16be3cfb94fa61fd6f2a5ef30f1e22b6dd83a67d60c156b4287646cbf5656c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h688296cb0f62d01b7ee464f702a6579fc9fd21e9c602852473c09aa9266b0ada4f9ee3f9c580b42d4a16bf98760171716961064d2c40bf11d99ab9e65455350ffd1260fdcf3eeb2c6cc956140a341ad7010c42f98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb904ad25714d3f29fafbd8e9d60424e7975c01f6541a69f93e62b6ae5497626a92cc201f0ad5af139858259f97286b5fdc22e937c8e180959375398960123341f41b27cfa85279f4966d29ea252a4d5aa1b234fc4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5db7a7c1742521b6ae02d770f2cdaf59cb6c7f6441e11acd7ba2e17947ff6c854a515ed0923f5a49c76dff46f38eed1ebf253c21ee7c5b0d2691ea84314e3001a946c1b12617245c9cdad06d0728a7196bd671b71;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c54b58f21b19d460bfd1262443d0e59b8988fe4f48dbd4e86ff17e2c964d4781a2609b14b584c4d5926eacb2a7d5d54af23707011269ceb90a49c5b8fac04383ff280d5b92eeff47830a8cb0f7178754a3ab3f00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0220fff8c74bffa2c54a6e6c422f0901e905a6e99da9e9b1227668fe14754263d1ea110e1e065d9f47afeb40658a3ffc7f1351e1cea6a6c757f823f600adb677cd53db0eb2ce830e7027d3f3df7d894318b2e505;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72db7fc396ebb79ffe3c0511a42d25010949da650cfe89a19617ef25531ac8b06f26879ae90023ca3b8eda078e61398ad147459ac8dad95a1ef4c9c4cc78d0ba98b588c6d67c4b2d07376466ba370c70acdb787cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56ecf7cdd984118b3868cc669091ba1891187f05890d1597f667c540a2b8f635a995a73831831a7999c52b6d68344feae33d6144ddcefe54160a4f20a3ebef36bb94c360eaf36d0586c132e19203e50b57896aa88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h412449b6f9eade7cec06cf33eb8a2e438a5b5dad8257e20099008ff50fe7642a1ac17e726c93ce5a9ad3e12bfa801306677d3a6c0711dabd7700a0e5f54645c2ec961bbbaf0ed88c9f651393ebece570c68c263ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19130c683689877448321eca3a7fd7b5f9589e552400ac51c78c222e6cac7052cdcab3b93f08cb80541ec8ce588fca57512fb54c542c9da3546a446affa6bfc86e3ffc08f944c76aed2b19fb91e4d49e588aa4652;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda653e7ce87b1ce2bad7903e4f273700d335375f7f59f7e469d0419ab0fa82d76bc1f3f39c6bc455b235c3108ebc59fc713bfb890c23ac1b24f167c12dec3315d14dc63838b75092d374d624216ace8dcca28c2ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43cd1e8b9e49748d120c0c4ba6e4c40457aef6e5267d79958c4552d23c40f2ed4b584119b4d1f493a44ebd80e69a5984294bb19a5bcbb23a56cd86c1850d5e2dc8555a90a05e2d6bb2a12d8f5fd6a01a77e9328e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7142a60e35870ca746902e6500fd4205f81819df57413c1c3e055d2db2bee89ecc985036c1ca12a21b804f4ef2dd8cc8a9ae56f51656e800c8a81dab5f9468b46054b608eabd29c9ff6b7da512485ca3e119bba3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48a5f15ef1cef96bd4a13003ccee8fa64fbded851af4fcbb9d4f142c7aed24928e1d9ef266334a99747d070116d480ab8954ed1f0d3c0229bdbdab29b7d4ff414debb113d40024b6b4a047a2a589e70f8770bd49a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8685d8f984e45eeb86df6de9811245e98713d90ed5880f68f8a3ef2934e62a75dbb5eea49b91c099f1588976525778d5a1bf7c5d53b831e707c04cb7df67f651dd92fec6f3b71cb18c6b226874940a6eed8c3316f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he584a676d0eaaf3ad692fe910ddef5cb866744654cadcea728630f8a8f3550ecbd1af03015bebb1052831302ac46033220686108dbd43491ebfad0a15e9162ccf004b510ac854d10bbae5cdcaffbfb28f73e7849;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf51882b422991daf1ad6cd640f2f3df17da6a2de87b5aa53ddddf2cc0e6b945e4f23b8f90b3e23e82e68def4e69e08d49f630e214f48b846c45ee339df3adb0efadf913b3e699293247ee09c7a57f4f57a69167bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c349ac8ba13c4a240bbeb40768646135f045bb133eed4d0e4a77460b74e69641f64aa13a1cf8f0ae10f6f759118afc0a5763fbc0291b9faa4ec39bc57febc0617c28cfe22ed1d8a5057b916eb019ce506011699f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23285bfac0caf3df88d01e36a2b02e33e9dafc37b19c9f435823354567649ff35d2f73ccd5b3902b65bda3cb31c64e7609c6eea0956fc2dd2e74aa6a59432af72b39d0a1bc4a7e0ffb27a2de4a5a15ac922dff8bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fb450d6447c89fca9d97729c7e55b912884f381d69c4f0729d091f649ce2703c031381a8dab6e0b7986d313fcb6ce73510b53c938ea5b8eac158f4d2d71a3864a277ed4450a08ef669f6829c41c79a2d027eb3a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1e9fea3851437a34d0e881cc1f1b1c6184b183f57901bdd6f409f1ff4147315720aefc4b2fe7a3de485a65f7733db9b6aff54ab2ab5f67f8c58b48910c886c4bb01ba7d6abce2bbc01d586bd93839fde84bd00cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9dfa000915e4e6f4b2ca4acfe8313385033ab54f30cfc67841315f0715f0d3a7297dadefc8887373f7b189a90409d0bfb27c1d63059e6909a7d9b088785372ae8cfecb5530c7aa90a7517d604c9377c03d75ce48;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h449a7537ae0460eebf718225ec525e4eebabb3113c422108c6a938b6242353c007f8afc0c8b31ad2fe7eb46a05383d74c5b48e92e36b729873e43088f52ab823f682dbc7b3b4278082a85c90344aab9f940dadb7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c4ede08d4559f504e9a3e7c7933de3aaae21cc395dd742711717134ff60ea2977a6645747bf3ee66460f83ef13ed81097e352c40a58d0803205961401f0488f6c00b8b5cd077321f750460ddc25a7592d3a858d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7330c7e2e5af3b8ae583d5eb6df45eacc38db3d81917a3e41e51ca2b34d1b0cbe775a72ab0093c9cae6e3aa23520b1724217908ddc29857bfd8737854ec6749982deb993bdfb74224a3f6037d97c99b8dbcf48e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3381a44e29c962512e6c63339d555bac217e9dd198f0341ce547a4b8b0453616418afcd0af5e605940cda40d006552b5e6c8561ddbdda5e87c6f9c8234c1ca1d6d971868ee400d7ff7905dd21341fcf1e72a175d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67aca95e81a213784ee0dc734e94114c74a39e709d5dda162953537d8540d0723b9d7f06837ba21394cb4405a65e38d382ee868112e0c025b9ced11453b01058778ac6a5d70c1f1bcd5e9358e141b9fbf28b749c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43c79933d038c2a0182f0ce636d45939a03b393f9fca88a318a88036de5042f8607017aa1b71c2b79834e82f4deae5eac96bcc487af45165f68a0d6868fd1e0b76aff57ae6181b5da36910ee78a0f9fe1b41745fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h796329d05c960f2f1f10b34395b6ef5bb9ed70542a85cea86234b16e4d9a79c34ddb3ae458eefadd3bea12e8698ffd091c1588708ce09f3d9e10d2eae45817c7b1d911ae8330cc635c50b4a7b0b5b71ff52b7391f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2365c2f8d7bc29559498c31ad32dbd4f94454ec04db83d0b3d10603a0ccce7d6166394b47b597cd065011e27d451cfbabb9c52ea00fa5f4f80ac0097b0e04bbcc90de642675aee2b7e0219fc099cdeb6f7d18ca0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb3048882e05d15fd44791e487933fa8e55c81835a3185bc28daaf7a4fdce1ba483e5ecdc4d5d0f4e0ebfd53b66b97a4755055e0dc2bbb2b085f580066b58450b9413719c8fc398f59916cb358f8bae2274834011;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82f3ab90c73d9c7f6b689693cb93985bfdfeb252e0d966cb034f890d9296d1541de321a4a86e6af7c0cc333c7f31ab61263c60d211f13b4cff9b30422d2dabe3f2fe371e8ca7a3895a1b501301bd57ff517c2116d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aa650cc2bda347b5478d42192f7fd0f3ca8bc66c2c17161c69c4aced931247e27747edf58637a13933e4ffca70dcf87245481067323939b83abefee34e35cd422252660fb92a014a1d97f55fcb8bd539d41e9494;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha05b31671cb94daa407c8ceb3fe2b39d522f12b6df96dc20b1b9dbb0e7c6a1a47b52871ac7f1e0333694e1042762124ff66f7e10e36848d8c9617e5c8eeaec2bd457d66b2c2d22176706b43e5699d7cf65d34d2e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3531108959abc76b9f3a59929cbbec9f87222cf3465a4b95b6e6fd5287ed06837e6d6b60e9c0e3a6a445993affc4847a84aa744a6ce39d0afd7bbbfbe1f596965594f5cc6fa2671f070a6b175bb9f5a4c75a5a69b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5614c00850dc87b990f623d8ebbf21ecebd94460b4ec89c642071f6441570d00bbbc3cc14613e888652ff49f228d91fc1c6ae8c02c67e96f779e1ff0edcf5d3be2a53589d59a8bde7418674cf5be7ca3b959dafc8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5285590499cd251c1d2d0f2e920ddcafd0588132b933309645e147d067276bf4e821308f2c0cf7e4ba123e68faace6f725a5760b3d1c6f0e9528e7ab2a7cefc6f6b9dbf93aac47e5dc8f9cc2b0f20e1ad6ede422;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8488c6ef4de2b31b521cd8589afda2331e23281ada9e8acde291f2625f633ad04d3ef473badb0690ece0cf5bf53f676991788626ac9d9301c909a354b393ecb08c8f15c7de1d3b240a867793107a9181992a80966;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5d88d622e77e535edccbe82e2b2f66341875bfca62338fdb2d683dd906f32783c6ead0f46a183cf34c182ab3aaccfd478f0734dd0c2e675e671831584620fb426cadbaf2374b0b8e67bfbd8c96972d331f822fe9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc34a59e77606a2b3b1be8ea2d81744cf08b76d4b6832b66730e745e6fef20893d94842c5b2a859aa5e3620ed7ec97b0408c075ef928656bfdd2baf5c06ecf88edaf7fc66a4ce0bb105f865769861c3cad147c2780;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h511bc93822cbd204002d3c2e97c4854bc2af6a0d0a7f1a4958ac6c034bd14372383df9c0965b4bc3eade73cfbaaa55629d1ba9111e40878a9325623d5504b41f2ab35828eaacb5090345490313689ecb2f39af3aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c100f78fb6868c8cb5552b7ceeabd280557f84153327234264ee9aa065a780b606783ebcf938cc1122969630202f6d9f239f90b0ac157f4dfb894212bc15ba19578bf8a941fe0d427d2618a706338bc2de0926f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85480ceed35cd3fd1bd6e77d6488ffaaaf7549a1d74d05272ffb200f89904cbfa7304e31acd5102dd32b99c8580161132aa6fde642cc2640651385ad5cb469dcd0876b3fecabbfa70c2c52bea123543b102288d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haea1efdec0295973d39708231bc36831aaa683c0cb5a22a92d6ffaad5867dc92b0556276b38bbd0f64499e45e7a6033d30576314f5435e7ce673b3ed65dfdb0af76d7571f4c7c1b98bc25fde853829749b77c580c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h626baa971d16724c527238a2a005f0bf82cc83ada4cab4da79da483afa3ae4677e5e7a68e478bacb07c693fdf1e2553994ca587ef9b2a358b73cb2e923052459ae406f01d2e56d742c3f50417f52d786dd12c2e47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h660599cfea31f6bcbedb25210518b1fa60cbe1af0085fb58019b9b4e19a09c95e583e76157429e23b942f9b4027c8a39b3e6b020609e2d7d02f9827948afe90c6daf4aa470e7f5975205e9253922ef38bcc837ad7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4a6dde73c64ad092608d270b86e7fafac8f96a998f16a045ff7756b3e503fda9fe4eadc2cdd15c84c39cef1f2192643deaf4609f239e7ef6fee8b912a277834be90ddf7c8e04995b54a792dff8bf783562ccc032;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d6ffd4730ef518c4d121fe04d000bfcc1f60212eb72ed846594495023267194faac39442dc5ce9d18876bde9e919c835c6221ceb4dca1608af76cf95edf50b121026e3e39e3f8a2b25d4ccf0f872637515041f74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf792dcbf9351594f14c10e7eb669acc4b49e71ea86c5e69fe8c8818251398097469d7ad8a142ef85232b5d508b37fac5110a6c07f82f8946cda35c942c66e51b9547fc055c46037051aaf4b17cf64bc3d00b2c56b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1780b3314e7b296b2d4d37bd4b76ef2a12db60c4f28a1a788e840eea6b1c8f3b59ded4a6e44db9a9b28e9ea1672de3166b38b1c79a84274a7c10145635067abae54ba87769350d7c339256662279548db6afa2181;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha45d58e2f50a125e55b83fb421a3707f4262fc5bb2cdbcbbdb3d9622a0e0e20b42aca4120dcc74a6447e5611f3cef2fe5ee700f3d81718a12db9aa3935dfd048fc9a007f350748820098b8cceb146271e0431bf56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92a0fc0b019bad0579d0004d8af9f376677653a17296a6ed0d010fe59091f91072873249d1252e60b3a3aaa446bf05c8492ccaa5ba1afb91471ab81cd64f50168389bc633ab96fc6d9b3453ba6f47a0f164ffab8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h621e8af28e6309dac5a86b8487a691045b3ce9ca0e7a3fc75f09dc659ab5970f4eea54f459efad369e70c480ef27c5898aba6dab901ff17227b5c708d76c0183735484e8aa0895dbabc933bc65b59ea626b5a0b4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6913f346b630db4e221e0190aebe3ccc2b626e54bff550522185d02cb22f44b85fe216f5d9be6647497f9428b583cf21bb2392e50880dc74e5489f03340e52126fc88bcc84c44e2d322a27e89104ca3062b2cad2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c9b673dea322a460a9b785815d5b1e808f49dca947466023944f0c2bd049e843a963f15e0728f5b2f2c79e6f5b627f9efad63b016a4fd5da9b8c9399d6b138c21a6339548357e0326da251744c6e8d93c78a234d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba649b742c2010c5fea1103d352ce10a0ee20ba3eeb9438061a538d0ec38d3cf06575a006051480bf4fca408b1d7f378ddfb2bb084d0f51b91533c31201078a7b01d8f3e0e5b4255db4d52b6acfa0920dd4e98b22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd810283e32958ed7944f61f7f2de224f6c1ac6a3300bbe2e4242f62242d1217e4414c4dfd64d5221353a596907bfbb9eb1632267bf5ef66b152c4bbc0de514b4570542e85656e6071bccf9d6812ce1b22cce1d7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63667becb6ed790cacb6324d9d9c61f6863f7ae2a34a9a22f31d687a39a16179e1097bd2cb12f7b1f579e18443cd1ff3d3a1fa93b4879cb8895e58900dd7b56e6c2fe7ae45aa4943f863935543a8cf6437836b4d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7325acf8397833a54b88e88b967aeabcb3e887a3246cea64868cc701c8477a9c0bf7dbb9fe724a4160030a40781eb37598e877a4132b8f5068d0a9448728176b41b4aa22f0e0ab86889cd0eaf3443f3bd5cdc9596;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haba06ce9fea052375afbe303eb99d6900bfc7bc5bdf775f74052e4ffdc8e84dda09465580413d189a8a7d68f700edde7a70f4a6799d123cd60e4bbdc690812567a9812b1a8f5c0fb3b05fdb186e4d2ef09c7ec496;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf14d568d52e56da06de3ac5a8a9f0d845bba17f528f983d1ee83eabb1850010e9b744279e837df23226e8d3c04eead50066894a02e3303b582384bdbd91e441a76bc3051b88803b72f718f39a39121f2d6d9b1b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77e7cdbb8d9a33b611f32b6821bf0c0da89ff04d9f36ebb9030d262b059563935953bcd2c87d554f670adca67ea0a4845627829555d7bcba3216be1e82b684879ee2bf644120866e35ce1e25c6bfb8d98efb687a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95252adbab1085d85ab2d5720e02aef11e02e51e79298d6fb124dbee932790856e808f8bbad442c8b10eb5b0d7219a8f718ae74a038fd21c71ff6b87faad02f09c041b985e74535f6be250c0afda208a0b72c2b5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf57d0de1083471e57bc0e56f0519150f3602a06c9d3a064ad810c4d2b89f17254c574608f4756d704c0ba101fa598d4661d502f0cb21a79a6184923419a104a18b94c802ce6bfc4b478d6022b2aa140a2c7bb06d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4c62defd78b617ef04b3df2aaedc132e94c273eb2fadff61b4b47c7a77d375cf3023bb54e7ed69205413de667f4a55c4d07d40cdb281555d6b8e0d7f04734a52d2705f0b9a567cf48a0904053e141e55f7b8fee8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35e98bf3df87085d1a364edd657a9d459c63b6f93f6625bdb732008c1ba141b73d4a8d9c5e4e011bfa28d1ec697485f0191e06e7a81bcb64c9b7e65f910b15e9dba459cfbc380dee4a84c232eb033ccb6b82f00fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50005174daf3cc6f0b3912fea8af4113cf43cf26e8f71c913058e7dec7c3998017b284da2f8f722c507078186866caf5e4a54ca0e043049b2462aca29a281b210d53841c00a5ccc7ba77c34be9e84b7488962b5ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb82f895c2e720de2a057172a25223e051767612ee5d192144a8274bf69cdbdf213ee1d444b915a5fdbe09a8db1c10eb4ce4c52f1286a877aebe9cf696afbb856262f155c4bb9c7d265c6797300d65fa1a43f6145;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97290d02f794e9d1acbd53a4981a8be8343a845e45cf873863a8cd9ec6de7a3e81ee24a77a33b2f2053713ae6acf54121217c8caa625b3b5aed1d1076dc088584a3111c737829c6c9b0e659f49cc5256baf80b05a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c1f7fef9e6b9a4cc570c8c25d32c50e9e1ea8ca3b444b66ab3104567b618a40a80d56ddb9c07a8a7a39196f9ad65b0e16bb9d154e4eb2ae81338e9d8937df1e832031313486dc10659e7e5407d732084c2df8693;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4fe9abb7f5a5a79f531c0d4fb679db35e2f924c62fa15c26a2ada91ce637f32c4c5c70641c51bff6b050cc462184d7e4402b66bc4d451e0875d10d8cdf4220c84ce22ff9ba8eae70fd07b07020fd1eeeaeeb3bbc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3aeeb26b4494d33276e5f86eceeae334237d504340296d1303347897c361f3a7d3d7a98edc0cd2de11760051f1858406508e5a372b1164198b4558f4803091df25769f6e52f80e9611fd7a5570f23efd0840ca150;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedb9c6724e49ca5b5418c3228b9a4e4e1928b0cf09e7f73b248c62ad1f9fddebebfda7dd82c69bb532ea4580d8daa1c0052acf71234a11db19da4ab57cf819243ad177b97489ac00ddd53c13634939759dabeed73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac42070c23151f4efc21299847c8f477a7058a4cbb9bb291ed6428532233dd8a9da642cd0a7b53a2ebf58fe263e18ab11b719bf36c0343a35df9a278cd4312167285f0305bcbabff9918f3cb53a3e3d42a5860bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c4c92fe3bd0756efabbfb042fed9989b102074a39aae579e741fb099e46aeb74a2e9a2d9f2eb0dc0b3e2f851c5915b538aa3b66e1450df8daf5ddefc75ee123bebaaa1ed3a04bfed8ad8fa2af731de842efc9505;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he65aea3018a9dd34f62dae592aad22a1810e0c6cd155ce3d6786c114b8160fc16251d26785d2e21eb55538fda25613e534376aa67f2cf9f4dc6081684e11811f0fb7e7b1c6e872e0aa629956e1a70db6fe260f7f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7445b044026edc1b7b7cc77201c03bac33d81317edf6562db141083e64412ea9e1636ddcff501f0db3ac3ef9023e646e6c3a28d2d313cf1b3986280259b29da3e926b0a775b5eb87a101738247352cf34d10d4f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc22f7a391a533a4b8db48a2fa66a6bdb7cdb8c8fb108fbb99e2728c5a14f2bc9df00734e035e7fbc5ec04f38bf89940200bf5d676bfbd354a656f295b06366ffc643df1fc2ab9132f65e4cbfd7b81dc563f76547c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38a579aacf221e1fdfad9fc6390b3c7e7dadbf2699c6830eb3598596d2f418c3d2edc43927d3f5b3b72a42723c61348b4564fc7a9fbe3ac9dc166ef421a83c9f8ba080650638e0cf24eb9b1e99d0f7b8bd30b6d10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2368ee784a10c20b35a08f417bc59fe3f11bf9ada56d746081d4cea9be78af7af51887bd19580d60d265cd0d89c95e4450a7f1e96cc4c8cd4c2645ed38ebf1b8ce86ca2c85394cc6db8156d3af042f162e32ec793;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88b924514e1e74167d22613317eb8a5b0e5e02621476097ef2d8d9eefb9d58b4ee8480408f3fb0a7bc21bdbf5432ff3dc95a2e980085a6aae852bc28f2fc79421a10a0e2d2663631f23816f183780c56a0acb8099;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2950a54e0519c81cf0e27da80eeeed7986d0e2cc09964dfae5fe6d3c7e3b33650d454c1e2899bd1a20d697b59d037f44035a4e562cf3a26e2b1c4539f2c8dc733478eaa3a348336327d49346c5d30db088bb53e8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22b7ce0e8e38bfff8070e0101172160810ddf928b98ccf1673773f0e0da8177f7515481d0ca79a7b97a8ffb66d4e5467dd2fc9d9653d7d685afee4e20f8c214cfcfabafd9c02bd6583dc8868cf3ef8979692e6f6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4609aad9303ade329dfb397c5e3e00529cb35d67c693ffeb9f0ebc8c355340dd8633745a225b26aca1bcf2e5471b1c6fe51308050f09151cddb76597544106c69a3a9c1f156948fb57eb0d67de3282e9fb582e66b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb622fa4aca0754e380dd7a26b196b73cb1d306c77a32cb8acb55cfe2f681f10c2a2bb9ec12c67d266bd0ca803fe94ccec95f688af7fd43fe2cfd40a5a0f5ec2012fcca629d9bff89559caf7109b03490b395c3b96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ca67906c5f8799f3dd06e798bfaa154c04afbbd3a839a25230d246ea4492429a8bd9178fa6cd091f99cdcaa6842d0344d3939a48bcf43185ed0f8ca69b642f925df6b80e241b4715b8c43bc7a20e82a20b57367f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb108ffc993d62ab4dc4d615dbe3e6031c455dff27d9e7dbe4af51f59782f4adc03b27df4cc58a3b9cfa58d69c3283b057de72d6363b54cc2c05d4589644cb91c1e5467a327d98526b61c61e9bc54e630355a80236;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha69a9eb9787de0987d6cfae503c5c9b337ce9691c933961a3cff3a80ab9602317f00c534c1fc7d7f8fafa1f02c7245fa433ebb6f5077f3ef35c79bcdf80f0f85103ba692a2c6ab724e6b7771f2bf7a86aac38dfc2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50bf076c277ff7da4897d5f1cb66b5dc44e65f2a115b691d858a358541accfdbe2542bbbeee53ee07c9194088ad069447a7116c38eff65632d9fb037bb14f9c9e9fd5bceea701dd6e32420f96219da35b50aa7b90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39517132caef267731153422dfcd1342af8fecb470687a55aaa231408319e9d1c3ca68ed765109129ded2351e9601c759b8b9737b20030642d2e4d7dd2cc010589d80538a94f67c8f7348ed320d78656b5c29cc21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed6255c899abfbba80f6b9c964004da90407138f85a800b6799ba4823f0fbed545a0c1822474e21a7a5e4190bd3fb4f156ad34499833e53b03c7f586cbb68e2ffecbd2885f7a9c43aeadb801517cb2708742d5d53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d104c42fc3981be72ffc48e9cfb6f2ff18fb1f7d56921c992628e16e0d35a8138369f48859a726070ddb89ccc7739a2677e7bbfd90a9101b5425470aa9c7cfd5f83552849ede879fe7c5e61baad7221c495c6e25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4896dc220619610e03b4ed329d523358ef84701ec23eabebbd2c86df437837bb324093a5fe979468adf4977fe75cdeb1f6317ae69f0578b87a60d2f7454ee272715ac9b30951b7d337794521488aa8b415f46d37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5e3073782f1db72c0ba00b4d056bb2016c45d4da5e1d80776afe370bc676a4cacbeae434ba71301b72fdea9a451943f510ed18daac489165aee03a4c9a1bc172c8cc2576b6eab402e8e1de50841e1e1ca1c2645;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13e3ba73f829d6750ede9fa07c80ca4e23cabf99cd6f4a1185d41417065bf20fbc085bfecd79c70601149b9da0f4bd167a55f2a6400874279b53405441fa61ea93509b6324989375c5907d89a33a5b963f3a47cbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf5c5a63fff03af304a45be4e5823b4ada188e09f32fc54c2699fde0530a774049fe5d92be7d568d1f26f38075a23473cec1a4d4d8b22b876214d8fec0eb5aeff0bec108ea04b03dfe0911703d8949d19d74e2a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd90f2d69ab765854f8e5d1dbca24dff9f68ad151811d352601bb2314a9a6e09f33857977b8d4cb370c5e6dcdeef0a538d7cd1c2baba7b1f0c82464475f9723cc11cd5fc67c7d86923ec2bf6f33ca3b9a005dbf76b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64f36e84319be8bf44a20d9047dc0bfab5241f93d88ca6351a34b4f6dfffd752d57449d009d1175f80995eb8660e734110bb0abf05837002b2ec8806d8494629dc3166e5d16c2162d6c7b08e822d5111421b9a058;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca7e6b0c19c2aa3b27154f8d3bf1f1abc81b18608b2623586ff19adaa1a6c6a5600a49da91e992dfd879320e0fd026d0a9308da91416991c5b246797848eca55245ea33fa6675b0435d416183fc7fd3f66f2e1911;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc8250bbf71b14d6a44d1f7e04b9f0ccd7cbff071cb84d84fde475db8e8a0a14527281835d72a6c633960cccf17232725e38a3729062cc645fc4561feff198491e6b035ffb40b915cd15430f859ab15975f0cc787;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92cbdd119f62bd4944421e1d4c9e6b9eceeb98826d1fd26899756bf1e7d9ce39929c11b13d3c0f83dbcb2b3ad66942befe56ede2a6f72c5ef5a002f3b9b7d03fc46a4f1530b0926174c03924c12d947fe0b387d88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c5508eb5392b2303632677a26087603703e0ba13e6aedfef2d3476bb817843d6c3fba47287a4bc8adcec4c6a0d206534c4f59757befc7d112ef8076c8bfe56fd179636f4142a65d37006c917ee20fcee7fad8d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h344c6caf567b477c0c646da7b556c1f925e3f4e097ce248723fecefc8efc6329c8aebc02e6784b949510184141b6462547f687b2ba8ea30d9949d6192eb163fb0e85608d148c46c5c2edbf77b1e7351f2b1a3dec6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5b06cf5ffd56c9ba9203244dfc65ab40324db054a786d56529a868267d79cf45a5f85ed2082bcbe93395b011718a03878866baf65f21fbca0d87d7225517f7b84e0488daac379cadbdeebb73c5883db3ea667f9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6891693001c2f28f8d0c5eb66bfbeb1ed285440abc3dced0ef4dc05d6195e6347b72dce096cfe5562b5b42d471b6076751aca9038187cb8dbfcbab74c631fcbb8733e6d14a53ab3e3729601af68b794fb47d704;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1270f83d5ffbd02155c36b8b6fed87bb6efd8483284a548809c3209e3b6ca97137883ac6998a991126cbc8d6d70e737dfb88a91f436c05e02fa19871362f310d8d43afd070f96d890887a1010b03c37eb86839bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de6935ff572678d40776046a8a3827ab1d369b3bd22c465fb4bc086b1667257282ea9c5b2a30bd16567fd2fd746a2d10f21e4d88bfc2af7e3eca4d4ef81fe5674a82c74b5abaeb5229e86cb6092684c252d2b900;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f2bb77a2b02e6575d0c90892c557f73528cec1786b148b499cbbbceca23351bae6d5bb41a446a99c474032cdf8ac5f8a725b12bafb845a9c6b1289bd9ce8db1b545bd63925590bea2f001e29760d4cbaf3b75b6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa7c54791dc6f89b039049b0039c538a9211628dad79eb7a5ac9895b09ccc96dad8ecfa9a3a3669e6ce922554955e0f83f1be4f74698eed97267aa17f8cd142f758108777731fe94dea278507966ac1c1e9e516a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h722138df914a75965603150584931922c887a41cf10a39b8c65fe966cce4abb59ba7557b245b3e97a41672aa449d1c440d741b5154e9e741a16ae83206959e05b4e10d2eaf9504b188de79df103a321555456c835;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cb226e44165438df4518876951c3aaece05b095492c9e8a4be589845eaf2ebf7afcde33e9c9fc69fbcfa8c2a76e34df1105444616761a37de65db914a7fd91d637808ecf1a3fb700ec428b4039759bb26c508e4e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h167a7a5e6bd4908c7ec98ea950ad20f0513d6165949cb038af8ac81cf8056c31264c4ef1dea9dc625b141da8ef9fc8a0165cbfdcd79ae181657b55982e6a35a48c28800f91c256b7cdce27a29e69a07d0d18c6473;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b71004479df653c46f231fa9b68ebc6f8353ec8d7dad1f191c7b2ec7e090cbcd933290009a83262fa65a9015d3c58f2fda0ef47ceb01154d8e238ecee8346a928db8556fbde63d2240bc48a203f2abc11a5675f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7eeda54e9e72a101c3be6d9b2ca57cae4d12401a404aa2a2b88035ec76840539e3d9c0540609e64e52261cc4ecffc3ac6f2789418db92451ee58894fd05c40e36eb6e3e45d01929145a1c47dd43617e649c496883;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ff34025b0771d3009774f447db476cb49755da60a33be225125ee2795431965a441175b0b07ee47c7502863b31c0ede2c345a578d69b5ef719dcf18dcad96000bc54668aa59d4e4c85b85b848b3e55e0e0cf31a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7613d6ea3ed8c4eb435c060792bf6de012f8b17871992e1d97f46428e29360192c5ec7973730c3287628a1ee142e9797b68ee4fb3da8f8fc40ce9aac78b880ab499898145602dfa274ded1fd9d855148e2dc9139;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4369285f34388f7d1f18f5b2063b0e41f3b7fbc84551535b7b51c56e32becfe2c1e7863a501c66860d2372bdd42d8b48b538359f2c83b0048cedafc01eb7f66cff142ba0f64fbdcd2100f89abe6aac2da7b3f9bd6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c6a2774575f5cfb070e409a1f9722b1f9265b7a5f216851ccd68870e656eba7350fdaf4af9dc992040ce4eccf6acf562fe888c1e698465575861d3c05943e26deba0f662790217e6bedb60f75ca125de0c056786;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2af756e4758fc94ca51b0d0b324d2ae1bdfda9c8d9a574b58fe4eb12deb342c4ce5e045460e614315da599f2520a1b7c5fb0be0793dc696ecf59a90596d59ff20b21408f3e3b1c7f549e31251f38480a7b9068c0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fa4f6802d2fe0357b5d7da7a8598b87a9c995bc2d3a86dfcf01b3d3c1917c27881e9b513dc75929ea4f9da3d69b3161b46475a7aebf6ad0143aa480d34fcec9f7b4121c322cd7e14bc3a1335ab1cad491204bc7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba98d4a6519af3d104c0dc592fbf1f0ea597fc23d05ae28b3dc636d9921c0287aaf9d6832672e96f1df094695309dc433b2755c1b5a81f4a5b5a9cd4940a0e7e6190778c1bc01a7d021643f3e36ee890dec69394f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60c81f4adda138def3865858c23dad6376ae6e12327b6be3a647e18b7c1f6b6201f5bfae4b3d9d94bd8248140092d6707e4d5d65d429c52b0982b0f1e9721c9205f6eaa0377d7d4267e09c548d9759d5cc6ba6848;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h639e439701f14b0e15211714b73e3e17f1af45b685c2598cc7921acd489ada0b814b24d8eaf4a700be32bc0921e7181f35eee0c957c9ae35589adeacf04892d785eaaaf08657c68a4d7c2f883dc7b14c34bdc0dbc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0be745a60f51c5a85a59a078e7eff0dc47dbe269bf41dc6b6074bc31971880a20497defaf8e1bd5f51fd057280180cff34e3542b6ad5422bc9624c7893559e8890e2a50e03a8e02c8015cdb216888e8f13069df0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbef3784979b6bf892caa61398b14d72512c27c4e5084a70043f345aaf1d385fbb4d400cc78c0ed11a97009abd3088e412885730e0042e855ce0472bedfc2a5c90f0269fa08bc3c3ec40da29b0a0c9d020c30bd7a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1f8c359c8fc2b702af4b8abc9de1316683b65c0e6ecf438359f7347ff497cd88bb085b06212a63bb72716ef396cd72039e4c667fcc71cfb9d13f19e6c0f95a0032aef2f333af2a1c3cc1ac40b38f1d882fb99637;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a2a2ed9b4aa26d88fcfe693cca2d5881dc69f57e17384cbebe1fab486d7c413716cd3d661713f0fec42f0783de004aab530eaef3f0c454ced820f51079a233b28843c9960e29f8c8de27efae292cc43530707df6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26ca14f7515a7d5b5b3b5fda5dda1d444d28045b32a1b9fe5d08f1d24900184ac9368485fcc3ac17e3a6d3e93fa568a5e1ab3c4074cc3f16b7234b14411884b81ea4d58b91b028f9ccc8c2804e6638b6f253547c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57edf8612e87b3f5bf2d9879897c6a2740f734ceba7f85bfddab258e93231df567d196e78cfa23ea1cedbeeb00307ad4d43721372ea3cd41e7cdbd04bea6aa8d35e74592a056dcc20ea511c0065ef59857dfc19fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42e03ff5cd2e4ff55520958d8d00c7b59cc8bbd7b365e2f8561afd5d58601b0c9bdb350146e0142db349291663074de6c4e2856b0426f9799dbf8826c524863bb801b3177c2f5b8d91fadd747bdeeef8d69c597ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2f1e00ee0178c0eabaf5dd593c399081527cddb7ec3c7acbe4a1892ee6b8f7afa293dbd352cc5504d586c2c3e94ffbbd5d4b01d48b6afcff06f2f37fd47ff40f7ff7a0f1ee2c014c27e9f4bde6192bedad62fc6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h659f5dd972269e5eaddddd19c8ddb518ef5363f6503ce4902e9a5b09340dd35822b60e93f727345562cccf09ef9df58c868da848e327affd5bdb0633877d0eb3d109b7457bf42140b07c67b2a46559ce31345081b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65df481c8301341625e88c4f339bf0a58d0d3e872efc0605744cede9e0b1c57339aaedc2ff9d99335015396459057fe9b2b9eb52b3b03cca9487bfc41cba72f4bbcfa15bbd673f698db42b68f50c78fe83d6ec548;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h732bc62b5e45b215b79526e891323eeab8e4c39c0188bcf9bfe781a4b65e69bfd1a8fb05f052df48b7035503ebf7efaff09271f5f3fc4bf36b65ec3128e42dc9554de477820b030e3c84c22785de984c9ad22affd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bb92568bf6a39136fbc6d04cf222c29dfffd596f720b4ce7194336b96f8fbbd06ab130845265f05071a12a2a97694495fa78d06b64efd04baf0d112835531e7d78d32c2eed4030eef4233428e2561951f7487fab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e7b1b79aad93f501441b4e0293facacda53512e12cc2131ab8dbfdd123f3800a3c81041c032c947f3d6c5133eb3954d2cbd5e1cb6243b4cbedf39d02f2655e3100cf120d918926639c6361f05f66aff4ed45d5b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdda66d5dafa717b4614106f58f4b91dcbd369468d42f9f5af8e4c3f6994ac69e1b47714d740a6237b77ef1f29c0683056d6d8fc621c166863fd4bd10af1f0b317cbb947e88309c5a58df3fda219a5ccc35c80da4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf7e2dd81159b122b1c9d80b98f92c06b8b3970326a891dd9f984c821019341a88a5e0b7056b2fa9dbe5ce424262511215af7f410b96c96fb071b5b28f861ac4269285c867cab36c53f6820ed6ff50b559ebaf609;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f42b4cf1e270c65f8a7a7de23440cce2ea8c0a017d6f2868e4a9f0b96d035eb7631c3a12c9492178908d5035d567819be3f6d7a453771d3ff4522a166620b3d6ed52243ebf7710e71e7b5c87e0aae3d66fe37bbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5784075e3710e41bdaf1a7bbcde7b112688c44aac6eaef1a88c9eabfff7b18d941c28525d86a5e321f3fa20114adddfea4eeb9e078edfa0f3b326a239a621b9a089d0cf1d144c8586857978d02128f6d3e0f0fa22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5908144760581199b319e3e42fb7e2a2371ff2e7599694555f03508e4613331b6106cba61c563fdacc7dc490777e1aa7cc4716cf70f6c4b58ca46cdcb08a03e3154b93c8a14e9f69d33d5b4b9657b405421242602;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19cedbe7ef65b6a379b2a791910802a8af5fcab2656543368fa955a77fd3d146a5b0f6ad82f139d3c859e7b6d7a9c9cfdb915d8ea2b2eacdccd7ac9d2c39baa8d75cb9265fa12cb6868958429527681f032c33fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82becca7ea39b5ca6b8cdafde819a13e6d23e73470a3b64a1b1a6ae28cebe3576c54bddf00372f57a116846b920e6b04a2bb2cbb3c82437e67ff9355692a2ab98b35224313a5f626eda18730d69533cb0057b96dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c2fed9fe40051b1477c06849c9465580bded93c67a55018d6b37d1c6ed89de8f795e5c34a0c83a863fef4b5ddef927f69cf842cf3d48b3add11c4130adcc7fbfde6937febca944652ae7eadb4f41cf58c2327634;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63fc0cbba6d2c9592a0a5ef39ad3ccb033dc35e29f5a36d4d30fcd9f834454c7ce975a2092fbfa7805964c92b1b1664e49b9691a68dac85247fd2c7cd9282afb788f054f673986e88df867cee40be7bcb443a67e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ed19f5cba67f4a64826da107d92505cf6bbe582868bc495c7a2819fb7ffe6e9428a5b49f7a525f09f724bae28ed37d2bb49be08eb9f951304b1817cf14252545488bb138b6e08bffec54343aa1ed55237bda3d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a007171e1332839a44fc90e2b5dfe06e32437f7b6c858269092bf1b3f45d216174b5cb08893cf0e81f93aa795774a2372ae39e67f50e0d7d818eec6472e0064a4683a90a84660a26ac0aab23348e51efa0847dbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46099a6cea5db5ab37dd6cff62d0db8d5b45d0246ea08a96a0f0b254df192612f6d2cb0f2fe91a5e3db518d5a82a5a858213ca25056d0356b7688b02b5175317c42146d4851e4ea5c78d6d9d37a7f9b7da6d3f17f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a2f9cafc0a0f7e335aa348b7ef89c30970bf3359bf76d20db69ef4203568c27939c813e01fabf45716cdbef49354dc2be45c8fc0d3610027833c5cf97da979ba46d420e235b42a900f6b97d2d28a9eadd6f43eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31d4905246087b9b09585cb1ffc1854fce2ce249426c7e5b16017bcf3f29782fa4961958c3270c356ce76471a806cca82de91b114a8ff9cafa37cc59e4ec0f77358ce8543e2deea5299e3acb6a365e3a0548c706f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb795f73bbf5299518c04bf07cf0e6bb743aa0b728befbdff9cb77b006d8a8fc83d44a0cdbe3983604765a9fb9d6d8830c0e559dc3c631b88779276747c70184f0eb1646c82cd1fe4af714d695d29c9e4611fc88c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4993e3c007978a33ea143179a54e1b0b21152cd8cf8ee24f3b6b9e029eac3596f2d6b5d3e61226368a7b40b407f0e1cbf366c4d6a890b1065a9d00bc5125ab6dcc8d2dcc2f24295263d610e1e25bac94b1e2a5351;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87b6ae673a3340b695bc48ddfc270985057a8dbdd3f7c941405cead3eb4bbdc7a549a08a049cb3834db083c80ca7a48174e9322743d2e546178c4af5176dc3b478c786e03e8beb431e4b3e47e5308ff0b0cf1b92d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e1068f750978cf3bf0a4d50273a01cf3b48eb5e522b8bb60d69c14c9db9fb21c0c5a262021e87453bf611b850bf6da1638b2972400114f750a4c1886498ff85d01d4cfa4331e44d6090123b33bab00af59322336;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc14499a7eb10648764ea98243d595b4b057053e067d1005ba3425459c04f80a4baa3ccb7b43205f41051ddcc68395bf6b9254e3ca59c2c2e2247625b4f4bcaed04dff4589f250d89a77bc995d0ed05adbcd3bc850;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ab91ac60cb9ac110b0207f49c8838bb7b6a3cc4f737c476753a861872220ed78291362a9f13a93f7260a8a86fb5bd573ea0189000910c75c9ebba6b9ee806f75f463f532f8ce264c05044368ee05b5f736ab7cf4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c6b4d789eefc3d1bef6c2e6087cecaab7004902fb4d24dbfcaf324e536cd851946cb2c893c413b05f1d7036297bfadda0e777a58c3f2871b17e90e697726e91a5acab43da6750c0f928024d7516222b3690e423f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50f48e5aa916a324470b325397553fbeef260f3a11a30f77a635518c83595d41820b4f00c1a7256b366273dabaacf95e4a51068ff901bc05f56028f15dc388d174a6f11613d476bc6f7d87ea7f48eb2d51a177f27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3fcbc5eeef5586d7a956200d7befc2403ba0e0b358aa12ce087db5a97ed8a518d0d0d72888eef65143d6dfd43252e06e2cc30518233d3943ec88c8c68e777fc8d15a3363bdbfa3fc8dbd1e356aa862e379a9c503;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7492921d82a19444d859fb364a07ae2f6f7eff3a024d3729ecff828ef9b016ffc15970894253bca456d2edaa74d6d71a4b285efe242480a96607755bb6c0fd01f5dc2e474d4b289503e811cbf9db66f07402eb5e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8928a51fba944c3c4bc7370ec7cb1564045c29765e09c4914953938ce28331dcf5b7041213af5fdc6d3d29945be552945e9475fbb2bf8527ba5cf34213ea7c51ead853dd59133872939a5892f4b367185e1268e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d3b9feee87bf01a16feb6e7ead6a2d1a1523f1bfcbcdc3a53e945cc72880ad7c0aa57e7b3b2087e3b754b51b543d039677948a6984298f3e1bb17711b2aede5ac26879bdb4292fc65982ea9f9941ead556b22539;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd031f672eae9b8d8ea2a69e9df9d9dd1ffd682a4eb0892cb000b71fc1cb13974d5346cf6d7388200c0774a7e0d7f63ce2986b364948a6c39dbe998fed9406c7eb75ac7a0d4dcc7b4dcc745e9289e20ef310e570e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd427d313e8031d37c018a7701b1823bfa419a6a5bf890eae288df2ec2063da8ac383fa98437449e54ab7dcfbac9aabe2eb5d04135cbaf3477638d609b8f5c0ab8bd2c81b9565d1431f2e17c4b070aaec9a907a0c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f3469b895ad7eed9d34fa56dfb05f8cba9a9066395337f4776488410f2e91becd775b3e15d91e7e1eb976aebf99a2c472db8cb96d7c85b95799b1514153ecc44fbbf6b322a1d1f7481127c309de39e8a758828c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dd34767d2af5de5ec8f2c548d7b43116e7383d368a7cdccde33ddf841261eae0fd072776ba62e74b4b6a1f6b959df3538e6c01272fc81ebfd7c8bcfbb88af6ee4c71b7d1b40037ff217d14406d97503879fa76b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c4d0bc680eb77c3c67dd56a9e52b6255a3b4f6e30f107ea11aab0acfd8aa3103352cfdca0bb806200b539863ac42fa5cd115804931c33c48784a1a98c5441f05cbf0119c367a807c5862129cef57565b20411fb4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36b7c1030c62195e9c4150ae3ef57d8d2e6a48177d0d3b5d7fc04dffc46207e6174b5fbe33d7ad082bee78bbbcb9f758848f55e86f44760c22b4efe83565b067ce89b720cd1eb748422213039a23c3cde09238e81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc091f15b56d8e98edbed0cc333ac618b36a4cd2811a5c2e08cbda5a36e7565ef09405905dbf2f60c7b770f00db3fee3a109a52d59b00ab312e25acfea3b6745bb86ec4c7b3b7c9dd7ca58cc3f455d8886f3ada67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbb3dbf8529fbc222d0eb6a5d85641178dde927b997fe8f147ff4f640c2781e7f52276beff2ac475b44c7062ae2aa285c5e990aa5b8ec03fac82c9db2393318e6fbae1ca9dd0dcc89129b5f7ebc12fc0a8a9f62f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha130cb26bdb05e4add569c4085344de4e649d74245e4cbb7630fe717d398298517514ad02b47485bd55dc624616f20c20197385d55061f5eb162798a64522985d99b8a0cd0a6640cfecaf78223c29a78cc2dad3ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c26da7ff3a723c643d9f90f85c393b6ddb1468f9b3b8262fa90d30c94afc2aff9982fdcd57a86124fa22b72522997599b6213a9af059ce98d0630c15646dc0374e9601bbc0e6fbea48f0dc149b01575d361a7e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7688ca08d11793f53786698459a8c796873c1c7ccf5730feaf57efb8455fa78a1c49beaecc60064927d976efeb1f65f273c6bdfa34d4718add5a8b38b9bfeb71370f02ef752e016791da19199a0d62e3f4e16e7fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c2002796a453d07fe58f37a9798fa98d9d8a587c57284b39c1d62387f0f6860c9aff5e8cb844481d2b4257442378b0a95655aec1666acbe96b3691196bae9e7dd3fd0db68fc65875c5853c0b78534ff1c68f9798;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h127e302a19d83051e847460c5cf0fa16ee846402ed6b7cc9517e7d6b3636e7b40da143056784757728565264b80b6896ee78981195f5763878b291cb6c77031d9b4626ad37fc166386fe924db595d5112270c7ea6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5f9e6f4eafcfb518c26b70acda20260afa6f35e538f765f7ffac9e45380eba43016bb855e3d3e851183edd969c4f8f42c2a798e312d42dc519d560174ad2ebc38691e962d5c0c7358c7ba1911ecae70c7f3ecf7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c06c4721ceed86185397294800306e6e22f2d6a670323229824b87fbd6d4ea370fb0a994b53b0d065ef96af839b27c59940f0337a97bd61bb451ff2d62858a1d3471c0ff01ec9c337fdb748fec107565dc48b2fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfa8a9444f9e681cfef96c749b55596db5ca6674303cec752244ee4e22a608dadfc05c3d3277f62b71807d2202c2d710413b745976982065439b2a262d6887f034f4bd9a339a8020f738ed0ba784fb84cfb5c8fac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haae82bace1a20a8b7edab8efd5002b6d11f523f9df50ecb69cabca4054c80ab9e220422e9dbac24c37229ef4f41285af7b66f09166a7c6edd6e09e690b77bb3763ee4bf39a8c1e7ea616c5af9281b61a10e58af6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe7cad8d8fca4a47a2e9894bfa5c4b945ee1b3759e826f0f758a1ae53a7e3dfc64e85bf0b8e09c6b9c7b4147ff40eaf171403e51b609596152c4dce0b30d97ad415588d1e0822f63f497d4fde7a15a3d5336b4029;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffa9eef29e24c705c043c89d68d00d929e017c934591e15d7c6b249578befd16f179c2c35fc30663e1cbfecbd423aef8f49a923253480e911d7e8ea3f0b43177310cf8501ea6b67eda27a3a1296c1d61ed967b5ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha29ead1a0bf2ef05c5d8668bb5ce078b499b9f3dca9e2c2c883a07c38b55a7c3f6c6013e027da1769e7f2e65186b994af232fe111f86ec432b8e634631a0db1f4275d9762b4f43d594d2ef6844f83d8823dedb367;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heee38b6f69793aac20a57b6bc12f68c6f1fc40bab2a4f855724f855982b8328b67c6aa4f3c65014b6fd685f8c0ec993a227664696cb274bb5c82600db16a787f64d57277a225d9fc2358bc8705187994bf2d27e5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48c4e68c3314824606f633e220488ab2c2e55225bbdefae1ab62d82843f32a2513bc3d2cb2b351b2ba6593425bc6795644990efa7a64ed49e6aa5f4c7f1fc99a0663d491a9aedbe4929ca8795bc3c4751ac6188f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he00e73e59d90a70bbf106fd808e2d2bd8b98c73dc5542bd6a6639f2a1f1902747597a71ac37506387f0b1da663664f0a02d17e49a4f3cc9e44c37f0126c811b325f62761c0e83ee2caa782cd97a47414f5dd2ff84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9358545560c5e9bba55d1720cbaeb6b3368ba63b743f09aee43ea7159c3c01253c77dc1276b8a2062edda2f3c7d60944ec0a20de459cae2bf4e31b46b9cdc77977426d1fe352db7f37ebb00cd08612b1147fcdc70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5bcf8c74ace1b0146dbdb62cc27cdac4b7257dc54401c6678b390a536377a68a27e156aed6d4ae00b870c7521081868eb5d99ddacd0efe5f39e519e79f0cc38a5a7b82bf34e0f7cd179c6937f18a8f71f6ec70ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69c277d19488e20c970a3e4ce1eb0afa6d95db97c8fbf6f4d583c8478f18b6c7a01dc729f02069009dd735518a0b66b44acb8ac04a4e2b7cb3aa10c430ba6bded1312e8f3a3d50f40f4b2f044177e88537e37083a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0205491467de1d06849ce250c827fb2ea6e43f63d8842cf6ae6f8dfcfa227d3fb844b5cef35f324b8af762303e4ef2de7199f0f43942ec4ec58508c96c43cf082ea0d886a89efc94f37076365e79251996426ce5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d373676c5ff75a2dcb3bde2bb7a7a8d2dc46788288ac35b8d732cf273a3f42161a1a69c6a199cab756f7ec5d3a6788886e36c6e24320678ce4ec1a13ff75850c607bd94df378dfd9d7f984ef1f0cecafba15d3a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfb77df3851b836c546a8252f854ea62d96a52d80240c136ca361f82d18fed7da5a7624f53984477f14151d0a1558344aae47f75909a0175974e50d7f9d2ff2c90d60b60b9833498bfa7ff580e54e2b0c812e5a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9cd04607faa33136869d2cbad6edb292624bfb8c3891b71e5a7af96ba1a13f0ef93f0be4d70683850b0e8d6c105bf7870432a54c1f21b19163c6f99de1e14ceafda9146b86bdb49042ea4110c261fb6db121b5c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8ed07981bfb7df706c85f686353276705f7d52b35276fa5f77622f51c1f283d2c1ba8c037154164b16449d8300cff35a770cf19b871a7505730405d9c9195721cca885459163ab5a8cc063dca8823579f39898aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dce16ab2b1b3d202545d0a97e6e5d9ae09847cb6db4e1a33e9410d9848c4305c6880ffe545dce37f5d3691b81e8d39feb0cd420b41583a4adfb5c5df2f8bdacbba34f879d0a4f0eae24abff1285b1a6271b6b246;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h660f4dd82240247432cae8dacb2b782b8154c2db0585ce1602537251541f856618d9fb074399e177d0e17b9e4ad8fa290d6f424ba85c1debbe6a8ba7080e64eaeddcb946788fa56b93455f6e4993ad120c7ba646c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2512d656e3069ef72663e8aaae9bba3d8951ad02923410d735ebae73d23f373f40f35f146a756873594b166bffaf162afb7ce9020ed7340ed300c5609f866da515ea962a9140a0a583c1a7db1ada15ca30afd2516;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h316cb633568feab5bfe82dd9bf5d2e98435cfdebdeaafa91be3ddc4cc9b24a76bb6468e82394c1cb0ff15c47714f063337606d2998e6dbc5c9beb2626c3a655f8ab472eca1a52da3f493392dacaf42e72d8c8a562;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h165ceab9663dd332600efc3d0949775d003ce19c594ca1afe146d240d27e115c57ae4df7f56c1709f9b7de6283a9a455ff13efeaf1d94e95976a4a1ace6c31d001a26c42185fa01f85a7ba0d5c157a2ab2d3b983c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf599454d52f33d466ef3b2deb363334ffc338730a728c78e07e575ca8333251e2ccaa4d522023cb5872e8f7958853c44407ffa9fb4fd01f0fcc9fce25b80193a6d23a5370b29a19e2b77c20cd98917a4d87bf6376;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7d0a725c2644e8cd10bb09eec716ab4734e28e7280721f213f0257475722798d4188ec79fe17f21bb7d9ac29a6c2b5f43970b400885dae605859848f7664dc1e71eac4c87fae3f37624b3e34a2833ecacba35724;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf6f4c535a22aa95b078ba584b98767cfef182d96e86af9a964d1347a5d3798c94941ee82416d1951393b33a5325e5fee471ebc7b55c553c88394aae1444203a2ce20979b7a94a0ab8d68c8a6fa896af449311b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf558397907278e0216e986f08e7a7cd0d81885b49c07951a2085d66bae9f34dd436fb2c1ee1dfeb3f64c610270e70e6638a393ede9d93f796a308cb84d5ae9bf6a15e5f2f3eca117ae1ab453662c5ec58c9250e6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a09414931fd07fb6c7fcadc8ef4e77e8af760e4ef5a19dcf06e08a8a092fcf5bdf5fe47ad92e5cd4a66579e89ff25fa4dff534ec923e508f4c2cccd039b1ad497d8e527289f058850c1206d1c4dd244426d0682b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef68d2da09f17e28415efe4ed8ccca16532c1f4759623c4325e5b28c1c0f80c6c1ba6268b71817371b9d1bfd47e04dd3f8e882c1a4b3b559015adb79a8cc333fa5f48815e3b5ce99a91213077edc4b0065ab1ea54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2721da0b762c4713a0c3755c84a7ef5588fba587f9de6a8efe159c4774d1b39ab63df1538fe73dbcc01b0ecbfd663ee72d5c35111af6628c5a20ff87f60cfc12ed290383fdb9fc43b051e16d42bf8124f7130baa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1761219ff5090dc425f50d42c9e0b019df7529d3f0c57b40243ff31e5441031c5b0ba9bffd99a370b1ec55061a8fc83e7c8a68465f34a5984e89c5d768d2b0153a04cb0ff95e40fddff73a60ada861fa5a591c81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2cee6a99a4d5f87c4e6db20c08b3bfe93c56ba1de284453315a4638902b5c3de64a34dfa02e92b45a57942972d4baa94c52d7fe40a2ec3d43f25e2eee9d92b7f084246c35faa18a5efe7b4f35dfc168a10f2cb3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb7c9a8363e420981475fff985ff3b18d545ed52c32b9487b50b84cc556f1e1b41a13f2388b68a86707859ee459f40d1eb50a48dacb2f8aefaae5c0c0fb92a4833e976da6a361b39250de9afb5c86174152711b24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94753f387e2c3dbf2309e29a92afd27b1c0064c022b42dd03db122ceb39cae0ac2861b904602d58c164190458b1ae15cddbd21a80e91f1580a694052d3f5cf4b4cf253f4b80fca316f16f0dd05309c3144846ac06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h543cb591aa306a80cabf708714397ac24e94232c83039b773f2106d44e0e0a5af8cd30490b5c97e2e52176b612775c31755dc6541698215dc9742daa9de9ab1e87bcac066fc8e8720b1715c4a9c583977358be5e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2cebf850a4b1875dd7a43c1bcfb3ec8f1136400c799d33d16be98c6c7f52ede80b6e6cf6293bfdddf69456c82d023f5fc40fa2d6ec962232d11e3c3afb978756578e43ffc1f6e6f1747440a1c97c02fc361da7bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33e101b1d6d7fcc72e83c3c835f2fd5a510b354c4cc944fdbe6c9645a7f755e87deda4f1d4146be4f42bb2d7ec576b52133ca1e2f9426a979701aaa798f040043f5c2cb8634b015836eaad01a095806013680eee2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b774b4c24bc0d433bfda8afafc27b62fbac13f3a073cc8733d901aa3d14bf6be332a9a32856c6f11963287994dc37551c83b13a19acc38e219d92c392700bbeb2b9fc24b1f10f7ce634e9138127741520298ac2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64e1c39bf9e940d1b6417dfb9896f1584a6b5bf4b5385e1480cdeab5c89dbd15960aec56f02009891d50ccecc394877e3bf9dbe1b0a14620b0f89b74de26dc25df3ce688ea69aec47ccd04d81c2dd2538ab651422;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb82ac06218a1cb6f14fc8b2083d7b44c50dd974f21a778be3de56c86abadb6ada44744226e647b01fed7ea26e9567dbd3b4b1d36941a27e41f144c11015a1da5fbbc5fada356b2dff6a03d193523649ea560ab1fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c76ee441aa72c87a815d46307533598025fad16037eee6f6acaa4ff09508eb27a71caa121f4c8dd601d67eac9b54032096263262cae65237231e2f3645103575210de93c4759841252e3e5fc0a3e47ed41576043;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c76c7b03a0b41cdc9ffa08a1b867e1ef10aceb6c495aa590735b5cb2deac950f93eb7b4bd511d0ff93a520e65fe0861ac142464b163b6da02acd9727167f79e6033e5a9a32da869775f1ae9afceca96c240de116;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51092f98337c222763b92db9bc6eacdb8ec67de7e678efe0eeb56e3332b3ece4775b5ea51b1787862d4f4b5cac4f56292be740d045d78ed20117d2918e440aaa62f9bcce521e1a709d14c3fc85c248a55c24c4f9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6b420d3e0d98890bec9a464cb45bd5f228b7b2d762bc7fc67d663294e2b89ac05680c1072e219f9afdcbb4518e1ca54e561a0a7f51056bebdb55bf05ca655b337933e68947756caaa5e0855575c948bddad71c43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8550f235cabac4a842187e545e5a8199eb0d281d0899755caaa64553955d69587ffc537e299a1ea4bf7d6671f31dc9a549c42ab4d6e71000f6da4f5bad094aab92a5fb7789c6bf00c6b6b4356ea437803e9cbcf2f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8c6ef0d117fe1f0366aed5894ba285bfb34ba70b8cd7d64a3d597215ff3cf4ca16fa0ab1c82d40e10125093844cbd76d2b681c9f54411eed4bc213f3b936e9e0e5ac9999468f808d7ccb985137b932bd60d2441a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75296d55c2990ca1fc365fc8f5fcd8533e96e541d2b59d41a34a7aee0401c5c12cbf01d9e3028c21dd0466f6a3ca7455b298e8aed83537d7fbeb5ff8260b6c40a2370bb1c1817d02438e5519c2d7a26458bcd6900;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ce1020f72c6ca62145c1543f7e16b7f72ca25627729cd3f5bda6cab56be26a55d959556771e871ded677dc3624a6927ff8e42704ff8d148b9d00dcb19e984ba08463396164f98f3e86b7c1f6e4df313d2734c390;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd51f373cd00bdf167f8dd9e9e1617b8ba9c6ea39545b5a0ebe57411e3f846f7b1e1deba5dc728734768926355ec5c71c806b9ee6c36202a2fef93711ac9954b5a854af3b6df7b9e6987a7b925b8cf0be1704dd5e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8d9b5163e731401de0a5b1063ddc1fbae5a4898fa8ad90b4d952b5d547aa99b2f025577b7aba3a79cd67493839f9ed643dfe85fe751e13ea67244495e6441ef26029904437f3212c592463a7a08cda77aaf9b133;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19c070f8b9f77647e13e7ae27dff6d8bab825b0df8e08b0824b198bf402800863cc0e5f57e184eb2efad7b8fd31d60e1509766d8c768c438e1b530f182a5fa907b6ba17ceb1f9604aeba1aba404730d5f43c60479;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7c4531ceb7da5a6dd2eae8158722e34f32b60d080f1749cd02173a2a7b23aa818e9ba4b1dc1f7748ef441633f3e8a04a5818643df4dd9fa8bed4aa152435c5747b2a8c8928a241c67938771641ed7f9a8bcd6744;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e6f3b040d4edb1164bd0dd811c3e72c5eef89f611829447327eeb960e872147d0f346345ab4e290c2df1277d275530a927b8d486461a89166165e327a07b57a46db7458d1db1bdbd9b7b4f0d25109f2a5cd09738;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a49ddd86a3063633a500c34615f9bfa3f26fbc5053f7385ba340ef746937f1f19f196aeb52cd1bca21ac5ff962a575c87dc69de579b90a0d548b4dbcf035a9d098325981234e22108f217f7b521476b9385228ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41e2612c5af6113062a7f970677ab121830984715a2902f9faa0c9d71981f1b4aa1fcd90b7b47dad9462f768f12411bbc20d3f6e1b9a502b8376699feb96f2268ff5378998f522a2fb844c274cb63610a7c46990c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha34d190df4fb75f78a4f44b4c8502cc293ef33e4f92b424b2d9d648871e84f98accd1440729b553a9b721fb2d6b791e30f3695203463eb73850481bbfe54e2ffa36d65b5b440bb7a356cec7ce2df1568e0e64a165;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fb2cdc317aa0296002bae61b77472b110b7e015190d98dcfd334ff330031df38ffd365191c3ccb26e312e1615bf81e31e854a99183cfd7170460bf19a2afbd4366e0e629d4bc15b8e6785a853a243c892da583f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc59a049633552011acaf28815dc03e1d3af454875110c3065442c91f2e233afd87427527d07635469b97514cd05fe789c1d6e46f41e6c10e08a732f6a5dcd82581aae872065610bc13be68a6d81dca2bd7457ba9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70fc7ae1e6dbcbd058f54efa309ef43529a193c49ad24fef2eba4c0788798e9a68f99f2d27b4e5465b027250d020132c896fcaa29fca4ac0e7c0d685fa4ae554adf7b44f62f32462ab3ed0f51f1f6142b6674ef5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cfbaa1527797e23510583f8cdf10fbd303667c9b6a9778a50407d1afeef54de47d88d4b0d1be4c9422de827fbadea310dc535743c954fb04640fa8869edaf074231324f21de4689b6d1bfb6d00230745937f716;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h239bd1e19ac5a7975dea7c4b0ca8886e81c1a5a749c596cc09d6de55c3693ec1b64cae76ae593f5a7a686e59bd53e855b5b992352e63a7ca1a66907312dd0053cf98db3396921ece844b6cc75f89bf966946cd455;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb31b39b8417a15ff518d86bbc09a7cddd5e978bc62406dde1efe4c2ef0aa8a2c61db746312833fa55a0435d243a71bc8267ebad885e7f6a8e3b032640036c3764da7f5f12a34c71ff2c58fda58d81e5a95fbfc045;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4848c9052e542eafff1bdceb0cba9b6d1dc6853ad4f21753aed46b73cde4636babf00a0b06ef73b8450df3acc41bf851ae76d746bfd0977870ef12a8b5dbc920be7d126a73437578a3843a6e4b5e270c8a89d59d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e781b8b2f9ea075d7e69cedfdccd462a7c65470342690dbe5fe87ae0c6126dfb95de68bab206ace62aa730a9baa30093b662051914ee45bc2d2b6b4d983e3f25ab60b0eafbefc72bfc60ad1bde5cd7b30a00debb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21526ce387924ae0dca9f4f4d3091199d9727b6720064f611a3f28e07b8aa3c6559f61eed8b31379244909ea54cd8459beb537eaf5d57fd378025b7d5b5aa5c0390e8fa188b2f896ba456562e9245f068c71740fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62c58714e6b4564b781affed856b464f91d4ad8f755d1e764b4865e2047c2bb21514df2527f0c8bb05a97f4ae531453910aadec1b4f36782aa64e7d7700cba3d42227a76d429cbb8a1b57323526e661e4e7c3f44e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h157b42d5fe638b70480d4fed9a96ec56f792162a65a9dc69f166c1f3213a1a5a7477bb9cfc642f3d2f001608d9621a4ebb896d4f20262f8cf8affe126ac7b1179e38bb71838351152d7a99d148cb4fc778edc1d1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb406bbae6b50f214a8e532c58bd2733e753601a0075c067092489c2e70561916852fdddda70277d645e9341d9ab55cbde93163c520f78f46857892122ece55ec198d44fd16db4d72d855c26cdd7ffac70bd91911e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3abfef008e0affc16dde962bef8fa485491f3e9e036708a2864ed0e9f9bdbb2b991b9d07a31553bcd0304f4d37263e691b3f407228283b5ecaf5059b6f4abf344132010b1b6e17454a833785e951c72b4f8dc455f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0e949f3a80a84ba43f873ec3af5eb0541f6c0771b1dba682537f6749248af05869135d798c89f72ffe15dd36055b3c9e5d05cc79da37963e130c8cc3c213ea7050b251ad88d079fd5ce69d595767049a88e28508;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fa16a10edd298dbb3dea561c9c0515a23e29e47b2f36b0fad325348997b6f1a215a2e19a041ff2c26c12c00d2390310c71cc7b801c9a84c9f92c7c85d98e7a4c0ccb6a8d2de08abd80ab64e0c53fc3d711788af3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha75c81d54348200ab93953b35760651c710210c4fad28269f27d604b8c2ec1d8cecae073c1d39ac690447413d22275922a680f7512eaf7fe573a763aad684ac83ef264c408be1708be10b240183d9eb0707e3f6f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61cc249e7e782aa8f67214667c26ed3a13c09a2f36968892963bd5d6397dc1b2669d464377bbcdd3b4246e091c1b2b3559b3ef866d4b672e10ac6afc6379cba621086c11e4b09b7954d1134a4d2d901b6ae53ddb1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55cb4eadd3055cfe86d7e3c13a8fc813f2e5d77d58d87145063059d8aa661a75cb34b43ce15608797c6b616532c68cb756972fe49b26b6dfe6b4468d4243af1b1ecc8125920b7178ec172e23aa477ec9fd3e3ff4a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h502b78692b2a5a12fb8e63e98338b9f1f055e27cf9d8b0444b407408d6c19a3216888a10584dac2b7f030de22c9aef9cf9814593ac341fd1ac6495c9e8998554b71448ee313930c21574ff215b3dbe7741b1522b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h205e9e1bb8af0269f65d57f7fd40002e58856147900fe614543401569da128f0878579616a1c2ec50bd47bb2e2b799c76b3e32281e802cc14b64e7553a99cb1f7d88061012be8cb10c37724de59d35337bac18cf3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f8309cd8a7ed13f531c98d64c7fb2fb4e48c146414d2354ab876363f1e9c98b73cb3a24a3fa3dfae6999dbd4d434ab279d080f29f13d2e27b74166e64f113d0edcb66f54a1019efe0a8c170067dc5dbf8702db6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h857f2d4624ae131b8f5f199f10cdd4cbc4b867414c48ec5898472ea8ff040403f6e9da1e4ace51d1db6d4c96333bcc0ee0a4c76bb73a6c6ff6caf8a41edcf67bcde96690844c861206b2f5327075ae46b4ffae537;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ae1a06a89c802ec453d97b98e7008189103d3ceb89a5e8c033a7bfefb80dc7fe26de2f6e9658a130fae7c64f615156750e599acdbd359bb5dcd1067c5068f8e88a079c2875bc257301ba6695ff66318fb32fda81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d79f4a6a25b3164a0ce7581905c4ba499e48cf2e750ca4886134908b99667990b1612b6d431e7202b65618793ece370198468d1462f3e442086eff1bfcbbd32b8b84d8310c883016b03885228990985969630b10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeecb30e5ff58fc7f6f9ad306b6bfaa7df5a073b2667390f3e0f757ac9d4a9ffc3bca4b36dcdd9bad1aa5b3df8cff97a1170d73d9e929be793f90af85527095b1c086bc66fafd5289c8f3c55f89749f2348b2be7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h194ae71ca43d93862e9529932665281314534d16aecdc226f1e9e7cf6836d23e95a74e01a8dbd03a977e65cef9a17b110626bad6e36ebcea04a6479c8096a0bca8c50923bcd783e3bcc3ae6c3fc1faf1c47539298;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b9feb5fa0ef8b4f4a5b30018b79c23a757aaf883ad110a14a612814c0533b96ff62d18707c2f2a7020d3765a5a2c4412aa8f159caa12dac3606aaafb02094da4411cea5f619b7018b4987e4a8ddd943a39c482c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29f49c58739a63565be1cc12b8e386f982479888c68fe891795a9c550c2629c6cc181290a676a40f18e40479e8f39f587c75c730d99236495dab853477ab1382d02df9ef0c80ca7df85f24482d0bf455eadca85dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e5fd406af33b852238c6d3c4dceb594b6417d8fd12c8d138db8d4db439c63100820b22b5aef21dc35df87883724d17716add2f23f705caa8ee1e43306ef716019eec5287ea356f6261acc5b810fb62d292312e45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h810e247c29f4169df215562b8d79ac6f4b8e0343ea6a42d22d8db39405c63635dc5e6f9e9560bde29db3fd99e61e1296fa8f597876340f31b25ff4cb655f7cbc2f2aa69cc24e54468d7e8c13b9b11439115832465;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa4461adb3914a4857d1e304f5725ac5ed14ea43ff936de486165218f451840e2f1b3e0ecc64ff9805575d489d621214741d146fde70f9fe7b32d1560a7936a66842e0398f73b82299f72326a39a01c5108ccbd32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb5915354070a76c7d71c644c422af60989ecf8cba3eec3b1a5653ae5f4b17c28ffa10d8066ff128d8149ba46c2938466034e1ed941059f35e3c352c6c4fba3570ad7da24b099a8a3a7de99f2cd9504b88716bfc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4af611fee4c9ead7b8f1a42ee16025861eafc8f557e8389c8189cd37d5ef4a8be59e6a754af02947a1eb1bb906fc02cae626db0b0ea5510cdc9a6f2d510910e643e106b1462f1bef671217b420ce904d8c1406069;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9646f0b0525c025e82af11954499c9e3743973b61a65cc7d740f7a83b39105d293d2a573ad25fa1aece1be5d5d45115d4e60c78ccc01a64d52b569112a7c9d5ed11b0e91e72227365255ba2deca041b01d3aa3ac9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h750d9d1d17c1e1033d225006823ba309fc3ead7a51dc396f668e3dac98d0a05c8efc5c41c7056b13b0a6f8271f170ae3ec8f8b24d9d216bf8cfcc3e674018010f116433540ad31375ce41330fe968a89952986cfa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fafc34d01242776186e1cc40021afcd24e25cdd46bfd606c5a16117a4001a5e3068e97c9cb1decc30813c5500ab3de394eac9799d2229089f4604b57c18809f8490199d209ac6d3c46e75f976d0cef2ddaba77f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h776bcda351c7c88098d4d04fa39029a9309cf16f605f333acd3d82c046a1299a15716344183cd0f680d11b5f6f8d16d99ed011c3f1add176b092ef6f78e29d8e6e08301422456d8ae43152ee45be8fea92de385c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c80de366da82da2161cb8253c0854536bf833ce5363b498376d6d07e0d73382d3f35ffb67eae035b42a3f54cee0dd626b35f285e2cc0e47aa6323a5a8880262823195eac17da3c287311ac2d4e58fd48258af2eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6474b9471bf7c4693faa5794b0ecb3f3355361ea4b6fa45de148aceef1b5e0d54369d72dd9ff27dfe1528133417eac657412b4e67c17bcc61ea991a1938d811db1a794e4450fe916081991d071031ae524bc7b9ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ced94c7468621e63ba229f721d62b5ecb9403961a73a834f640784667c08046fea9ba64424626bf0b7ad407025a785fd4b867827bf4739e174bba0cdb57ca83bbfc78873f45b82fa2c4d3aae91fcedbaf01aea64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54661c3c3a2bf197fd40aab189ad500e81e52b8faf0604e34e05ee80d87e6b8144ad839e5d443ae58d65e58a02b1c7aeedfbf0fca74bbdae2b4e89d7918dc953d1a988e45be51a02dd486accee20bb6037044b073;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc149d02745fc4dfd7cee48bc5cbe61d5482d5ae6dc5bac91b7dcb9d3afbf7cf64e21cb63fb5e2eb3827ad377df9140e055b52e3aff7d030ca37dd67952ca5c24cf49dec7f1be42eebc8e9c822189def8c6d4f4e7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha89d86b6b5e3a789cdbde79d4beac53808d5312b539b26f00531b1d73a2606660c004b78f5943449a3d4a5aab33b03e97b5ae2a4182c6b0a86bf025f95a631b441c5fea97c2783481acf95397dfd02a24ac84357e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf477c03bf076d622de326e1c6099294e6c6aa8dd236d259328db288d73d08129c076c94150a9cae8b534fa6a1949ed36ae98a8b20e97dc90c5dac2829c1e4173bb1e13d36971521673ce505107d852a52ebcaeddb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3df35706cb786d2cfe368d15e74e7c59cb038a25c1a7b7f7a3f4c7b0718264a6f572b8c11ce8347de08a5d2b42f7e79dd429a8b7d6a061af8348621e4b4a6ada260751542be2c643b9ec1fbab22e9fdeed58c849;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2b5e1858443aaf5c2503ea544b6ffc04e7b9b48cda0c69b2b149cebb62308f22a5f058e95d1cec97bcbaa73611fd22f9e319a4e4ec8bb3cb2af76546fe17aee59f15dc0666d23dcdfb214faeb2563c623f6ffd32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f1b2b337980b76e4cf3de9987a3c3e0a95216897993605dddcffc00fe7d92b617b8697c38c8165cc0d511c06e85fdef781f8f8aaf42f3dc1ffe5309cb7fca2d997c347ae139b36cacfec28afd16187b5b3525c7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd85aec75ff57761b8415664facf5eb2e83c1892cbce9565db8e06433339b32bf97dd3c2383acd8e270b94b4b85b53e9f7e8bf267ae4fdf456af7f42d53320355f3c15bac1b982f6c0dc2dc68e463bbc88b59495d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4458a8c8e77539e49feb90bfcd6d934abe9cf56d5335e9629b37b0c833a5a3426da6f2c190a7d7a72e72b7bfc82529d5e34086a3008a9f5d895c0b343aa17313f4f4ba4217bf3f7ffc4abdb3444e2e39e0330c4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31b7ae5b810d93959bb59b8624e087a4ed70ab4aa35c54872cb951481bc6ed040a69622e85b8f20023570eafc890623edefd61d9e5a2774f5a57372e125dc1180eed6f5e17818326ce5689ac692a9a5a14667c092;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c9adadb511365d5258a58cadc2533e1d37b7fbbd5c15dc3a42177d87a3e2a15c3db9c45d7989eb33e96f9569a114b5752b3f939423c076bf8b079d66a5322d94aadafe65c95277db59d598824533a67c8ba4139b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23bd22ab6b021f4a892ef17ee8d6d464a6285237e37ef3d626d0eaa991c49a606d0116bb6bd6d78706f1cee1d39d10be515c45e2ee407e8fe8fe871f3497bec12dc53191f900759883854627f4df32bbfa54569fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb849a7e53a4b440ddbe7058847771f195312b26c59c7ad872ee69a37fc4c3ad9c8e94ad2c78fdb311391be5f4f227efbab2de1e31a34fe7641feb69dc3afb114f625c4529ecb440f87d07f6672a48751d3f7911a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha972b9f90361130bd13ac1f8b36a9fcb58dfddf0c59c0b64d08e266d2cb5af4f4539b5aa7c113bbb4ac9a302342be55c3e649ad7f62a4ac25825035dec5d1ed886586e2c746ca09e2e682f99ed1a040a1c3f8e0d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28b0023e371f0e72ce5fff65aaf4f9fb15eaad4278d3e2a51b398e767006832930098521765076876b6b7469fe61bc90d3ad10d4858d692ac57efb7fd213c8db93cdb68d48cff488f86775b4e990bb7caee9d70d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea7b9e13ff609096c51bbe52ca6b566bc06530c25db896bc02ba8900a5454eaada10a4bfcd821a4af47bb7cee161e90e1d67864018ba4541cd04f66ee52578e52bad7e9925825a326f4cc524668b449ca323cafd1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4c79b1f644105cadb06a2a8c2254853639e025619a47a7b7956467ffe4efafbea5737ca79433d6e755c26804d9dd96b4fcf3debbe250e6ab117dd366265f0ff599b0935fe6ba4bc5c7350a4ad2662963009d71c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35eabfc543131ef070100ff8bbde29c13a40345c24d2d77aa075d3ae0e6e920b97760911fe6ed6bf96939977eb95450c3a37568024fc1e2aec7f0221f4063240f50c9cd7491d6b3ed6dac7424a2f4eef0cc18e630;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88eff5cce802c4e522c75f2dafbcd44817112f9bcb336995c869dad1383ae612a3db462e668219104f64eaf060af4a96106061153a36ca5dc169bc6cdc6b3aaa0d06f91907808645d9bf7743c6847a7eb95f2d1d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3432df1f75b910e00a2cc27425e29a6376b15f23c1352d091eed7a7fc4009c6690bbf82d54d5727ff92d3d6a507866bc4fc91cf12f2eb49c6b297026a6a3db007c92f239e32337139e8efbce4db20a9a4b4e7d4b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ebeca3850c2eec2698762bed6dbcbc1e1947a2df2a82c8e0c868ec5f76a74e1779f08a16b94056f2e024e4c8bb6b90df55a6c2c1d2d784029a21a41e7d2741b7563a6aa21085c62a01fe2346bc574f0e68ed71d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3fbc32063a3d77d748c7bd9ee900408f61794be45ab285c0e2b22978401fc13ffe627676fddab9a2110c026de56a29512ac3e222ff4bbb34d520a3d3b596d6d90e7273c86c4232b9848a7f3198230ddf9239d92d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5de04d8c896c7796b455ed645f572cbac6853219196f296ba276425b76f3315f9bf53c79f2cf36be718a4ef000f63e9536e43ac0ff3b7780a8b2af3f6512136183ccf42b44e38e63d774a54b8e080679e99e7b765;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h941c5428af1ed72f3ec6cfcbe40aec1acbeb301e5b9d29c8f4a6ec52691d011a50b38db1e17c420e59630279b5bde555f84bc306a5c7c72f86fbacbeb26300b5350bb9d1e47c83635957289cfef0a4db356fa8dbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h120e5140c94216144f8e6cbbbbe57198da787e72dde9f412f1750138f7f0ef6705611ced2252e91974744e2bf0255a59e2e1bfd0bcb23cf45faf6c6ad604f0fcbd2977bb23a445bb8c66076bb76072ca673731a63;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc18ad6c3e6ab25b79e1ff948c422457eed7d40a831c83caca698aca9c51bb0e0976ede9b3fe0b44c169bc3a9b3237591562d88d6d4b243a1f1a80a980309b3af2428bcc161826e512f1935b1195afd0f4b896b325;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h610c011b93d9dbecb018a50af6466d206e189c62f741ab59dff0af514a25c4e2d718e7eda831e197cc51372fe33cacda4356ca0aba79084ca417fbd5c5dbe43c9a1476f56041d91d6513e59e4f1cd0da6b8b4aa35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d5ddd3cc64fa7a63403af181332c864335d9395976eb77d9ca11e3e900304cb33afe200ec24214753238f85b4f072de5b02f3b4eaa6a123b74575f67122ea1ad009500262514e59a9b125f1d7f09de12e47b9c1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h700b15f4202b2c6c8d9f95148d83be0595b8b844f9ff50880d1209a757826843932e95df52409009713ea3419d670cafbcb815a97bb913613cc5f7ed5f9b0a84c6f1efb737167dc679c368ce6ed686178ef7e92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20c45f5ae0567423fc391e2a709a838a5b93c8596ca9ebd8deff643d3a0179fce23729628897796142a75da864dc338bddef2c782b68b9b9bba9cc99812c21ee984dfef8f253891dd8680b9f9898e190d7b2e535;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30d38395c815f91343d39123990007e91b38d839d97c07427f1ece3ccf05237bc6ae5ad2776aa2a7af608fa200989d78d5fb3c9554a108d0eed9d5ec03a9da85ba10946e34c224e2bab4bec3d343d6858efb97dc0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45fd0f6ea4fc4de49b91a9d8c89cd57c21379bf8798ed8db0cc4d917506dfb99b62ca5075c23c0a4677c74f1d5c0c728f1c2ecc2818976192fa3f4a9056ef332141c2afebd1ff18a179134f5899c6df2a3d53c4e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9b13ac5e5d790a17ccddb3b335f3135c4b1ef7f265851832704d6be778f29373dbd570ff8e7219c1e7ba384609c68c2ae3175006c1eca6fcd4191334a950aa06b7296687ad80e13bb73905da69dfe8b03642e788;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9506613c5eb008863a63b23050492d566f826e112798fecc0363a4ce77393b2abfe4167fa202d97ac1810bb6274bc4cc335f2bdfebe05598624936c66c5be8a8af6691fe34dd351eb48e50891b146ac59b511104c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc52b7448132a01025f2c2726cae54bbee15440fbdcb2d831feb0ed1a9dae16ce7d05ead4fa0d55b9699449cd62dc654fa4a433aa312c4e14f1e38f943da24eb2714e530918588a1189221c5dfc093a0a8cbecd55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h117be935338eb628770124491363f4c8274c8fd2d765d625ab9c46ebe824bb0283787d42ac6f92b2fcebe4c9c29aa055cb34a0b8c9739393f8d611000380c821bb032a4bd6c6ba1f975396cdaf873a27358c00bdf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h626a985ca3baefef9acc862fccee30e88f5907b9e5dc5405aacd4adf7477bf96c598eb574af08e67cb1072f0b4959f3626433bf12d97b1b4e79302e6e1b0a7d28bfc986b9e1e4d4366dd79d90416d94404660b9cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4706685b265e8261109b927efb55b8f9662f8aaee33b3f883d36c9d1eed4b724edd9fe8e097b76500f3f9bc6f4c9758a673cec962a78d56b80b95e7304866828e9bcb3f6abd914179bbd2b16e455b831543e62ece;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd81b095857bd12aa720d135287e2589cf73f3ef640b060c9706a16d56c638cb7d1e457ba20c7f023f6d8585eea5981c6d777b014ca5dda44a044560f1ac9899e510a609d75b63d29f71d78287846341d7e26c099d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a5450d18be56d9138836f5fd93caa3f22e821f1357f5f9c7e4dc042d5594ece44863e523d0f87fd5240373e703e26adf1c71247c98bee009447ecb2f2b6379c71f06db7842a5867b9abd26724e0a7b974b6ed207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c08a12138eebcf0a23c9b9acf21ffc5a31b6073587ac2b723e9b1aa9e632bb6a6013d387750dfad3af98965fb3efda84fe0bb93b76eb0b73f02e8993c7ef370da70730d6062393a456fbdb89e96d987f52d6f50d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b98b38068e579b9a36171e406a0676e19cc6855e6f2a927f87ec18fb745045c67bfc7e06044cddd04aae4802ba7f159f2c72cea6b022c315e8c4fd96af54345e88fa710cd2eda93deea4429f5a147340cc337ae7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57747a6f179389d069f9389682f0791a59b81db3b40ce80783dbeadc9f849a389e5c0f09065a3d78b192979e6c2523c03553889c022af0fd2248841b22bb38292db255c9974532dba1a5f1ef6d467538b9ba29d04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e6347be3c762f3a47b01a541c85e7280ca05b4bd24ab23edb68f8fdb1bfa9c0d9d54aea177877a464cb89138c73480c155af678640e18ba96e0d1ba132d4b4faa24049cdaf12aab90cc4306f6500ab2abdcfa42b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7b37b5133b00298b01f13ecf11e86bbb18973b29d2c7702947d6545847f736de03639d88f2c6278f00a8e3ac12c6a70f3331e214121af8cfdb914ae072f56594c88ea6015712dba3cd8c596433cda01dc20c96b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a72e0671233acdf183ebe7143c8973596ac7ddace3fd60db2d2c8f0d642ef7d01f99f4c33812a8ab96b0fee37baa0c2e23da60faf26b9d29e200c49aa1f36a87cebe8e44f9d202837cccfc23448acab3905bb01b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b26d3e5653898d16bdd973beb77d5a1129beff751e39e7596a770cf70d236d72dcd710610dc1636aafa202cce863262f6f8cd3248c725d8324e1a5bb1854d08072bf116312c57b5e81b7c648854c25261c4ec907;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8678d4057b30ee8ada5bc14f1392efc1af667f1c9d0a100025cfc3b855eb3878bdaade1b7c3723a39d50de1d1415c5f8cd7128fd94e2f6db9736810802cceee4260739907cf58c4230489ed2144fe258b74bfd8d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9943112d757c4b96f945c59f3683c277e50832b1b17b7f999060f81e5a81493dd4a31af8ef4699a3f8b76570acf994d497ea91ff4aaf44c472f60b295db95cb45707855d4c8a1cdc28b7df479acfdcd4b3edf5b6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h358bb83b260b551e2ee99ba1dda4029320f37cc274c404f5c32636b39e9a04f1b8fb2300971ce9b3102ebba555bc4b2a7a7845ea2197f1949272cd30543e1e18101a0790af82079ca9f5773cd390cddb0aebeefce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c8a78e9ffdb8719ed2792cd6ad4736c9f0413c200e6d6cf6ba89de9bb6045c57e18daab97a181b3481e4e82d22bac09035bdf303c9b8d16db993a9aaae9351d96bfc6f22eeb22a062db5beb44c28b31787887fe4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6e58e7bd57945cb04a7e3b0566889711863424f65fe8e22e6cfe7b58ae95f0c7e934b7c75f41b5b2e68c349418113965d9bd73f6a34241257b84c1f564400f1294c88f6736b27e87c384637b5e5c8f23a1e95ae0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45f199872a854760b88abfb06e8cd0256d445196e1b6835dca8f29fcec63e3aa6c3357e9aa7731995520af923c21f28a67f11e250ddf51efb912fb16016f7c8df360f590e37a355c36d83598874e4229aead0a19b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2acd89491a055e18f95644d50bd2729323ca34e388ab1c9ff27abeff3f337599270186a0b103c527d221fe521d1fce89c5f462490db1e07f6d84f7b3b5fd26f2a2d33de6640cfde74dc229bff82080de56d28396f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45961e7561eb6bffa814ea16ab78018d65647e7d6b9f2a2516462afe46291f520df76b2b34308837220bd8d358fda24b6365d2198290adda930fc444dcafc684bd28fa2c5b9367f587447742368b26745f027e554;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fd5b783b0d0479be06c43085d962f6c0307157f1248f4a32f0efa0e04377999da5b03ee75c2d8fddd085ce29e273602801be3b9f1f44b07bf948fb448f56fb006d94768768fc47e6fd2f17802fd4bb060279000;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ba8531079c9dac4ce983026373b0703ee4c4ff197d59b954955e952fa05dacc4eb074a5496187c5c3a284af04c27585fa8d383aec65e667799c29d111ae3283cdfff518176dbdd5cf441dbf1acd343f374e0ae86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7d1b1bdbfaf510a30a3b90cc39c63ee13629500b56690e914976751404877f089a751dcc8a0d1a34e3877b22b9daaf9e950c627cb8e9bd4f08517d547dfbad7a27ea63eacd6883f173bb0f770a18b3ac9ec53951;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fffd9369d0bbbed7ff8cc04ecd7a72af2426e3d4de225af440fc546bbbe1ec262eba7fb906efe275fa25f6b6efeeebc108c659e18073d60f9107ca86ebd110c3b7e9f5c4863ebfc0d8903124efaa059e362e9e3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d7a285cd5292ddf74af9d9f2211111a285c95f14facb61dad590d3eba20a3f30f99343a4407fd7b5a1392e159892abd1014c082161d6cd1edfe3f23728a1b5a3ed3e35d36a1e5c87155f0f8b27c174f26014d438;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h341c2b9ae88260c1e0e97291791b71f203b07a530fec3b7ce207fc2ec32df05a640c3bd9a75f5c19d183a93af8b49d902acabd253c7a38b2528e26bd38864303dc8b2696755aad961e2403a4639486efed490b693;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ad4e011ce8ee715ed6ae69af746861b261fa497242137d4f1ff565f02103b650e27b9c1f178f46ed0fa2d9da335756ad1ca16e23d05eb13c9ccb414b1ba78258326ae9d2ed994883a61ce082c85a4b8018e9ccc9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c969fc2a112174abb602b29ae83b4dc981dcdcd75b6de062189a380c287d058a7f670aa068db8f948981f80682172ac87db9a8a0b9bb4d2104a7dccd523bf1ac007249a3da7abc93ab12bf4468eb901299ef5605;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1197de864d4567a8a205f8c4fa0947ceb99fde3822596d990e510867f9d75b7176a7d79eec42d34b6f962942f571dea6603c3bc147ba025fabb1f7868510d468a884e188291da57589c6f81aecae7ca9c76105e2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he32a228b3cfd2b801db28b4ff3e3bcf567f0b52f688320f2e8128da415a603e13aee384a14b9d01ee4021a7044adabad6dae84e2f534202f5638236729a6d734f72a141cc92a46f72cd6f0dbe311c4bc696e5e27f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ec0631353ac9ada0027c9c576b7a41871e349f191e79a1244b6966778318ad4f89da4c913d8ddc6f8a72878eb8a5f99e83c1242fee37e839cc212c117868370cc605f8c99ed0f2ec69b3ed8d358582514b93fdc1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f627acbad4c6b03fc41256f496f7c136f2747b9b5bd1dcf22388762777651b1c4daa8130b1e6cdd5a9945372409e9c5d6cfedb94b8905659046ad49bf2f5f61f752cf4768af165edd7d49e0b2998eb7596f845f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0dd9fdc9a52dd295e32361f117926d8bea1406e26399850331beb5f4fb48e8aecf9cee5c6f86c8fb8b6bea742d73f32611553e48d8957bab294bdd1eff4665d43dd43a1affa9897c183502c5edbcc9cfe661aa59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd39da619bbea71c956b8c93b91c90b6192f0de67eb55b7c1459ad1c9e37c52fd64ccc28d961b6e4f146741f8c9423288cb94d1068d277d92e48ca05258edb67b6627b1803cc12654f27122e95d77f29c140d6b9f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd007d002b42961789d93a0fb2b4c2e034b631602623efc48c8266d12701388c42663560977781075f934b4163d06ac2d382d9e4d79e2183b596b1f9920eb84e4244e4303004543b0b72aef5bc540d4297c694c8f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9958b9d0f344468b32b36fe3a5e8e9e0900ddfa68a45243c3f95a376fabf85d5e3c61036a5b29d0f9358ef9ad629e08bc79f06c9144885682fb121d38ff5bbac3528f1d38828955815ff3adbed63f97f10dbc980;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab169085ed6fd1cc08b6dfd6b1f3b24450e2be21f201b07695dc3b56a257326665a0df2272d34bc159318b6732e98e43af6d450643aecce80b267648bd150522ef165f6a0f46f8d0fdaff3afdf6fe6dc82eac170e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha98bdf3b373a27c59cae4b9ce892bd459cb28efd251754b4440120e7a6e873c54451b2848aa616401dd0c59200e923915aa2e7d88734cbb4d973c343577a24f6076dde4ae20fde3cf33a6d4267b956bf59ad1b8ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc9b71d89d3fb34b17e74fbcab438bf5b489741edddcfb5985645756cba55a8cb51079452e734ac75f425cfb8c51a6d31969dcf467a6d4dfeba405240c0d17a628f1e7ead908ea07d4d4ed9afe9b7e6e0ed3d80c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d84d15e7e1d7bc380f5a18717dce9f11f9efc2ed6a52669308256367985d46d740d55da3c76048293a21c3956a766b8b7ed04cd31d7ce15c1480b6870601e60ca53932809572c4e323384fc67b8c524980203aec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h521df21321ecea9ab2cda78cb54dc98582cf6d6b485480b4ee2b4723dc0c736879da578f30daa3c0468e327e75ea3fe445b0b680d6a5947cf41b6582b5f7d8e5b224f0f16db610cade42885a487ce1ddfd178aae8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba5d1201ef8add80cf5450267f00f95ebd9702daedd7718ca4c4b811d830e6c92db70e4c19608fb556abf8efdac78719dd1d1085275f69b95e06e6403b4602ca22e100c2ca035e1bd5f91eac678de52d82f4787fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3096f107a4f8a94dbf8cc26f173cc53b8b7737e85d7ad7cd341e27fdc2305a94541f9595a5dbb617dbbc126809938ca1cc4bcd19348cdad30ba85a45184af1ab6a1eb42493dfcd896081337edd1ba697859b2e775;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c6c310cb1f2fe4269422725779a0380d3cad518b84c698a52633e3e2bf86e88f4907ba23f57f004b20925882bfda267613a3d89d3986eb7d3b3f4914a3fac693acd3b9664d3f890b1500cab96cc5169e5ea5a847;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5212b2ae2c93c8fcf990e3e7c79a3baa0eb99d3900288f39b2d2bd90491528f62f0dc974c474d8af50d4c39013979ed4991d18192b1d05846b0add5b4e8ac6087496bde14a36377601bae0f8e5d8642c1f7f3bdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc04a8c5e4be4659d8beb15e62553b450210a3a8e5b3cf21b1c79a55af4e6154b9887aab5be4a4217547b02152c73b3a9d14601b0e7dcb0b1621c521a96534123237c29c18171e97b3ad6c0515916d123c0137ee5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b6fa853240ed72dccd6829f88770ffbf3aad11c91167359c4011a8e62a8b33eb709031fa9f4fb23a9756e3add339940a826968a6fea5be6167bb56e702aaaf46c3618df5a22cf39996bf78944409076d21e2923;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefeaca2274682f68fb48e5506d56c9c54b8285d4c8e1e977c024a33b1ead18f42dfd3d4a32bec6f49c3e93557a8ef517f48f16c8e474755e32510ecddedcccf650551ef0c9e69ff4af5703c9637f3b93f8120f589;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56b09fc2de8c02eb93fc96037574444ea080661a79c8c7a4386829fdd36b7789491080747605a6bfb568815a3bc39e7d107859df7eb083f359c275dff04123fe60e162f9b0046cf46f35a980176e66c00752c3838;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff1805879f1006376b2483c8b4f735be46b95f3d87889af5034af2f7078bc361be4450e77c268c1bf1621b44e7fbdb73beb84b3577d0aec457f801aabeb1f59f66b9f4b9040fe924c1ef86f39d587d172ff3e9274;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24241f0848ff76e9bbf37922607e7f3806fd8d8e0e5407343acc2fe524fc68df82b4732afcdc499bec5422f9ada9f5a917ae795c172ec3d28ec866d6cbb97135a8e3671cbd7edf6752745acdaba3f9c5096d633eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc48ecec342093bfc454a77b48aea527b7890efa1e52057dc843de8e709f40a5211719f830623ad1fb852f88c87b0d3a4701855b3d72b767cec663c02caebb6f5015855523c427b23edddaed079e21f35dbe157cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14c179e16ff76a80052c476add97815e3daeb87115b06b49708f9a9ffa68211521659cc76e44423ea9c10adf4b1dbe492248524e9720b4d54ed46708acc0f768198fad1bddad192308bc74bdaeb20b6e5ac822363;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h184a64fc2c14bdd1e9d5a4d48de60762f53a47d6345ad0d71985d2ef83ef54aadbaa7204b60f50f59456cc1c842cd87d8c149916abec2282aee3b5fa1c23e8d582534ac6855b9d60869d490a54c497483f99f506f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3a52e81a149c3a0fc56e6372a8e5940eddc55bf4f1c42bcfe8f9ff7672f5b8c26df9a44241400ca29c11f9c67667ddf091513ecf6e396c9ac696235237a265008d473ecf6f0e523e30b05eb438f5f264f5b07b56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h907fde958ef618b826efef61d8258d6a65c4cd615285057237f22d6f944b2a09afea40c728a8ae2b5a4b6651b3e5730c45663741f205f02e707df0b2a654427cf8065433715daf85deb95785dc6a827520fa2ac1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1c36bf38c8b4105e42f1c4b26c056b5e08e348b4db8c7c1a4ff8090331ce782bf9709dcca6c1e8251e32b938fc0dc60124d4fb796390c6f0c7dce83e9bf9d5752762630a509d6d5fb2e5a9b1bf851deef797bde3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbae581b44c4f3c20fd7450c6051dcc1925345f511a90edad593510ae26a19ac210ea5469d462f540657dda34a0b0ad01ea6538c5d45aab0a64245b6b9d82f26faf595658db3fc850dd62bd04f0472adf2351a0f08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5708e405ad7be119d2aca5ac958fe04f7d2ae4baf7641b84f14883efc6c12a9a70b604a9dbd5e944484a86353fa6695068ebd11c0c760f01efbbcade2ac2c08de99a9028e41a7a4940777dde881c175c52174b4c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4851f6cc8884930f1872189d05720b6912c98453cc032e23ff18049a1d4ec986b7c9413fe7171736eea5e5a1e179efd6f8f1a9f275f3a36ca41cd2fba921ba6102e4d4e699411c43c1e36b901cfd8dd2c95ced5ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6550f44e1a1f15b89727578638011eac576ecf20b68bf03c53a9be4f05ca811dc1caaeca78d4c13a23d05a4794751e2d7687f44017eb219d9165dc79cadc9b1f6ee893694581488e41e731cc226e9931e7c8bc6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd26b887732d8b548bbadce105375fde026f12be86c45f45dea7b8af0d472ff17f6f29eea9522976c6b5a8322dec7a546d5c7842561e9efc39e416e0b1bf34aca0907b9c01964f575f114d88141001f31b5c8a742a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27752ace21362e91640551ef9976392a892baabd7f38f104e0c819dddb7483e24bbdf2ad32ff2e9de11fc77a084886ff53a99fac60229072528cb4baf5eb0222ddbdb2e793823182f69b3f25328bbbdc4d270ac07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf17965ab4940b14905e3bab9902ccb6941e1482ca5cdd96eadf6532ac333117b66ba43e3bf70d50b967ccefbe614c8c412366671e439f403027347230c45b87d89a61dda7821d965e951873d347d3e3ea3c8a0904;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7fe792c0dab3a68fa06dbfa8911291effa50178eedd7f9be6a172f104833afa94026826ddb47f323aac740889395eb2035fb7e84fc66cbf7b0bac62a029cbc855311b48c6efdfb1dc8749e088ce89c06cb1fc4bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39fa8cebfa06947c010db10ca21dfcc0d83a7df5d4bd276e573346683d88003cf25d2fcc640f52f65190c0575179bdd7e0df7603188dd7892e131a5476e6c0f244af239dab03b3521b12276c3006b797053720f43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6145b1540cde6ebe1e362f594edd7c8c9e62890641a7544d7ff4874d724a665710cefa54780df4a93201c69f1df0ca0ad040dfb691fd981889df98505b031f11c61f49195e2a815ab6eb6799574db3ccdfcd5c50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89ebd303148b1ec25b5af3d8839dbe4c05ff3f96f5e27d60d83075fbc39f31da0b18c8835ece0df91952e6bd06109976c684da30b647cd21984c7b6066d5f228936b9667ce7c64ac46dca8ccb10ab7ba788965059;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea01da7ae09d510c5138b40911f36f41a53ab1191336169978a88d6484fb1aed753f629ab084a74fff1baec76ff3e9884ac6b84107b61c1525ec08598f296b93a77b5e45b1fb06cd6c35492e057a1fb70d410388e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaa20773f8b10fd8df070696c92dcb05cc2b7c1c958a441999c68bfc53af27496c3de635343ed9dedb46d0ea5c70dc5c34c1f4e0e079628ec4ed1bddb5376194bcbd081bbfa0c83c0b656bc2068cd287e424af710;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had2aeb50b466ada35a7efb392268fb1e6a51b8d78fa8c686acb9d31c31323824b153860d378d7b20bf9e59d5c652604a7bc41e48121efa25b2e22f51c0aba7f27504499ef4e705d32789746cc73fb2ba178ceb516;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96fe49725501d92fe1379fdda829b8332b9f3afd95647174e2101f94f12a6491a6170e62f658dbd3c2cc4435cadb18e649cf6f493d6cc2497bf4f84a61e1c027d34fa1ea02a816b05605221c702fe39a5dc0bf21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d6bef4e007c34a3ca94e2d7c8c5a6eda5596136c247be7eb8faf1c424152893edcec9add4559eef0a6f1a7b924463d0a6adedf84ddd255af5a7129503bb3bbdfcb05074aa966f66f3a50a52cccff751a09d8489c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c165564b10081f0d090de8196fc052c0f9bbe3d95e61b42484b839380367139490836532d3f7215fc42b08d9c34e14f33c99d79aec14b5eee716d983311b95bf24f8d6f6dffec7fc619d02de8b5a8739b6cb3fbc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38f1d8610bd83cd0e16257a5cede9a52ea6ca0333e92f2cc56312179e12ca47e3711945fa38ed1fae9f7a51dfb1ee027c9b86d6f9483f8a07616dad42ebd9bf68ad64ddf03c314fa6e8c9b389d9910956444e6649;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha21ee0ba6193ae3ffa2737e84896ef135b7310854ef511f241cb285d64a5948e9219dec6c31eaef9c30a7641d419789031f2a15d26e3c2eca996f84120dde45583a25de37123de7fdf6869a47996b9e4502a478d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf691ee93549065dbcd185bbe09612f9f91e67d945273967fd400df3f28daab6e8af7eb6ca6aa5bfe84ac9c67f8ed716e5c66ba6ceb1fa092384d6245436fe62059c5dc948d7bd3d31e172d8a8f0debcee2126d4b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h454dc01bd12ae66246a458d8dcaa61501b56840d4f5aad6e78f8ddb9d4bb44b8993818869a2381ebc203f94cf13bf6f3a4dcdd33717501681e75fe2a48b248ec398f3e07da4bee49c90942c726b7d56c0b81b44d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he93e97f3358dea416a69a37b28bd059b6712e60bded3d1af288c6b09694a4b32566c6aaf69b00de6ad50005331d31f950ee25126e898a9f1b6a02f487cba641eeda017f2d34979aef0891accc61ba473d154aff9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b2896faff8041ba22945b8d562d875f486f61d579428cc0c580a69f4573099c86000828d28666f9c9b7ab7de596cb94ad5dc27b1d6d2bed5a75b274c3e576f5d2e739e180e3ce100761132667629074320c26698;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a2c75eec558e62d204ae3f187fc8b7092610abd972dec7b5ce2e347479e49daaa1666b97d2c57dc0592b5f1956a6ead76ab0547c9530a026bfbabe0ef1e69844e34ecc9993fdec54496da7fbc9968a3e02420056;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef598014a34599f79d3d2211e646940d1905b745d4d346b53d7eb87f8f25fbe4cd3e644fec435b2fd023d5a24dac99aac41872871e321b0fde9bb452957e076ae20e79b0c3fd778873fd9d28c4c48910c5c1b98e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he990a02133ff2f790b60b22577a6142e77ec11780c6f28f5e78eff94e6ed561ef802854028b9cfa11798625ff700eceb140649c06cf30af45bd2603d157603a54ecdc86fceb7a3d73731b36fc05479f56c1a78f6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d4dedb2d8b9c0919a439aee8433db091cb130dbb5862675fb6b5e577dd93b2be1fa494dc71a4833d307fb236e1b579e9355e1445417bddd60d81570ac87233085b0001b98b047765619e4f0e09b855ac55c4f7ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbffb38e35b0c1aa1077c989d70b0560ec3ecd1224b2e67fd2927dc43f3c9520c2f4109660d73a8365d31f38168d8c0df61a4c21592b07631b841398f1ad293d441d813403496fa3007b3bee357344d3ab63a599;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4533ac393aa47b5ee410b8dd501f67159b15db23ef3922c6c555b4a84632603b65c0ecc44e901cdcc2e6000370544ff55d6ceef251e1d80db2d4e6812062bfc55d6578364437ea1e1e3b42970200b332efb5466e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d7b10a8232cae7e2468cafb3357b4d80791c87573fb207775c2c113ecab8bfee08ab36dcdcf8f4753a40e901c46b1eb20c4c89a0e4120033b2768972134d0683ecdb14fc861bbe423cb890731bde782ad855e0ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ffeca157b104e62b29ea3bbafa5c4fe501863d296569027b3219a38caf437af81c760e4fed0900f63fb911718b2c5bda5db4753610623d649e1d8ffd6c9afce2c6933f602b2b22e0dbe8c4c048e2f441e669b6ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d606d69e507c1abbe8c77cf985f828849545b5f7fc6493e144ddea9bf2f3ea18695e1dcbb674729c0a3e8b2f3c3b7bcd997c7932a40c309a4e7bc0a41abf032291ba20807a295fe68b5879f611e00b56cf0d4c7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd804d598a29317ea61020d9d410c068c43f421a00c8518e949c21fd0cb34302f5cb7af07c2be4cf32569e0a57cc35af8baf0cbee8f6726258c03d5df27d34a0c5432e91f4ab58fd6b7b4ff1eedb32e90237d48f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7af51f37cd008c12add3cecc7f97dc28ef8d0f2161d3bf1f1ff381fb478fc051c83fc85e0d8e6bfae25fccb276e9a0ce626cf713e6231743365d857304643a40d4618e2beaa6483ead3002d7cd6c0dd8bb5b7813b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h663d9b6d683e1d72943fc5ce279532ea4c35c5227febb1616b90270d2a3e6fa73369c6477774504b359828fa5ffdc80b7429677b9c7ba1848250f617b8909d73d34e7695237fbeb5c155234a74582745fd110e389;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a591b396fb13704c92300bca8d318eceafd743da626658a0be2646ecc5b3793346856e370fca9b44c7824394fa4cabde52d7e67fc0d2dd200d7c98f20f6d914044d3da50d36d2a0a5c803b6952523a59800d3790;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd62d96f7b23ba2044493d1c82e68ec65b8995395a38954e23d8e497225049cbbddb3d9386a27ba88b1b32bcf2dfbe4a893b277a56e322eff075aa47037863a7e2fd98f48e2412965a5a4930375acd32e9b2290bab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4395006d40f7bdac365dfdc4464cb93dbe6c982bdbca44ef516c4c26d3d8ec0d800b407e7e53e191d8f4241757e372c36cfd56b3bcb6153206f4f8417acd0ee6f185abae8c6e159b22aed67031ba114b6f8ee0dba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92c58195492005d65b0370e7ce2e8ac1454f66c016ac1b65c8edc78366a60f85e3d54c0af708c0203f331e3756a448ff7a6c62379034f34321d84b1c0e53b3a69d009e993b1f1d14428896471a6b0b610434fa190;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1228ecb873ff992845432caefc4682d45119eb3729adbb155bb9f528f1f6b1d7987e4ac352c05934790d8c487fff4a2f67222454b5f2214617803d41dfb0aee5e1e77632f2977ea51d4ef8fc4a8aecb2c6af670cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91227124d88e27c8370403903dc99af8967561ea76704b84645a2173da56b219e90ec89ec85f315865772e02aeb43e7be546782363562e3ef34c25da79ed88964dc07c8df241bd8bfa249f53ec4807358c2f0a09d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e99f59ec787f7ca03ab62946409f7f5f981a3eded2e1880fa164b832e99ca061c134f7563032b007cb925f82970e0de7c4e6d5c4e89b7cd0b957f85ecefea7ed283a54dd9dd23da033f0bce9ce75e9139ec4bb7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62c9ad948d0ae4438d2d445662571e0454ad77e7a50443e4cb31dec3ba4118f5f7a3b5a935321d479315bd88466c89a7c485ce6eec2cf580f2e67c12fe7d00a79055d08bb671170b01a6d3d01ec431e7dcc539801;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fc147a84f33b12847d05970ef1ae39ae32e697532238d534a2a3e19017592ca03cbc1a209220e4df6a4e2cfa40bdd36f9061c0f10173e4d88c048ad5e989561d06bc068987e51f917315d01006b9fbbbfbe1fb86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb8d70377fd1e038d7a4d2c116944123c7d32253139b19e41681cf8434592ffbc73bfd5f7d2453e73e2526e6232401f582d413addddf072a1f6b5ec61125e5d83efbbdf0bf87753c6354354071b68aa28f425067b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2a3121f7d0f5ba38a1a87f3f7a984ecfd520b48ebeb6956e6872a48592e40da1e34e3a8bfcd856e7cd59bb1ca85080e00079a0fbfcab6d542ca2d2830d766eef0a38202ba00b4edde664f660eaa89e01038446fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heee0365d1601785999be51a370ac5ffe0e5a3e959eed33e3896b0c709ace3d2e46ff87d2f2475f365fc2fbee445550341748fdc7ea4b56ca5a8efe7498208c9fdc9a2149f46e251c4e8ca521fec81b1706c9e127d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3da89178d1763b890319803232e9236dc9e54986ee6a67af85e99521c9ce14fe7cf0670873e01e03dcf6770031ce25385fce88aa809a699ce8912ceda91f7e75a9f3099e70c029871b33602ff9bcabfc06c4287c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d4beb3afbf4d62e338255fe94a8e75e178f430678b63fa97b3979523362a671018d46b6ebb02e6143e28ee92bd5f6dab313bd8a54e6be1345a3d7b7f19540769eed363f963c0b4c0e5b8382fb0c188cd99695f72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d9497f031976dcf1176052945847637c190ef977cfa0a4beaa844fbc4c5e39b7db04b1ae8d9dbb918d6c44a88a4b7f841c02b945d3fae6782d273f3de699ee84700f21d50a4fd58f696098e9bbdc872298076c53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fc3f369ae2daf6ab9662d90e6270dbd1ddaa332580b843e818b84f88a34564ec8e6502e3224f4d79310c715e7d8a479160c9608d1323f95b0c3bc311690812735f9ce2a73493adf743f08151ec9ed9ba63b076f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fb14d58f775479437f7fec87f8dc9aadf6b53df8995b050c631cd77cd0fc9dc07680b3946183d47ba406b66804daab5f941bcfba33a26d221dabe443ef820aef74d6a3fb090b3ba035022ac26021cccf556eeee4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec4e1a8a0786df5561ca746c57dce16a6ba2ebe01a4dd83add9d166608655b646521feafe84f3f0f3003e5a6c67166923d814c10e7794d6c1bc2375024548fb2f026f7585cd6bf76ba885d77c5edb77a3bb0d2b35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a2b94b01d865236788ea6b4310670b800e04df2a0c2080855fd960be3ee51056e0c98125a358fde1579fa5ee30f37d07938a42170341a7325a8ac258a7b419dfc05fbfcb7e041d008032f75c654ec83921eebdb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2450e15e50feb3a6b651584c86a064a0fb79a5f3ebe8b542856c46b6b088e87c19432aa5232cf2a85b2a0ff2915ea6353c226571e1ca40ebff2893990e3f46d051652bfd75041b4aff2a88bbb9c7306aa8eb668a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebaba1d4c75aeea00b65fd83ef47e608e236a9f6226d10d43766fe48c1fa0464c25a66812068e8296edf4d2cd16cbd7d4c267ee390b45d03f09d75a49f5a9c5065ff15ea580a64fd5ddb24260bb1d6216f50f52d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda32cfffb4b6c2296c028339ce52f15fd51c2a2ec7c5208324b048e9c2fe902e0ed93ec0373e216273fa57944298774d5bb946c2eef5a964170b1dae61c111d4728d132256a74679c02337922433d7994dbb38511;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d473a851253c2e6061203522afdd68950ffd172a003f1be8ab6b5cfbb7e804ba9d10e75b9cb766b01b5503f326c93afa49b203ca90cc9453598de93b30125974aac171063fb73630cbeb58f8bfcacee6a931bae9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5334aedb4df599b6400d3d494ead7291b1dbd4ad5c91a1d58d8fd3cbf14f5dac117938b650819e883a9d9a48db4e5059181d1b6c00da58ce65559e447aeb04b40d312b903b69bc4ac333df097136051c0711a75d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha30d78a10cca0583bb5b3869ebb1a24b50d60ba389bf3fa7e477efd8f00c91f0de5b882bc652b787683c5cf5381f78a67efa0f30ca58fc38b40cfd98fc06787f5200a5f96f2c9a44d6da2e809b3d7a99838f717aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he87c93cf1fcf1ac26538a76ebaf225b4f5ffb9cdb7a1a808143a0d58b775effd286cad0a1ebc57d1394dda2bc5bcbabe178ec568bd411dffafaaf063b6a1d2e288396e8dfcaac4870988bba3890c3a30fac6402ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a4131189cca364130ab1125bbd7d1ef522cba7841af7e5ae2c386bb916b5300d762ad02dedb428f41771661969b8d5c55c30ec6f8b9f46d62a7143c15da6ec47f2778274b3f75989ae7790de3daebacaca12a503;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ee13840abfb2d3f8aa4fbcac3c58bbc2c2ff34893cbcd5c65f90dbd1cf1118075c773ba73a4160edb532dabd49182726b46157808587526030ab2437532b3f8e1c8cca94ea8d12707d4a3f11e0c92f4a71fa0f37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he483c34b1bc9ebdeef0a3fa6cba4efe91b890a1bfa20ffcae174bfe4abdd0ff8dd29ad02eb5326572e02a8f8551f7a633a64f3238b68cb93b3f209fd6625f8d0419b20fd89d8ab571a62411ab3f675c511dcd07ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99be8d6433cce383ad9c95575a71c0ffbc88d423dd479913cd083526c1620ece27dba2ed58ac0b573fe54461e3702a4fde55edc3ac65505632fb5fcf2508dad6f2982a7c2f05cf65b5232f88c77578fb0cef6978c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb221400d6ed95564535f8de072c005b0aa889bfeb519f95f1026b1f43bfd4d1337bf79d2bdb20614f62c81e49f82e6e091e2a3c6b5ea69d80806a8faa6dc65bb64cbd8237de8109358e66cd5ea6281068d856017;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e96569e209c900e980b2921f9da79ce04296d32e1b1961a0c193920bfac2b984b05b62678639d40457569d6f8257ec8930b0c6d1e75ecd4e15ab2650f7636e1164cb349902886d9d2d1fc560ba8d62cb0e10fc9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a3a7808c7e632df76cfa30b24e0881f817366c64541193b823771bf88cf363607001b59812e3e6c4eeb58f2ebde6388d732b0ebff4083e82a06656462d9d6f0e651ede1cba887f1d9fffbe6c0cd269edfc48d7b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1661847ce53c2ca0cca9c8fd89f381361cf7033066f9d3a0cc2d712845765a1fd11f7d1b23c396d09c9b5d59e67df6ab548dbc2006ef7a421d97abf037f307f4a9d7be5eb8def4dcdbd6a0e77e8a30c81dbb58c6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4c24487c8d61a6da20f36f61da0cdd41a0cd177c4d55f5334de8d7a020855a129ecfe386cf6458c5292eb7a91c58f410d88a3ba0ded821caf172e208df3a0614f8039393059d52b68d1dac1f3645b21afe64e79b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ec9be4512b3fe7c6e3dfe81c024f716da481cdda9ac4b316ec09af574b7a193bb4a4515a5fa2d35cd814731289ae2301014ddcac9eecb780aa751b8d2a6e06cfff7c8bcc70e4fab538a750eec535fd15f2f704d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d39cd7123cd00a747179a4a1ad391c87b47d8581a7630a588f94b147a8928cb1b436d7682af593fb7e498128bd0f4bc7760e49b7859730bd561481942713d179dc71aff24c77edf73e417c181aa19028d08baac9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bb93de60768558e814df82bec9c1cbd93f2c6064e6645db5cf2e192eb815d9bd5da5015701ebd7ddd9044410d74da17fa16cfe311b2c7d5a9cb361c6830daf3e0fc418f8420c8a0da668003bf2422b77246618ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bacbd34d80b2e6f2c85016c498e2185409c7571763b51542ad715ac8de30fc587eba684ec02b43c05b5078b8e0547373298adfb91a0992410458e48ac8eceaa2b8d8803a79b09f96512d27cfbfa9aecf86a22c01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34a6ba861cd9f820833dd1d715e53fd8b204ab6524fd65f2bd7fbf774695df76da50fc7e3ed5b826d07646e7e94685af9b44f50b2d917ada8bcc4f1ecf20df816c9ebbd2aa116f2933b45b5ae6f29f70561a53fea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fb7c65789d2d477151280b8f8ead30f0a52a4720d58a348c34a355ecc994bb3d8501be8311de0db06c53017cc893732778a17c2f762c88f4541496abf3d3bc59d548e5202410cbe1fc7069030acbf13f4e5b801a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h234e8dd1bf9fcd21b031d9aec5c1250befd5c51a7be16fc9e3ff83f7e1d1b450b6eb2750fb77df1e2c6f599c03d3e5ec6d31d31b077a6060c00300eeafe3de6c417e8bcb3efc76eef68b33d596aaec1b4bd29125b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf39350d57cf4f57574b246b559141e5626821ca2296a4e9218b9510b83701c28a78843b2d011c8ff7bd665cba376c35ed8ac36afc6a9343d1d02138480da6bba2d987613c0bea10c8bd0f26bf15aef0dfc0f3c159;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4215b62f722e8f85730f28320968451ca60d94ebe1947169fe9c415b71aadaeb8a098abff85bee6b94f1e2abd34eaff6696b26d4df0f669c329a6fa6394e997377abf3af53eeb0d574817203de47f86a90825314b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4adf9221e2a5baa36479f0ead39f4d9b4b56c9c88e81ae6dccf26d95be09e34e16da5b18296efce35d7c54aaad53f9f4530a163b0a8982f488b4345bd421dc11ffe167fa1db211c007778a6306eca6f05f147d670;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99e0e116a0c33a39d7998e851d78ee7d0d6f4a9509a9ff6718abb12061dd504b54893fa5cd36c659e5e1d960efd214ae495e2a2ca5acb2a7c55833f5083989a255fa2bc41bf91cf4d57f94b6491ed4b440cd7ecc4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ca4eea42d2d167888d0c6e6800a5bb52ce86729461adb36f135eec5b92f1553f8f039576eee40a855431b764640eeeb206aec2c803080e13fac4572a29debc9c9781bbaccd72237a99c04066a28fb4f156df63ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb68054f9eebf8a5da2f672559dcf690108de37bc84c2317ca262bde0638d9f3748fb9262cce59e3d38d17902bee8bc59520654a545caa4c80c48bdc8bf6a3a8060410cea21aafb7b6608167b6455af643d63db;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1a6d3bd3534f364ad33de4309c44e5b03774e00a53a78174518f689cc46a38e239e2273742239c333ee683aa2691a58265dada3737061d6737bca13ccde7d75307a6f41f8653015e1574d583ea21a403989eebd0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22eca80e014469b61390eb0702222e7648e3c1abd543a9c7b85dd52892a68cd3698c1897dbf25f773414a3b086b9ddfa66d3e076863cc6fc2b96599e13a2db9c6dac3b7fb4f073bbde4f353465a11718f891418bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92c885b56a1b9807c472460547215f1dc3d28fd752d50977337926c5799e248d44fadd159dad40858fb5a46581b47d6d56df948ace370a243b9fc797283d9d5472c2b48af0b39f082b5d028c1736d7216582c3220;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fdfdc3ce92f8a2a31b21d5333fda9dde626851eead82819ba32cd4984fd7a2d2f63c1c13294eb597759ba6288f9bd77504a3f851f4ec8e2899f2175f90dd3e6410c42349816317d07432049bbb0296aba1960973;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fdd09432c543973a34b8f66aca93b1f151bcc692cdf89bf7b60272ed814323112c02f22279aa662a8724f3449ad33cc2d0c374fd6fca5078293563f7d173290bed824bbe9cb42f7d41d803dca156e1b24cd120a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5a82e753dc90955304c62b98badfdf1a5b97d9d061b91a0bdc8c46d1a4b2feb53cb93a7624370279804e83f457b43f1925b4696ab0139b5f1fa2ee44c13cd3168333657751f26d8efdc3a93d684173b60ed600ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h648c5c540eef359381660dfe6a5d3e382b73841708f60a5bcebf471d0265cf12ead4f5f7c6c460be375521743be6c79ba741e035a068877bfb58381d0954df6d5e9e96b5be31d10c8640919bb39801d1e5e493807;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf93293b647ed7cc6382d4e1d9aeefd57e5b70babd66387dab6d2e79d2937c02b768c2b2cbb0901e051a63a753785ff1fe56a4166d1630b69c6a92347ce63743aff40d66a782b4807160c3862e47e4e72225c58d51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90398bb01cfedeb454c9fdded46850075e2df9beb53b4ded90863f906a9f227c389ef2967b6b03c5eb0763f6915bdd1104cb910a0f57e251bf330430b3b5ec9c1c8733aa8897a0fb98f2b41ab32ce008999cfe87c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6899b16f0cf08be6b8d845f851f1f9c67159d95a37771b858e8c5b0a9f388ddd872ec825f46cdf4ed328beb48ea528d371061f43da98ba4bcff3b259c371e79d17e2bca8058d422b60af538ce31aa98c12b06ed2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58268f02623be0c4782c193bd58325ae9dc326b1a731013715faf8c5bbb1c34bc5f741670f59af5ade65f659b7a269541f97677838097db5e70988861634d2cb4b17338d3e804c0776588dc1fc5f039bf80fb1027;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2ed04dda6a3609771dac693c0bfeec4524fc7bcde88f50dc162dcffa365e5ade530795f3e8dbb345311d3e512b8322f967e6d851bd53e609de0a88674057bc3509b9ae33eaf0ae52392d79afe01f922abdca282e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479d7ab802cfa6de092af0407d59222fb504d2f7cac4efe327ed579140027aaccaab25019edea7566fe5496b7dcf3588f3584a6540e0e8168ac1d4af7a58cc275bd86e639f64c23027be107b947ab1d265c8067ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3720d813ad29f111297a2d1d8a9ecc648b709afe14062ce8cadcf9d052cc88c80c5c7520ae54858c6e0afc6e6427c9198e0f2e0e085f1670623f7115c645c2de9a49618104c73607b689c92da7af7311d2be94edb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7eccdef0875c6d6ab0ada7a60aa421ee6b9048301ff49d508a2ff0fc8abc470c8d8e7ae9b6e0820b0d798e8b18cd1be53ca299513e7eb8ac24b91e3c184a3896e53e067b0efd19d32e9527c4c8ef5e6f4f22a87b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79c00ffbb7cd9df4bab35d83ea50857b63b5f7c8a4daf93e2f3de3e84cb2f7029baa054d589f64913b160b7d87bb4eced6e321b16d5b976ff9ce3f3a8966a28fcfc1f2451931ee795274a150321d2c677ed295fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8471d15d06565fb7f69ffe48192fbd4f4c17ed1aebd104d561682414682857a81b23c6210a1fea93a45081a48e1a6436e325ef6765a30b6c4813c2e879e3f9f5c5770196a96a168f08631a0c844a6e5432fa1c97e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb0e6966b5220cd56f1e7e2746596e09afbcf652ee0b1cb88239fb603b09d43de2046725c081b32e6c5da04a56a8b452c3d6f29832242ecfc3fd0ffe7609aff7944a06fb5ccb939f19052e4d37100cbb9ab6d7019;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84b148dc878b6b2f23f479c3154932bf1496a7e1c84c167628f41341dd8492e402dfa92c212a606f887a3d4b8887c8c403c48eaca0e04ea7375fa82b9b3eb5f6f218ffd09abd3e3a67f8ad62bbf387bedd2521c02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf12311d8ff20403dac80179ec7ae66e74363a755e63500435e47b89b0736bb3e0368f28c95d031bdeef038e9eb4e09532b1fafe6849f39d4a5424c6cfabce4f3f1b3fcc53bb88463648c3d003a768e0c18efb97dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd363b0afe7c07d59aa2a27960894e3cf1ba4f4bfaedc981a73eeb79cb5d12e1547718d90c270f12a9b0959251ad166feb9e6e319b408f8edc2bc933067735785f03dadafd8881787a4adcc5c3795f3edfb66ca0a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb607f372ec5af0a5cf4d649b560c7d507f3366fa69e73eefc5ca4d39f81396bc10e09e085bd65067e099c027496260a97d890b0e2200b6dd4041987c77aa229a4ef944f08fcad3238ada8c5054baf9d57e7c23146;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f05efe107254a12128703f778d702ae550246b8ac72857fdda6911a2902fc90a659fa67d2847f6ec67a662327fe3fe427a0a5239351216cc66ab46e2b391085514e0b0fff51433e4e074051e1ad36807599674f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25897fd564f88fdfaaf5d5139e5b16b082cb78ea3c6a14bb51f329acd711d62de7290c8d755898321f9a088f4375010d259d586ea14a792b41ee2d7a35257e7e692e3111da2469f329bbd8bd1a9baa89db434798e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h808ac9c327122875d5bc3df7980517dc1bc2de03ef6207f3fddda4316022c28c54b6bdba7c913947f327ac32097ce84611b70ec16dbbf65ee4bb5a0ebe5fdcf70bd2cab23cb3b790d24216d1fdb55ae9ec188ce84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ab841d3fd4a2623892ad2b0918d22e1eb391aac1494c3301cd6ea08d94a0a73959c6b541c5e22a0fca536ef69ada15198ae47e80a3a565b3e59c32aa7b6da0aaddf6f05fe01f1fe114fd9d635b0c3920cc4794b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h512e0702bda5f26ad54e56f0920a885ae10484cfe8b62cb47ffc1783b7ee584c8ba04dd93e59adf2dc9b952ba1717221f0a2d4ef0371b85e32bad005171713f19be3a083a5e6c9f2814af01c661387919d79eb569;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h725704ceee1522317b8d9fcaab889bc51d139d004a828cfb4dccc5080cac35c8cdca6c8db8375de6b44967351be9cee3193af8f55f9edee3d932f3bc0734193cfbe72ba23310a440348bef8e28854ff2694b3e8b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd03d33ab2ec5dd56702766dd094f0a8d9c2a513c345dbd6b12bdbe55f3ffed5e5313aa0a291c358358073dcab4393c7d157ca826b405ae55675f48ba84080e71e374cfb9085ecb88afca1acff9dfee5c089f08fe4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2a7a492c188ab1feee949cf4c5e124549ed0379425c7445bb418bb4dac10afb92d78af8df0c940882990cd82742dd3bb4abbe9413cc957aa08e1689ae46fbe4209ac40c2522999279445c6d3517d951eb118d5a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f58b4ec8470c54a7f817f50ea5b17a59cc9922f85a0bf49c552e02edadac4a96df741fc2fdc75877731224f0e5014aece6e15da5d87f4b1e269072b8428cd96b0397b6d19ec49b168e0c448912909ca7dafdfe36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3aaf9dd179bf580c338035994f1b53b58d55ebe338116ae7b8623af76a2908f66b4b41e1821c0240d91f1aa92c88bad76662811d6d3685ebde7f855b6e026a67c0520b35055aca34a4f7fa7cfb3ff4037f072080;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56af7e05d20fbea1445b9d5a7657eae44a51b066f427ecd400d69f4405954a06321ca825c8f8f5599c22f8d466a81b0731bdd4bf0f1f7e30cd6099c0da8cb4746498933589ca7318884986b6979be29ec53643b13;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c1c6a73a118f4d900ce228879ed25e6067d6ef4024a465e2a2993da543b9379846b53fd7fcabc5fa3d38f729633153e092078c0975e11896a2ca94a1bc999195f5039dd32341b70b0e48363942a3cbc6289ec8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fb70916f250298eb0d4f240f12631906cbdf03e408133ac2033defc6e16296a9131075c746de147d096b2933c87ccfeffe3f7f86d8975f718c7ac7fb47dbf9885586cb24223334a44d994131665a32d6e18d8ecd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he03cf40c47645c7d10659ca1971a6cab03f1de258b7bc4f4d9ebc5a7d3a87fda26d64be4c4baf8b79018f96016d5093706f619e945796712897cafb14b19a51fa6aeb109c9611eb032112a4f11c4e0ca64cbf7c00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4964e2c3c5d330721c3e476a798bcc61d603a147f1c2d11ae525c1681a585b9d7f232d444161ef2afa6f86d659f6c365a043f30d49696240cfdd31f1e16d348f2bb815d09f26cfc8ae611c281cc62eb546a94d9f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e87f3ae934fabd233d1bd8cda02df9ae744a6b96c0a91d44acdcf1418669e7d4b2a4c9820e4d0b551eb65810981161afd76231270f52c2daf2410d63148f275c9ec27909e8ae32557c4f407601bcca2dd1095233;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a777e6297a7d77f17f3f39b6956f30483b7b43a8b96d9697d824049d853acc459ec8ac9665d972d36da77aecbe03c65d757ea0950af81b63e0f9d45aca086036f8db2061b7f5bc0302011c5188449bb4688fe7d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha14b73176ab725c591012bad0e1b0a6acf11ecb535f2b73b3dca2881c63d567af46d826689cc70c44c7f67a77a9bd85a3dbaca7529944a8b2a2801ea5c0a6b2843f3a9d0795def1af78011dcc1e849f8ec85464cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae511b33bb5899a163237c8dca515ff968d89df5deafbc1340efc53baafa69accfd7efa378253f6aaaf212c4dd3a476909c81406fcd3e2d4ac041b5447ede699aa22c467df9e5e07c2fcd653ee51c03e0163573b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32dc782a33741d8a91da9090bd769d449c79e9472d137258ff4f777054597d9261e0503cb65df25593f88a16e67ef0d28638758cd46986338b448fa38c352e50e5d7a068e7934671be9c6b682747657af5b09615f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5aec732c4e0f4c81f6c5cb5d69814b2ce48fc88a0508f8de94f9700277a9681ccdfb977f45a77e06bfa1beaa22f82e43fea8c5f4cda1bcce83c43d53c867e71978a5ce200b279293658581e056a4ea725cb997d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h633046e191551ebabb674d0f4c936eda7fb4ab0cf5d867337977e5b857e470bc5008fbc2397aee9f545cb4554f25359f8dea2f46bde3ad394e0d0dc5c104379f602ddbef08fd704f0640ced74a834a29dfc9da144;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2bbcc15a02019615faea09fe7cddabd4be6fcfb520613e71dee3188aa544d1fe57942ccef319ace5d2b8da2bc71d07d9f1b6ca77b9a5b043109564a320354c79b3dc4c8bb943a503f7c4a2b52a211bc0d9c6b838;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f1d1a6e3532da459eea8204b921991407cde3cde923b5e856ec3df53045f8de31970e7446b0996395eda9f0dc0d95dd6def66c41f808bbae03682f9ccbd116968c687943bdd66385a9f38bf18b012a0001cb5f24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4ca9564ef468dd7fb41871fd4f36616b72f9a78a0e5b35e5f04afb20d07a7440aed50996c45500a8b73df9dd69ae1e283a268c7492879177f969689fc63d8ff4c45fe5499632341a3e2d2dc2717455dbc1eb8ed2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he73b1bcb0d67afbfac7c2519ae242205904eda527427f0d2a6b5e7db911a0183fce47efe2dbf6eb3ab2fc2974c81a5b026ccf126d685031809375b6da2af05c04d341085b1e0ab24b0551db68920576e3ab452d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h724dacef9f19058b45f75d90731931773ebe23164d182393e64197c8ecf5a0e334f11e414c40136a60b506c94956513914bc86727d4481ae905e0c82c099ccda1283d53c195c5000b2e81b282be59930678a79ba6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f61276106ebb3a63063fcdd9306cf97e9b2227cf3960e37d24ad014183d951fc1a5b65d958780c5797f00a256fd8eb0af7edb17a1c668e5414d5b25144b14d904e7186ec8181893a1217cdf5d88b3cbd21168fca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec53af656a1ce50c3f1ee0c909f8e55f2b2ce48466aa72f8500f6a8f9741ecdeea0cb76d6777758580cef4487a432454e4f1cd8f9a7a169b9c8d64750fe497d19a0f90ca4ec731fdddf84b0ccfd8d873da6002d4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd15bbcfe71e03efbea5affa9945fdf677a92b32663ad099c6ebd5b4a2600323a262fdebd2cbd5f793813817f50ee2cfc7e39718b0132fa0fdf21d9f7060b9547721cf69416d2d67c71c11ee1b3e8817317002dac9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccfafea95e38920cf3c4a3b62ace187fada2cc8768e5e416c32440d28e172b3eb787ac38eff446ce4118b3a13ea5c2593ec2b4640976ee2c0f69a488e17235c69bcf06c9175ea791645ee6797537cd41476a1ab46;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5e981b5210af1c4ce51fdcd87fcf6eeded2a4904188816e6565ae40d643d5ec320e7905948b2d848f0881d63995de5d251d940c0da6a425bb12372d5859ad7dc8d7ca665641f3e75a357af30b3a88994dd56d93f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60429c76e96bea425c81e46894f8335fb75cdaca74c8e706f1d5b2f5de8477b76fce5eb30c6d8c9a8871932e66edffc34491e41ba5bccbaef9f3289b41fdfaf13e22b44df7894d0e2ed23ddcb1be8b9a2be86427d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1675e1cd1696fb69b624ee25342539e53a350406a2cb9b0879337a7aab5e8f615bb8859cf0469375ae214f3fa61882fc53b6daab7ebf70af902bd59b405c62afebb9c006fe469356ef36e9c2698594ffd4d2a7b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7800f0738d66bda62b022bc3bc73b395a2ad08a43850090ba5dd11169a48972f1b11596d8d2a4564f29908a7bd71090d10be096bc95c9e12673992c6907a02457e9cc6e4a8dff5d7bd63a96fdf474f44eeeb74ab6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29bbb42ecff6247272e14e27364b1ba8dc4f3e5e3ece281f90a896d4847ca0531d15c8134a9ec992d81d4c23d0e2c5e23dc0ef9ebe45d980de53a8d85bcbe40e80b15a3319241f57aa5a8c2a0cd64441ecee82808;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ef11860a5b0bf7bdfad77633302edb9643b3b2fc3d35b7ab05a9584cc2e114c15478874313cd2070910cea2d0d4fe8ed78a713e7307fcb90342f31ee3a66976e6b01de93cb4a42f44f42cecb4854f24c8dd0bda9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc935d8153a561150d2e1957473c2879e6c18d34de8260d86524e430bd046532129e1c21de0a5d8d1fc9309911860913a1cfce4758dd937ba10d81693499ea36d6a2839fa53fb3f4aecc4ebab1006ed1b2cf91c2f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0c73cbcc97b23f2918cc00677d64d936722eb7ccb085a9833a2bf65e6c724f6a0fc052cf797ec125eb74a56df0a33fb19518aec4b589308f34ea434b32081d77efd40a580ea3b721af2bf922be7c4d9fdf89c8dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbc3db9971e88a97f71930f4f7963bb3efe61f4e400e5a7fe4de6b4b4fbdf91c196fccec9182425fb33a498d69a98fa4b812a67fee36a498b3f14511830162fd4bf7f06ba53b43c0313077265fcca2a16f707b678;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a0e38a3e31dc9175cd3653b8c36d97ac3eec2bb9679a3c48e48b7eb35c238cd73afd921ba1f424f685bdf0e43d4aff3246e34a01f9768fc653e1684004ddf671eaba6bbb89fa20156f22af4ce979d88a8b7995e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1ead1fdac8812cd79e4957d31727b1b193d3abe04299fde8a0a77b613d070e17f725f60309f1f2e850bda9cc19e7a052c8b5886da8e3495f28b5f9586de60f2881aaa26f53216e227df3450b59e781be9b0c90ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h503c453806c47f4d3030a8c8e8566e431c6a6c765b540595b6817f02208f5875c963b5c2ab260500bd278fe00a51d83d523c950b4067299290783ca07879c63d7ac9cfe65b057baa5a5124416d8c22cee225ace08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88b5c6df53a671c736011e1a8638430cb64f55990e09ecdb6c585b7c9ff753dbbb09ed221c0920f9b5f951ff05e1779c5355f7b59a58eb6f83579d4e7c47cb31797bfdcab6a99939b92fc9a5271c0e2bedfb21c87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha30157e07d11bcf2df4738e9cd329830ffa685cbe67b0c35e80eec4bd7265d7cdabd654a59266d5a9e51fb6bf7d680dfe66400f8a789b38b3eb97b4de5ff8f8fcfe35171ed8c6af0287163738e045058b74b30462;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8efebcd9300af78e47a05c01e7fa8a15af46df23ec1c9eb7f330206f9b8c7688fbb98d740972f22e8929cc6ae6dbd0b7cd8d310446f322cec3e998f8151825a394004f0d8eeb99fc7ce992b9282678ef27128af7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1f43b920680c292b00fc709149e118f46c2079615a74a0b6e5d3cda2df1e156972b3295cb4c1e44a2ff68d7a6d6a43cff1602f8263290c3fc331ff24e14f1c986bff5178367d5c5b35318ecf452fcaaa1bc54f1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5d8b9a18631fbee2aac712f8db2b5f2c6030fc1c9f9944ccad21b4b0c75e88a457286623bb42464df5a455a655447a75d5bb8a5c72c4ed91c0aa545733fc4bfa835a14bcfd7b8fa13b7ac7c723af470da4b89a24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8d641e0d06d68f0d76f704bb2872eb8a65b2b4f6050d528b87aca3807af7ccc8511b91fbc34ea7f1ee8f6eccf6c4a984467b796e3ffa45703778b615237b3fd95f985d72f33c63f2e8d3ccf4d03875b55e0c9b7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b7467ce2345c7e8422a539d8b77c902c2df1f68bc1527efc04822ef7a4faf134e58fc598a0be419901a216993742d13f89146f031ba9f68fa3d62e6bfbc0affe692a5883ceee0809a3685cbe691631dd459022fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f15d5bc37822938d296047710140653ac11e953da853bef57487668fc50aa3022898d5325fa5888bdd5c682e33944fe02b54652d2d9cad0e4239b8845761d4e3c7afa2e92d8e8ae09099f0912f65640a03806540;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a1fe474f7a01b823c3f2ce3c564c4428ad2e1e3e463ab0033da11ed361600cd22d123efd23dea78ef103c1a5230c18ce4fb383c5f12d22b263bc72b46a3892be520b1ae5a20a558c85abf42b6393d72a336eb6cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4128c44e410d4eda1259cf4b15c613385cdc64d3ce2ab560b0b2d1ce201a15849e5608a693e7dd6b178f87013a0df110504e14a1ff6246e14967cf7ea786fb21c78caabd8802cb07d5746d0059da9835490a534c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3c8c3fa435b6cd8f9207809e07bca21179394ff77bad535aa58a6113981453ff465a732bbec4e1fa6bed9fc24a59e06bfe819a523320e761b63eac54bf3c11779a2ffe8d0e6650b93c81b1f916d36ebaccbe313b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa3f26aed888ef6e3634fc9556092bc430e827d3091b3f2b94890aea9cff4da04146fd1bd78916456b4473b5459d5250a5f65aa9af10a5309c1cb0e11ea4402e46c335cdfd90bec2758a1ad49fa56b76c508038f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3eefcefcdee39207577371e1a5eb1c7f03db02e0b7690ad72a6a90abf20ec4d3a2038c5c3a566657b9c616e971b59d37d9cf8dfd096357b871f5dc8c418157a06375f7bcca289f18c8f0a6383fe1379eb1c0bdb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h518b73f296d38d72dd8df487b7b6b2898f997cd7318cf7e267b3e789e457cb513c82b05254e291eed3109c351f5b1dd6e9c9cd08fee5ea12b82b6443a316de36a52b38c072b7f2f74b253342633e8600b67d8edb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he62fdbe56a9a04c4db5a76bc3bdb7815cf367c8136d8806322d5553e99ffae930827cd20593ced26e6f65207dc11c9d13fbb8bc72869a8ab110c18212437bc7aaae6d92e2a00ee7c30b41e3a9c3b47402c4e4fda5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h527a497ee86a9cd947b1a57afec19b01fd2648e5c3107a15fc5fb00c9091fa98b4e14e48300ceb16d1cfaa841d9a310cadfb37ee16bcaa681e43e3bb3e3c12edb05b0161fc3673268ba09e37d1393b7adf3f5818;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19b557c78a7aee955fcceb8ea939b82601622ce0f06f3e13fb9b5e70f3ff68e3c2f3bb933bd9656ff2f576e9512d23390ceb41119f43f38c54c23832ab53859c52eb822e0104b0a87caa5e765b7f45f610e110ebf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d7f3fd3505ad01b03099581a6f7cc3f4b2c3bb051ed252760b348c4ad1a87632817b1321ad9682ea9e61a6239b69c813fcdd220a06f25cf945aff12c964db5e0ff625a6b9a947f3ac359ee5f1bf292b21929d03f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h461d8e8767f8d9695052efe322dd78f856d128e51035963703917d80fb1f9198408fd057afd417f2a546916242000b9c0cd3056ee81cb96ff8fad750b47fbff340f74186196d8f7365f5f8cd84d3c9de6745ed052;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8882e0f2abf63217af2b01024ca2fcbdaba1ca1c75f33eb1ad8e1778d2a84261a6f0198ecbc80fdd93193e7a5ed94cfe875477e52b4bf7066bf18b6e96dcdb89d6ea8fc5db3c62bb7773d4c57dc316e56dc691d74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8e2069168af8e5fceb83696ae58dc9d86dbd6622a01cb381ddbdf0f656dac7ee1b20f336b1d8b77a697580261f6ff148c605aaf1149f588db306adfda17e6e2bf95c291e0a604183bb328d59da7844fe145bc2a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h255944511fb7da80789e57dbc585ac6e9dd1579ed8041db8c69bf08dda64d5124e65f74b564d70b44f596a4d14e338175b3da040abdd7980c90bba024ce6d51d8e15a9af085266c886235f4fbac9004c12bf87df7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba19e43f9676a36ded534c61a3cbd8244230a351a56d964e92ac251e425918204bc16dd560e8cf7167c4e6fdb685d2a463ddc708dd116c6d7d69a39e7c451e95e47b1490e74eccdb8eea787c8de9a83e8f680792a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h161adfd599ed79c7e2ce8d6dfd425deb31d9a9c9c68aedfe9d1d8e26aa93ed8d809e6873f22a7f6b9839541a728d28fcb6bc71838694d1173c38631cec48efca2f6fdb24df0ffe140275b6f473c2c83f69a968d4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h743ae1fa69ff5f849239d50c6eeb0ba3fa1c2e1d1122676cc551bee9b4f70ae475415a5b770227f0c5f269e7e43a0e4b55c943c587010eaf1b7212b3e328f4716087c63e5748abe14ded1b28bd6f733bf6d5be4d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d2de03c5e54e6913cfe430c5a2e92d89f466c7709ea7493a7707e71a03a6dcc07089def32e3e450c2dc90c2a228da35201c03a2db7bec57c76e226da3ab3517097519b0b768bcbce175cd1bc15a237ef4f064581;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26d4c5c02a39dba0eb5f426b989efc863f65f4ca611463f21f829ac90ef2a374ae8aaccb2044f95cc8423b00c263adbd91056d143baa7865f055b56b89f4704f63a933bd90246d5924211102138ccafa3a5326a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a499a072f794ee3147aca728fabf4fdacecd01579452a3bb5089fed40a6a082e03be74971baedf8b9d61cf482b8abf073a0819c40bd66fe816b6039c35dde7f4cfe1d2c46874df1620f18fd7a3c619c1b5c7c2c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h611ceb9e8d9b1869e82e0bc7e5ed44cb843b090b8782f5c9115c2bf4bab6dac2fd58bb1c22446264a066bf873b1abeb9d1a36a3e8dcd3b87b9f81fe1fbfa5987b2ed67c20989ae88d102e09ece11ab01cd10d2e72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2a649b01ecfac89c0aa6b6f18824da33c6eef64f0c687f0650790ed5f9d9e6c05655e38bf8a96f2cbf44e563b170acebd6c2f94997902c18bfd189bafad68a7e6d24dde1cefe1a016b1a14a4d8cb4bc4ce86b953;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2361be022c1e4be5f597206b4552807112e10569cbbe40a643abfbd242d15029684ee594f073598960c6c76bac1034cbd21f412b8124c21ff1fadf7b47898a84b1b3e9ddab9d61910b5f0fdde30931f2741802d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63b3a9b2adbea55ecf1d30d77dca1676cd9c54c7020e377faedc7c7557ffc822b1baea0201a7b8699428ee5b51197f36bff0b7f3594750e1d4a49b2986e9d333367cdc9ef0d475d81a68bd7f5a6352bb84ed82e94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6c8202a2b354fdc435d705a473bc673736c4906a88141888ca30c474a2599fb931e28393e6789de33ef6570f2687a0360569b36341e88b5d1c8023d355bf2d3e708b59a1e20ee72196d56e88fe169745949d04f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e76818d9a9ce408fa3bf8ab1cde024ac0762b15d2c02738d4c210758cd1fa76fb93288a19cdf75389eedbd336a37e646665941816be8260c4fe8a9182dec37dd1f9a6b52041fe9990cf9096d0ca35b4580f0c24f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefcd1fa54531fe8290afaaee2deadaf521351ca37ad6bed5d280bb9fb2b4129b6e7627b2c1ae0c9bfb2c96ed307dc9f990b1f1e934fb870e1157e2124e5d45a5a51d34b2edcd39997bc3c72890652ef58396cf632;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2eac8b7cc3876a30fd47941955fa0c8710e423885681ba693854700b9a60fbe0ee498d7106e724f5295cd5999a8951ca8cb9f75264fb91bccd4dae788c81cc58391408d1c26ce8934a90ed3de0776f1d0be0c62c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a4341e6242767a2ccdb1a94f4e3fcbbccd3e21843ffb56acf4841592943c3e751bdb308552a21bee48247f4b4fd420e03ae61d18a9f16b897df8de982eb5f8c01ad02c70d315e006cc487a4f3a9535d2587095ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17556b41bc40875064c6fe4ecf5d5eda85f6ef13ef5b1860ca121c1ea070df273b08342d84fc68628cb3162467e535c106c3f8ffa52846e2beda49855a411a1a5ea13751af8295c6e91bbdf95aa1825867e9710b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbba84041bb62b5d53f80fd6d2b9707dbc107045e65cc0b0637cf4aba70e6120e9399c99b2ca76999763a9099f1e21199edf457a19185dc0fe0ad2ad9cea16f33bdb80ceb26fa69973e4cf0450abcd444019538c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6473e58a46156c9f7a3f3907f3643327926083f70ceed5cfcedf7cf33d72cecda1ef73cee62ba5b82f4864962cb00236deb5f97f5261e8304aeac0e005007c6bbd3c8c945b4c1a2595c46044e81cea76b05b208c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfd1bf4e2326745189102ae7cca6c8a0861bc7b8ec2b5c6f9054457e6650581aceff5f065df3c1c7cc901abd4e75b10aa419036d3aa4426b35c002b87d42c79d4813e47463633aff093e2bd10014a87c1eb38860f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf87271351fd920bb4b6b8c1958c2fbf5cd3875d05985882fbb6bd6b6196dd5614eb738f303b87624ef0459f8b8a055fece512af30f2d3e5b9aef337016c5e43f58eeebbf03f7cb830edbcfbf4e9ce89467f0ce27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee9f9b7fe2f59c4702efa2ff2f4069db9e6ff951540ca3f0d35a46371e9a08364c97bf809e71adcf772668005771b4b04035aa613f17bce1b084cc3b145b0d93b460c90aa4c870fef18cebd1cdd878054ba5bd679;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf27efd1b047135979b3c4f0fd79ad954946c67e3aa544c4fe910177cf3337e8f814a0c181ba78bcee274b0004a1b7d775b346f23d2514666de49fae9951d17ca9333331039a960561abe497d308cd4b00a58ff432;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50604628b0a229bd46bbbe816241376119c23c5b1f8457471bd7e03e412aec3e6cbad37d645b3d1f6663bf345e5ec037c8b839bd1cc021c9452889a70cd3b4c464faee6b3e5f73e4b1205ffd74e34eb3a9428dab4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3370b4ab449b9e72038705d0907c939da811bc8bf93677ca7dd7ea634974c800799a1843fd64d1f79be8789b316a534fc9f73150d92c37d07bbd4478e915f7a2fb464104b60fea61278ae0847f513d09b9fc102e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbac520e1aec518f72d542ba80d48a267d1f307fb0205d46224cd6b9f2c876e0a53dd1301e13d5f13b7142e76b0630d3be91543a0d07717e98bf0b6258ed8b43baf42d5c65a4e987506f83889890adbc202ae7f10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47799f523e3a42d5ab78fb827fd208308623a5fc083d3fad4a5565ea8f4aded838419c1e247e79283d809015abf95d1da3bff6158834bce2db39639a3d6c1c1378fa67a05763b8fae985e08e11e3c76fead67fdf8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc0da2a3312e7f9f43303a1ca02cbce7a623a90d3252b35156e6d2bb8fd5dba94066079181240e562db524d422a02e2c0a4e9481eddc3c71d343c09e8a6bf8c06b1cc845db976e571ae5c94f32b2e4ef244c1e65d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb8f35b26f996246da5ba868ad1310b17b2f752f8940b696fa11af6c88caca3402172df3c5113031d763a1de982ffc67e25ad95bcd18cfbff56e569f6f9f9258e7f437c184e3d85c1e750fbe6396d16f83c2c71c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e833200049804882c40a2909050316e0c5a4e895937b045849950627d616f5008b309eb02a8ccd3062c45074c1281cfce063e256562f4bef39ff64d1c666c189af8bc324fb717ad6b10c7a7b177a7a21f30a093;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h338922b9e0f328f46d4c59988ab7374e33be3ef19428fbe7c765723a4110f8c04714d9287fca40370f64b1b461064495a41937b2d5e728ae96bcdbdeafbd7cebd743cd1595bdaa0327430e5fd7b6cef87a74c8984;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a296079f3ff264e66687d2ca86eb35a9e0ce88bce4b580ade46de71a242b7cfc4f70989f6f5b12b86cc691458fa8d23e113a068a0f10943cddfcdc49191b62bcf04c489b8dc511d21c4b835a773078d49aac4344;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc20e58532c75275749284adc54846b62f3eaba67c6dace45e669179015f024932f6ef888665778268e3b3997dbca2ec23e5faaf82b4a2b69101b9e08bd8a03431f231d0b0a75ec41537b3affa34f320f42828e450;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h199b2a6785f1194213a7c9596e7a5904407dd2e885908940e92ece5b6991190c1240ff415bbc3cbb5d4816f507ca43ca6e393f207e62ddc20c60acf65de8771d1978cd8ff2d387ac5bd40262c9fdd5d1a5a8939d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf419a8c9aabf3b1a73edd8228af3dad239c7b85b2144df8c828bf6f46dbffcc2fab6f329d7b45285f30f4099ce21dab35fa2cec853ff16e087db9caffe3fdc137d41fcb8f170b37717a417942a7113e312064aa5e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93a5e041c303123ac8aafc2550cd45a144775856381f81e7e7f5e87f80e5d4c27517dc73e3ce33f116737fe6d62e626dcab6249f1d3f9f034934a4968f92ade2461969a87b1a1833b7076b382fe046b6447ce2925;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94954405c98ba634015024b550b9ee9b77454175a714a11ecd654369666a14fe78a687976295bdd98fea4092a4d439ea7ad049dadaf7f703f17d2ff8251025531c779761ccf9f3092aaf7345697ae774eb91b6d89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc7c04beb85f340af7d27534146e171169be0daf630b982b5726d5ba08b929b58e2b9f2810f1d83250dd2b29f0780ca9629c89c9d775120631329645b5724af320f271e25b4e43e97df5b765be20a56537e1d50a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6b383dc4c32b77fed1e4a6b1946c412194ed34a37ed030fba067ec6e02cb9e6f6c0a4556e54d21bdf93b8f9478c9aef21fc2ef521fb9569280b90b841dc4594e6cd3bcc9e841e14e6d6dd582674b5441d6853111;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11c164b6dd97067455e19dad7add8db08a4cc15ffbd6f77f9b749988006d79f6899eebc99fee009a122d81f8bf7e85371efab5c5f1cf8247542d6e3cf4ec409934cc18f0718ede897ec45437234298692e1d6f43a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d91471391c078538a57451d8c33639df9257ecc4e22fd03c5c10e03c0a7ece126564733b7dc0927aa51f6771217f6ac048dc2267fc264fefa4152ae62ff3854e27c57533e8af989170ebdf6b48f969f9268ce6e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c1a52a3fa5254da3d98a0142a0beb889d939230188ee8ae51e9ae8115e96238543be7432d0506aadecc97d958211ad5b567099a4ca6a7ad144005a4c4ea91fa4e27fea217ab0174d5b4f98819fd3dbdead141b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h756442de5baffdfb8776bf41542ef21082fdcb6507e2d112611b65075e52a8628e8a6c9999b9d82887660b40794f3a82a6220f23dd90812eb01a8f0fd6c04b733c917dc0ca93f2890d6704ad808d8350cf72e81ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e9f657e941ef4d8c1cc977f0a0c42ab368e94b6cc3b13c8a3b539c7ee4b272c137e8f16e732a8ab54b674742ae4f5cb79bfc658faa89c5ba79777819931e3e0359c2963decd0f8851ed0b8f7960953bb2cfbd82d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haad9bb49e5b939a91199fec34ad0c02f7e82f00b86ddbe5cb25332cee1ca56618e5af3fadb74101df8f24245f463ca31fd2469fbac97a9d18563d6359fb18b54e7db7a58038c8560ae39443688c6a1c713a66b323;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h195f33347b15b60bdaad462ab93feb04b3d9e3b552ecdb93b13e59313345e6c3a02af09080426cdb72b398aa102e66042e96456bda3923524e2af064ac35886974063951d0436ec6af7b9ea8f9f003ef7ae46afb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44d2ed2bb38fa8ca36ac6afa00374017130dee138d9ecd9c11d8f46cc69971832f1c1952a18035b7ee612e7b24b278e6598c3b2e9ad8987857606f2936278818333fa6567939f12ff6b504b217afd5dcae9cb1718;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8f14c1fb20f803ba8630e11ec5d42c6a42c6458922d0b72b1e65ec6b68e243cd7d6374f02bf1626baddb0d21385f5840913a38a9b4e10b9c6fa6a0738e64c72186581b7404fdcd7fe01572cd739b99f2c79a64f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h691eeb75f8b0d11ccee1615be2673a68507db7d341bca849725ff7bd516dc03d482c85c112e8539be760883b2a48a41ecd9b2d788d0997e1c7d39b35d1ee799aab4ef1614a6464b2c3e471ba736cb5283e6977a7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a75e63562288dc3164d1973709f00d89ca143cbbb26303c97319dedc487a5545a9c8bb2d11e14cd3844b49af15e1cf4dadcce4aef1fde595d38ba5096f7c47e337f0d9acb83d60f467f87b802b49dc8938b533a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd10c2773385f2c7923827ff31e5e066d4997a4c6d3efd41bf0f714e2f92b46a600eeed387d9b196c58dd53f950c8e7fc388e66bde9349f25f0b68d5abed2571d78a0e74c86c4f032bd8929f6090c0ff0ee7b0170a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35e6d52384235ac5fab8c0c6fdb0b471d9bba1dfd9a59bcf04f9bfbf3f65bc9bfa674583c0e42499b29bf64bfa6aa2f23842143d1309b57042a59db3aaf893a4e2eb4f6d5153e72693cad88562a1ebcfa61935a19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d713c97bbdf3c3e2d9964ff9a04e6bd1597621bb8dbb076d286c5120cdd8ed1d03aa9c69ce6eefefea0af622105a84ceba074833eeaf9dc5806387306ddb60ed26dec8a2fb92b9f50eccbcef425e2d2cc9719d21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb65836ff932d6c33de8452908b7d3d6e8f8051aaaf564ddf9669abf71081d90be8ec264881c5c1d4bda376199b17aaaab645974eabbaeb6197e19f89cfe7f5729d8ce524e3e11c229d75c8ef22632267d25a6943;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f8e176f256c47c07b319c22267b78ff50370235cfb9d56175e1561a46bd8ebdab5fd479a554fa5d5fd3a383d6c4a15e846fafe6f280b949b73b5032363f30e133e3ffb7e34604b3bcd6be0dad1870a7fed0aa5f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ad566b7ac3847a7e4d960b4d4d0a922f5877416452a58f5e48e7297dee7bce59aeb42b2c3eeb7c162de4e717ef902c8401942ab7039368e940be39140b90688513d4607c96e6db3a5feb374f3f8eb21ebfd13b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa42ab2be24a16920761394152487cc7e4592b07d8e3848db51ac38878e423bbfa00b5dfaa51c2fa927dc8ae4878efdcf97f57444f2d62115bbd276aec09cbcd98892584463999b77391f3426e4efacd13cb68073;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f183d12961d568538cfbc1c173a164e7f424a6135e39e560b7b326d23d0941cbb2b43d91b6ca93ac158a0698804114b86153ccf7106ce8ebc632de8d68db7e4b76a13126eca9a4cee68a0088e6b03934b5ec074e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2fa57c7d7dc60df140916fe681dad792d673929fa67ae7dd3d42cffbc3d6e0b6bce768c01786b59243716f1c8c496666aac1551e7de83d4e9c338c0d464a8036556faa051f9a3a671e6e0e2eee4b4e7dfc41da49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89940f2eaff5d440ebca9ac01b3dbc6859d82030e1e0b55417cecd897c105d1920079e3510c43d028fb933a223d1b493bac1bb3c59a289c4bac56d757a7d053c825fb16db8392d199b15c4e5479c001f49db74994;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8f0ded42a485874293928d6434fc0d27d46329ad14c3cda4f9cbdbc2cd2046cb352a673e29cc0ce5f4cf0ca5e35882d7e03b26e3626d540b68105c25d80b9e97f3538f5646adb57327cc6f98dde601e30524955d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c7dce2514f3812011f981d16e92bc6e1c532a529603d5070c4a8407c852438f2fd4e4e881a6a08784c25cf8fa247c9cc8a5e402cb84db2f2e9918c0fc8c4793ca7eb4f81ed0f985069bfb7d88608ae1ccc3fe9ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d7f678a6563d53980b8e821a57086d19a705bac6533f4bde1862258eb2d667590a43e0787625734851e91bf27cb3993f94905f0be5cab000f9ad453bb4f3d82fe939854ee54850a04921013cefaa647e091b7450;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8751e9682e0f00b7367a2f7dd1fbda48e5dbffc1b29a3d52193e506f3a05582798f551e7f80204b6873f2608e247769c53908228a0d2fac68973242fca3dd53952161b0085d735087bea60d8d7c5191647b234b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha858448f4da8f4bc6ef938c81e1ec1d83506456defe1cacc4e2979f57f5df5c60dfaae548b65ba74eebd54f44443fbe0af98f2c03a9a7cb3ee6988714aca36906f2792e73e6a7244eefe6f0cac8c47ea5ef0b7c0d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf4ac856bc3d28a7bf1fde0e8004688caf21b821a16b2206d7bfad5542a7ffb462265c312ee3a62a5ccf3af3a7ca8bce19c542717e05794f50048a2e3bfddc8dc2d71dadf49d80a6789ad593238fa1cf2371f7c9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b9e13d7ccca026ab52be50f4a2f77ae02faa915c21a689b5508e0eb79d729cc2beb02351ce78bbf4f7592cb4397d6042269d4ab0a71ab331e6440f17093d315d068e7ea1d7cded0d40d94e2127be561c937d2d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6931479a46dc4872bad735f70fd6ec9cf359a699376e09b74c1b2df335dad3cbe4797dc9e84a5fc3e85f786329227e6d439d8dcc4992113e5a9879a3d5a429ae0d28b6763aa6d714641a637bb55715ba344beb7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1760f033845f1aa1a44585bbf99d4a1ee50dbc493f377fbbdecc72caee5b824ea01ca552f067250eaa27dd837a8f7ec936ca31b680a869b9dc251dc5e2631e924bd51e1e99fb713cf1261508bebaba7836cc2ccc0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bbf32c4039245d513f9304c88fdc44087df65f70d69bd056b802ab8ec1cedbc91225fe7a42a3c1a1243b786f0229b262d3df0b6c7d1c5f4d4f36843096dc0ec1acae51d162aa76d50a56247de363ff1d4f63f539;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h879a5b9be61b7d7c0d0b8e234e4b68bd323adb1eee1178384776d61130a3dc57846698d902da04f1fb7e3fb33e938379272c3991d92f7f99e32ba2f877fe192036e652ab75e0620364b9f6b0be066d0e74367e51a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b75122751c59fcef26087c242085c360e6330498cee287f98f2f19745a79f86a547db531987e9c215e63ee25111961b1d6fcaf5147d0e9e52ec4fb8772a5064e300ee2a035bf184b9573940c203c056e2de17d9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h484cee52a8e7c4c22e2e910ae0e92a0f1be519d58e0213ace6af0e525c536ef3758de89469f355354cbfe6d444cba7e8531e45e7234894f7ccb51ded6d881e9c0de4ff7b8bde9455626855d049fe83aea820dc174;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h489f87a96b6c68ed6e92633434d0081cc6f52900619f053f8ff9e1dba3cc95406d8181c0d221038124c226c5868792e732481b97066d184714c3adf97805f03f1f2630b46f447ac9ae5e00d3c8bb8e936348032b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc45f2e827cb07cbae650cb1f64ca349b06eb333b6ba480d7ab69aaadf44f00391a0b68f7b23da207343c72f02c05cedc4f430efa34e91a789ce076a8f7690e0cfc06cf1a2520684522a46266063c9ab18568af702;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea0fbfbdc075fdd296a3bd0df33ea29cd9e92eb72c7a4c3df814c317be09711af53d251517bc44f80a5940da1c8c5fa58219c1afe19fe15a27953c872d4db1a4d53195f3bd418156132bc85c8d5d9e9e7fcf9cb95;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c4fb6c5075a3e813fad32252186580c4ba0656f77dc103e3bfc97f19e81861b26fd53dc9908143c43ef3950492933956155617b28506c40d70ac8658a0a06270dab2e284549dceff625246ec840bd7e85dbf603;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b1697d0e20d014fdd402528a90931583b6e2ac048d2e93b739495823e709c2608c7a5743536b92342cbbeceab44cf1609506a1dd202875a4e85e67bb0c2c52a7be46555b4fd97802b4995867580841c5986e0470;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h151ea4a415b785ff086b1ecd97f0601d04d2115fcc61810334add9fcdb493445078e2443e8df955b069feb6485294673034d154b6fdacb3e99c954aa6bc0ee5ec7d003f55c15e2fd2fc83468287490a256e7a3788;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h368d907e6de36c20df66e07644036a37087c283128fdc0dd3ff63de78dbd238ad69af6585028fc4747ebf6ab4da9ff81323ea75f212d178a54537b90873f8cb291adecc65731337bf89b0544d0fc358a33700d3d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he79a34e07b3b2cc4c7a1b0ba21406ee4685d9e83a8061e749d1d81c9285e46f2ea75d9df98d6e15ee197ddb39016c40d08015c4f2d5aa2deccc44abb6257eb3f680875448c5f113476a33a884f0260e4bb9446942;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa4e6bd592312237700102698a7851e7172fe0a1b6bd70e497c5bb66f23a346e86eab471bf0f1ace8c9c2cb15f9e5c5f1836fc1e8d48300b30051bdcbca16605331f8f0564a75a48d28615e6a7916d36309250ad0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha39556079e87b1d16af538715e2be6c2ada95271da8fd8161e9a45b0c6ea0885c1287f21c6b81a15a97d71fd78a05c441e6585fb161ef320b2b89f9dca5172ec5b34bb428a21c621980aac3c97689a845e5b2e769;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83cdb361acedb041b6317aa8fa565a443714348baa5b1fb940633ff3e54bcd4cb41aa9462cfba7d7b38732d116ff050363939129d72f98ff355ccb33be75b6a9513c3c3107ec7462d9c8185ac699c647b6287faa8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h413352ffbc600363ec3db4b542e8a455c1f53b44c87b535d0c7bf14a84479e29e839c1210a0b3bc7752ddae4539679edf0f38e730b82c3e337cc87527c38fde643af42f4789694399c84c411defb0f3f49c87ee18;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87769d25ad2a4881ece57fb57bdffe055a2acf0626a6b4add7ebd2782b047b7133d4c524c56c7fd7117b9a67d2af0d00cffb35e9348219325632c8e706dae41bb8dd5a5f8429b3ed42168248b67db22605ec7929b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a4a533e9d6a88cc9fb3661ea17bb641af6e15dc16b2d19ebc73741eab262a4530e95f760ca5df18702a3637de6768bfa2ffedc96ae2e63755c498ca8bd039477b6ff255a74689a8a3f90762d357b2213a8d47ee5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba6312acd13e2943a1bbe287c9202a18b4a5486eed95124512ee107ab76b5310d3d23bc930e044e558efa3db59e196e58fc5598f59ae9d2fd33db7825c0b8fae8fa3446f33904b87dfa978205ae094513dd4a25a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67a6d85c499157cdf6ebf9e794ac728ed239dc946382e8fafc06523952a168f14813c74ec994d23ae3ab2e415f9ec6031aba246bb9477a19d1c9b744a6cfc861d3e65a59d65c08862a68b6cca3bc8f073a2fe7df3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h267a3e20ed6d46eadcb09841afb1770b5f67ec7245c7a5553fec87259cd6b765744995cedcf64b8d058245f73ca9fa5865e990bb368f4f2fd539010909c6e6e5ff77293181606af4e457aaf82f1fe6f1f97c358b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd8ea64614f3104ef97e8f3667a57400fbfbae7c7763f6c9bc5a7d9f48ff403c5e241571c6f68272fef558247052e010af1924751c63cc4b3c0a4385da75e4de91c0413f065beaebb71209c13e1fd870d5ae5724c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c499dfef66bf0725b8256115464d99bf11d5fc88813e095784a070b4837678a4e8d10c678f13ee4ba79d97fd98bd9aa0f5bf3333ea6dd4c076941b299d478843653b795e2ec2111dad786c4a22aa3a856c4316d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a3acb80a1809abd474658d95e213c4d6d6b1e95dfb96095fa0b93a71f4e9e023e471debe435f36f33302d744b2a3d5bf1e845a61e34c71a80a73ed5e63504ba206e5b91898221b112d58f21e1a328412cc2521ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22aa41733cb25c962aa31136b4ce827448aa9177d0d776633d0512bbd61521171a3a3074040a9c063da3cacac2b436cb07506482f343370298d72c76862d7c225dcb3db2892c86736ba7bb10ce8b24d39ecadc888;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefa2548167ea1b020474bf0a996acfdd57f43cccf5dff61e8c3bfe35b620689e9350beb2d52c41fd557080ac67bed5aeb5cae642439e80911c7dc3413a893180708eaa57d0240d9bb2713b9234c0d5ea4c3b883f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ec34ab24e0b2e3e27dcfc87e0761ae0f1aa483aafaf52bbdcd2fc122af3b0cf02064e0547087c9631e8d8b5f70dab24482dd331e2e33b5f1e9eebd279642a3990707df09abd43984b5e9da7a7adf117beaa9d2af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71095f2e9d24c9d06977e91356bbcf9c843d19f8534f125dd6dc2555b209a49f544fe11c287fa29201763f94faf4ac9e800fe5ace3f511239c7bcc120436fac1602302c8d4d375ef28d0ed860522a99024e7b1c7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d6bcbd0526d37566e8c2aa35b5f053097d7098b673fc53961999787cc3186d777131b2713a5548e8cfca9b7c32abb7dfdf0956e5c5bbe879e9cdbe19e27913673545638c9fad5841d03565d613f062d7574dee48;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef50f83bd70cff0c5d3b5ca0b0d2abb062fb84c5fb893a73b3229b6eba0126a5b03c9a531fa098c37638f3efac3096a8c65aea3e21544658898eff1611d5aa453ec0809a3468e5d87165ac15902cf4bc7026ed667;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb0218af84598cae38a761ecffbdbbb2daa67d1969ac28b27f8d246030cbbff8c7296059552eeaffdd6a7302a67f45f58e47a9506dc9c7564e312c7a6bf4599c16c98c982866ce2a23c85966c4a77f7cfd85ac42;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a27b08928a19f332f056a6ff4f7d409a7b35f4176660f110955dec6fcbecf08f87e5f62f330a3fe19378ed77afa75dd40f8ca46cc134e4dbe6f18d6d508324466628f31e50cc5466c42d3157d91c95716a0e550b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d2eb3daef16a794504d037882c26472dd061ef9e26567b465943d6b85d28e7349307bf63a691da4b458d4901d350dce2454144d4de0bd2710c2305e2d20e3a47437aab298e86c942ec890de7f511ea8b56eab1d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dddb271f0bc2cc36b5770e42400b52bd57126e306762eab0099b07a390f17a5e84091fc6c4ae4d6b1328a2303e28259002949be04429f6139588e810dedc027deafd621ce592ef32a6174f43c7043a57e36abe23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4e34efff2569c916919683cce885bbebe0760b55a28550c1ab2302c86dab52ea904eda369b22c2de29f99c31ba0146fe89382d50fce493073e70914cd08409ae3fcfc4973ab428013d2dcf10158f13244dbf26f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff44807a6e206cd8caca0f6e07c863adba46e2f1c4dea70668f45aabc0af3c22dd5c59805e75d02b01eae77824d86c9d1d195e6cb10f51573caca4108c7ffdb244a66ce2d6230bc08b55490a54fe02bc402796975;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he13ff864f7601d5584fc5c8a79b9e39ed7a6073ef64fc78910077c1c4ee6abf29109ac5a68393b5bbc4e2778ccf6cae58640fc23a40a01c708205047cdad8a2e100efc100a0e6a13bef36d3d63acfbdd2ed966df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecd527d82b1fa0d0497c70503633025fdf855674eee952deea185b40d1f5fb157bcd27e6658796cdebe4728db6157bf207be62f3552547b6e9ee94e1cf6cf5eea833d058cda34104ba188b6b023501c797cab5387;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2658d7969f171a2df795f49a151ca0e142065de9a1d91bebc1e09f09f7d5bd54ff863d831a545f405c5c4b4740ff017573fc5b021784506df1b99328728b4a4cb08807b22f536922fecb5dd64c956c5ee68ff8295;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72c33119ed2fd256f9863de8828bbd005fd1ecd6a29fa6a12c72f987035f0774e25ba748dbaaf4f11f720efc3d78f7746732206936b66ce28bb7d200da6ecee9b190c3de25157eced5d05e1fa694b0215ddb64d7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6429928078864e192c0fb714cc09892ab4858b60954e1c3a37eee27ed45214ca7c30c0d4264fa6d5fcb8d204931baed94673be176615eca5f16cdfa4bd0d2125b6570d2151fbe081716d0150243115275f9be3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f3e6304f7073b0f7a3eee70f782804deb13405129ce8a5ff2efecb789099625041e3763cde75285a51b26c6e789419a3bf79338d26613e1b20f09c51449434bea727cd4e61c7a74ccaa6da494627793f50b8fb02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b4cb22a8a1a65a2fbd1e906cefe7931c301c55256f12ca6db5308cc25e314a3f1eb7775459934c596ab2a569fe9d810b2114f0a6fa29eaee66d0a7a3138d693135f06a00cc138c90f578ce5fc756d659d1360591;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ec635eeae0fa1a580f3bd984edeb63861a16c3149f7b0a41003211871c6cf798aa2c4c53791f2c823c4f32667fc29a266d12d9f0bd760da10a452ed2b95fc6ecb8954651248c076d6fb6db2430cc06302b6973cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e2e8ad2cd70f47b3f82011a69eb4a1f34a01b868c35b041754fabd737cfb8ba1b83a0e1a2a00354dbc5d5965515fa5313ff74f545eb66eb8ea21c561942e7f9cc0f551e1774aa5d0033428d2985fa3eebaf82850;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2521c6c1fdc384df4f3114ddab7c95c9f9bd2097aa20be49dacb0d7e1d92af09d61060f287eb43161191cb195934254dff3b7439b039405f1cfb755c93661ed0e31688630b018602a99e43a536418ba66a2d4147;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800c5ef34fb54c6fa13b7bf32ec1c6f918b55664442f61ee9fd219249e91bb54a2c14af2dd934828080a48a7e24bd74e1c5c445dcc61d996f95fdc3450c51c7191d9e8b476f87aa7154b0acadf0a98f32c1d9ef39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a1d0107867eecc532f82f1eaacb9f5139a4ae1a531953f4473f066a1c5aee1c0203953bef58a5a2537150aa9d71d4ce4d68f68082ffb50568ffe5e4183cd680aafedd783ec88546a729fde914be8fa488d4d209b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0e32d1f3511119f2fd73ea3c8b5e6e8a46abe1cc8d80643a28886a5e2568f9c35025d292287cd1a34c18795a32a471c057bb7c07188afcf0c60dcf536c39d51e38d63b3cb04ba56791f076c215f80556d75a1c9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f04b7b5973249ef4e0b6a07353590e93c2e3590eaf0599ead83fb2249957f749ee92ab58760058e90c53835b1fdc5c6ca39fc4043261255b6ade89a8bec518570f5a08c9ae211152362cda6a84d3342f0750cefb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1594dbce8d36ad09b538855bdc6cea60222a9202b6a3f95570f06447786fc6dd452392378d59544b564205e5b41f46059b2981fe81a5a0fe1fd5fc89503dcda43f9b8ecea22fd5cf1cfc72ff3149bce38bcf5ea45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ad80fd7fd866958cb1115b1dd61f1bc10a7aa777da499b4ff33cc11e7d5e3f1a8f11445173dc548efb67c5837d5f65f41f05c15a3d78a3b853541425eb644a5c6232a473047230566e9426cfcbe7bad232a499af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd611e95f141dfca2201dd96d587790540a62d9c1ca654baec3bcf0c413a2186d56bcb52f4bff71bb94a95fbc40eb4ed4efcf2e0fdb0f678d76e539acc26e228337d44a5929b77972d43deaa93e28d50e9f4ed482;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacfccbb6f1c6c34cc0bb16addfeed70daf895d5f8d2ad3f7e04f9b27d2639a0230b0179ea02a8a8fb34983deb0e062c0b58a2277c13b451e6d370c0e26e133309e29d558764fea1d535341b61f1bff8e9a4a3019e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h114cef993492562a0d73a5a5e4de8bd9376680d2d5c13b836e611e5aa03f8db79008339ca62e5e4c6b90f4d73b8a09667fec994f9399652bacee68e1757803225632f705bd800531a9983cd93a49576d8dd5c7e2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h733d477b22fdea37ff9d58f46d345de55345cd49b96812fe4e36bf656cf17de150de56b031474d0e275eea3b41198511977f8cab60ce61a9103658606496dda16a2e1608d03a3966268cf5a479fc22e66e122883d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21c6378558d64df93304611ab22ebfffd406cbfea271685aa5be49d9cdf2b6e4c9f5d182f8fcde1f3b7337cfe8821dd494d4defd6f4ac274fd6e30db61e11281446a0f0504d2a2f2898951acf74a2065f3ea9c893;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h572ac3ce2eb60464406eb05e0b7941bd33e78b1e3e457ceba6a48883f6cbad1f9423d004bd11e83b813d85c20437592630b409a1964141357b4c71dbae3979d9b78f62be73d67572411a12cca61f27df711aaac98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f0cf4ef1eac5e4d63d4b26baf18baa35d0f0ca874b31807af21529b3abe65c3f0a35130941d40221410519e84216ffa905fe83df7afce668d33cac86412785d3dd130647fc15fff8bc96a21a975dc05119e82936;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7fbc39836e1340cce105f41f07253d2606e4b09d4bf58d920483b4ba0c020ebea61b74d8e0abed14241bf1629deee98e1bef7a2ba9f3f1fc6c111dddf7d4c627ea7e965e8d94093ddff69f5b183e09ce6073d618;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0d14750242506c2a1d39417ed2a8a199c172784d7b05b18ec2388bbba8fb74245326c0bf663be560104f8d50ad46d845e60e4a07713e06370bda91e2103ca6d580cbcada53cb25e7eb31029940b588e85e00ae28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36d0552a9435d47ce852299bef2f37857b5adc97a1071f9abd594fa771abeffd36f24b77013d4e3f3d794bfd75f51ff6499b56a800260840a27c89996431f61d67cfa9a036adda2d5560c5a209807312d85f5398e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1318f5e51e6366b673ac0591083c70a421e907b20af1678bff05311e02796470ba594702bad24b64f159778c8290ed5b4e8959119c613b0337d145ab95f3a50a9461d47f9656bdfc9dd4a668b87e7497ccc1acac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h327f64f563f8a4cd0e986debe13a4e01026b5b9415ecd12081bc34b361b5cd2b55e64051254bae35cbc8eadebed1f8d0a23832a979119e1d1852231b7dffd1713aef6be412205cff6bfdcf37b9d946a4786dac15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64ae71bcb6cb3f7ecd559514a1749c922c7f9c0cc865560bd16eec0e9635d172121627fa9b5ca9968f9284eaff89c48eb7612c2a1d0fa055a6f77fb0ce8c6995f3fabeff9f72745e2712fb004aff5f84f9a1015f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2aebddea04d668d927728ca632090fb2c17b39b1f4c6dc047339274f87cb264c1cdff42cac725039f63f2e9bf99a1e17c1d687ea4237d5a783aa143b197ebca281036a158aab1ca7e4c5b7298d9a604d2fb24cf6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35044ce89752a260c167298acb43aa6ad5e39f525857171dc255918f60072436f62cbccefd9db556ce683c04635155c941c5a6422189aaa0711a322ba5a131041a52a92de97c77e3748eb6ec642316261cfa91532;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf41f11f33ad7e88f265def8b4513b45c90bed42f15959e08bee2dfc68c4703cf607ed4331faf1dfad90d94a4b6551ebcd5459acc8899f47d85cdf35ba92f7f22c5e6d434a2482cff717b9da8cf40e9c5f9ca8af09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e53797fd128ef97fb4210a599c1f7b5983047ba794bed0ac2c1b01463b75a628bb97f7acd12e68da044974cdf69e4307f42b9982a4a75ddf0b2fa1145af74bb4ae638b4df9f0832184af45679765ff06ba1ce40d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a4b07e825242e905ebbb7fff70f48ab675cf48210a6bf650204f39d7693a3ca72cfdc51e94071c4d7abe7854ea90871feb58e606b0d62e087034e9cf188ab5c7311a11e6a4b53fa13f464b56091ac0ae1273a31c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70342d7ddea7f3843c8424961eb03dda69451e9e9577417112cd0d6f9aafb735fef2f8d8b03507b6e065e05376d7ae17df506f5b77fac0b26e6897a5039509bf591fa07bee1c7955a052e29e4c866cec6f101bcab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb182d31210356f927d7254456925ebb8216a121933a033bb638f2e266fbb53871ab6f0282edc4f244eb510eb56c0aa8361584d248fbbda9c7e4e7dca86473670f1e774fd8ca457e7757e87a0789b75aa4fa58ea0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c952d87cfdd066b02ce8f74b94dacfbb590a20c3a655b6d1c795b4228785702ee61801e5c75e2970028fbf7b4dfbdc26d702622044050fde5006c007cdc3c1eaa7b96bba791d1cf98150b82e72da7591e915cd9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ac5db0af0ae173912f1dcdada01be595b98d36597ff3084b986b7971914d87f0119c4583ef6a3ed9de7610435a83c88e57179e2f7e2abe6ebea6b27c5f674a41e546ec293ad16d43189ac253b10bbdcb2c759ce9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55573549e39f10ead8867b52359cef3937298bb0dd92cead9424f503cf1b2adbef27b83dcf31e643233b9ae9197a22da41f33ad95e6caf5fc79a49e74312cbeba781145e5e09229ce240f9ccebb3801f94d4f49f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf9cacc193f64a8d5f3c0128fbe628729603ba62ba8fa9768f8d9cfd753bd7505c4ef46a9d3b7537669419207e60bec272135b212f6c479912233e1456ae69b28a3c1cc75ca3260a2241d1779bd4b0c7485dc4f6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3f64460e2b8092b4b8b5fd8e4e1325ea85f23af8381480ffaa0fd5c78ad679d33e3b577f81faddb76663c582479c27744c95522d531bec7aa6b4ab5a3e096f63dcc65440e2b3deca51570d3c4c379a351e67f6d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fe33e2805da36669e7f99affe359438646d6dd4f4d25f3601e2e2c7b76721d56b99b876a001b3185771e4011301dece11d541402457403af2afb67874c07c575d9d54b59e84fd5db322e29def8e2afc7c0ace6c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc826d8e552e49b076102aa942550d39a043da9acc5454262cd2e0cb1a1fe8f3e70cf082e9a03a3bb6b42099588a620b781cf1cf4f7d5c7e27e89ad766f47b5743d50a823f2ffd064126e0601dc976e8719ea4180;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c0b9dea442c80b24dc7a94dec13294b7feea674fe6b506af8ee9617917d98c5df220041abd671f3f8e05085d2399c24c920e9263b10b18361c9ce4d71a88464ce768e33b020d32b0c3fa740c9c38315e5069d4fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2bcfc3039bfa1316d0a5faebbcd84886c5f8c6c8864615cb2a554ad5dba9dffc7c69d2e3b6f640f21e1716eaa6e8afc9ae0f42d35ee0849793822ecdc7ed18e9fb55c528b80d300a1f0cbcf939ab0877c83ab6fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6886b981448b585db0c4fe9310f49aba7f0ca4937ece9553bd1132495002189e7925837fa1665f3b1183f5b37bd74bf3d9d1b833a688b80085eeb9f76b16bfd6764ffbeb72d0eb7bb3f7489e8c4287f15bd59a4f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40f6c9fa990719e83e416082450fedc92487794c59157c377bbfc48ba9c29315d4f0c5efbebe6c53008f5f54037240873298eb27f2ca55a7a2366e1111b6ddf0c31eef703dd4074ca0b87625a0c23b2a1e6f7ddec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd74c713ed741c420cdd68c53bf0c2c093ac8166c0774420a0b04affdf93f59de3c5b9dbef3fcf94499e2619b33ac7b1a723ed19246dac4f84aa4409809be60b36e2ae7311932bfc8289fb7f5095ae6c79fafccb9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9992924c5fd34f10b6f09690ebd3b028213e59461c62ac993bdb071d23b1d4ea3fa42ed5120a5db4bda191ff721a69a52ce6e095baf86d2b5fd88527b581067788606d55f8b8b133d7177ce212a66c0c313b6be5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3a627e14427e0cfc5c2322fd78d49e056dd26272afb01bb530f177aee366b0aaa5a5b44aa8a944e116614e3ddd342302f609a3c8c0f75f773ba8ebdd9bdf45b491843d4695b11a7a1e2cadd33b1ed54bfc226271;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1af0820a9529f86d668c112f41dbdd4b062b0be84bc637febea489498e87aa23bf70535d70680dc932980696dae510cd9d4d089c7d38016b40daab6405e3a7de1e0feeea8800f9875522eb60ef0c6522106312544;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7c2ed1cd11cb20347bce9d862901795d670ff55a7431ead56bb1b9d19bb9329fdc335829aae8adbbe2708c5986959bc7d2ea8cb90157cf284d3c68ab45b8a3c16d04bded21633be53088ce179b24faf6fee54e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h484298a990f5731b8bac33b6f99511513710df98a7e051e480de561b1e866e60da2f795ecfb5109887918c3fd53e79b6cb1b733b08f3321c8527e6cd86e1c63c7d3f2f733a6cdeabf2b81ce8457d70ad94007e505;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed1730498417c151b15a38e16df8093d94d911fb18a2680877df8a3db1901868c50331da0d43c2e9e71680732add0a71c6eeb08a4e62c13367363752895c4977ea4a8a1eb17a25c458805ef77f96c6b36ab31a13c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93bb131e9904c3ade0b75c40cd10c291ed14f5cf1ec729fca5fb76e36aec30bb6a084cbfba657fabb2e6c300dc0a090e47c38aaa930131418060c51231a0a5a905a30c2bc9425b706c26b76dfd5b36834ad5c99a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92b539e62bf1bc1719e20c16205f1c0645d36a84edfd08e05112fea0ca64353a718d6b69043eb063ee0a21f0aaab63e10015eb9348284230f01b6f2eb13be3c9151a71de92585312f76498224547affd722de35e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb21d35d51dad35502b4bf2588e12e4260de7b10a5d2616f00c1ddcca13063bce0ae9692ebe7e14c5a4d34e9fe819bcdcfdaa71819b9bb007f3161e4708c345d0b9d697c8578fecb445787acb3a4f3c0c64758ecb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c87470be01c94fe8fd28744cbd179b5d940644bc226cb849407931ce8536c1dba186560b5eb870d672e8ff6642e066cefc3576e1f97f7b06eba3a96b9c221a389cfed6c57850c2966f39360c58cf8ee954e98875;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h791401825e50c9920640281df621682152e2746a57759314e78434db5ac7bf92ab85c5094b7d34cd2fef79681639166b22691e85b79d9d21d8cf454dead60bef8dfc1d6d6865a0fa3ed847f13ddcd95963e2d3e11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1a79b591fd5949227acb3b94c8a41b44fd8e9b64c6cfa28faba60cdf2e5e9b5559b0f88a171a41d822fa48f3ce0878f1f9cd82e6a24c14e4429e933ba9390427d947d2bde32d058399baf371e9390ffb882c120b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3cecc6a61bb840a04a0f1f4601269516e84f598e61afde8a3177c84553c43ad91fb207664a2beaba969c540378e127fb59b7b63c86a02407b94dc123d8f066eb5248be3bcc231615e8abbd6e507e0465e9e4a385;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h134e40768c1869d64f25b1cfc89172b4e7455e1f277f748de3ca5ce9f0d964d893f529768e6bd523aa476ef1e7395907e132f29605aaf072aafff595f0a7ecdeaa4ecb2450a0d7d04fffd3355d05edcd081ad3b1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf351009722c0c3423803acd72f28aa94ce8e13e72df6334908b0bf742f10c713301cffe5c29f4c0ac80667ff63fa1ee1352f7c6bd4495c189e39942cd708d1c371cd7d6b6f7ff02cf1dc3598314ddca473575f5c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f9500abc248fae124591deab543c0ca954fe20310d8c96ff308edb970f15977e28d33f67588f93d264527c361838ef4452f5cf19d943000cc9b24409cb8d38e1e9ba134339307ab9744c7e9f01d6ad23bc8b6f72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cd2a2379e095e4b625520da924944f160991eb413a58075fd9b071d18d401ea66d331bd2943e370153c16a1e079aab658dcd6d90a2da10271ddd8ec80d684739c93e4d42a9fbd20957a1f325e9fbf4bd7dedb3b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d8809375a517f92657fdc9edec54f4e5019b71b98732f474bdcbaa7d15bf001b7273fc28f9d9e3c261097a5fc312f8ccef805fff61708f7636a0efabe16d514eb8755d28989026051f8c6dd0595b43c91ec5bd19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c33267fa7788989db021e0691b862475915ffa84c47b3da8eeda957b2195b4b3a05ea97d5fe319bc02fa8a344400d44c49bdbf1f64f72a308d5c3926c26a673732b4ccf2fe2e9892e4243f8ffff04b8f7779df92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h136840a36489792c28e06e552abce5ac8e97d79166e37cc3b8c4d7588ac2ec0cc8619d626a39cf59e0bf04e270ee83c060dab94bc51750b0862a40b9a4519c7b96b73776f18dc45e762297bd0ecd3f1e4f371a87f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2726e39069ce6b3e02435d3a8cbc9f6b053a82c070b3efe88526140b432cf3ff62e5b451a0124ceddfd0b0320eb4c59148841c948b8fa87267c7365aea0b04399a10b3c99b6eeafb4649b1e7dafd4c8d62c009694;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2634217b33a5df60d4c7166ff32479bb5f83762c92c2f37e997ad44f0a026c739a25b303e23db1e326c88d555d866bd7fef120d5c77bcc0caa95c340099169ada945ab916114daeb033eb0647da15f4a8f6a8d6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he07e4f8bd1b2303f976a7a98f5c63c68343f6d2af45774d15a95ba4453cd198cff0edbf60aad50e2a9130dbbbc0c841a64757008254d99c519a8b0cfb93377326aad6d739aea83e5d52d38685984ce6df7be78118;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22aa79ad761e3febf1ace609e385e7495c7220ac0f4c04b2f61f3781ec58345afb4857ab14fc2ff7f6d9e81034e77ba7450434dc2ac3d922aaf154ec1904e94fed94d9cfe46ee4366c0d563649136c5df08950e2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe90e483c485d3ca67eee59700d7677580b958a6878c34468c8de71e7db919987e9630d8c257bb31a46bff6531f1b85b5f05bbe914ca4f6d3dfce2bcf4647f32125b7d554761493271af36b30eb68916b22d20412;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0439db9a4645d9b0ac33da2fc924e70c10e844647bbe24065f6c03322f31ae87f7b9c9c1d47d34f6faf9927d8db77e8eb9abf9c1ec84868691fc7bed97615a9a73abf3ce5425634abeedf0f65c1517e14fca4ea5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h164784eedd2905fba3823dafb3fd328e775cf70b8b09cb97270cb721feb7af3a13e606c09051404a1e35dfe71cdac69d22a62cce2ede8374f24e188f3f459051b1dd8614620de3d74bd5df00bd14b393eff69258d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d2aa738b6ce0edccd6feeead755e72357a198b86ab407078aad3186e5b724eeb804eea7391a77b510e0c7bc67cf5e606b03d431bbf45b1806a65275a1271942df7839d1a6ff436f9706d349f5022d34efb97b8fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13fd231b31da5f87418ea6a4e3aa7d642f1d034b05ebadb68ecb115a1b80b74a8239c6172da83b28cf186bdb94683d8ed5efab270dc2e895eb5a74126df5c9c985a991d31b7b1485064f4d168cf7287ef2410852a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc08e36881d724d64eae3ce2c37a4dc7369e6499b45ea14526b4c25c95a742dd8405417e0e365cb70515047cd604ce29feebc2bec15a931fd86e501dc624734539900c502961803b44c53281a9d537dfb581fd6e98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h656529b205d29c6a700afc37d02746717c1958ebacd9a752f4cc0499d820b7f32ad4c266bd5a09d9b45e0cd590bd5fbcaec68a773fcd23b851950943bd1b6d7c42962934b5ffd4d26cbbfba7f32a02d1fc22be911;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37eff7c69930c3e85c3b6afbc1c9704be094eaedc1e4d81a3ab37cc0ddb33be658e720c166bed88094e8042d97aea9131ae11284bc91bdb396bef91edb3e3543abf89136a4272dc54491145216ea7cd3c6c16b597;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e792189458cfa026468de6f2c2162f5da08a920c6fb6d53decf5da4cf289adce7c41bf2999fd1a27973e8a7b63ef56b07e90578a4b882f366f1413a947b961e79b9017ab3b5f7e4490d550b793b5fa8b93459e20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf68224abe310569848f7b5981a82b67f728876b716c564f8933e49795ec63aa6273ad1dff2440a3ea2c16097b63a0b5817b57bf06384b6bb456071ce24955d9f7ff063eeb7ebe7d9a91e72812a224fcc0000a8c2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e29e3a3c69560af37078e5cbbc06f8aaf69c5cc65acec281cb437382d44c25d5c41668335d24b3e9a00f60081971436264faa8feafb7ec13d50befb473c5e1d63b0797c2764fdfbd90a7464469fbfbae6f16a8df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0c58adcc3ad74514bd40955f5e66f9151a015828eaf7cdf616e02eaa75c93f0dfa672b8fa1254b436ebf149e0bf76f4065d03ce20144ce128185af4a621617aa3b704e981f163cfb4c3b8f11fefddc0996457925;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2319145befcf12b9bc1046057966f967faca18c44519d2f3b8dd16c93b7cb3e8e86a4f2ea25ef4777c6c71c69a73241ba29c97a06e5c926d1e5feceebba7de62066a311f6cc7887e11f5774829f2b48f127db1cad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccd439ddadab2478c1bd94eeba4f59eb29588e48f1124c7681dbd8acbab1ce7b23f36acfe493f8105423890ea7d6c018dee754550b83b46ae06fad5388ced3d6364377aafb0c30626b42eac421a7ca32be185a648;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6713e21461e1e19960df4abad907f9f823e113e194a6598cb81fc9424059f8c3b31f95a1b3713a9edbe9246e530bd00d5c4d0e0b63f6fdeabffee6550b2ab3a06494f2949517bd40bb282d3b1d52669472695261f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd731feae3c3d4530247c0aac23fc74cadbcd4fa821f73a4b53873538c866dfc37ff80d5ea686c20ab6143afa10521079308dbbbd25da10b359b90c63fec8534b60348a548d7deedd61a21cb5cb0cc4a7627cbe482;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28ad923f560a51bdbce1b0e77e6d77302a413c387cc2fe732274f9f60c35da13d944553465e589e65d174742a81b71b8a8e5a59947ff9ec756b53a5c013a5bb2b8b0eb05bbef33cac2b2dfce70e7fed1b106844af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcb457f86aef301fe719a49083ff8b2156dd080b6a278d3e7175c06e1204261ddb275cce785ece729f93eab248b6ca6c4dcae5509874a8db6eb630e2fc3dfdbdf1ff8825b043ce5d83d72d5a13caa71cac34313e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2df783f57f69fcf0119fb69418252a870ef57a2c9c874c0f8d7cf8ee930fed17314e1e2baeffb15a61d11cd86b44856202c6321cfc861877c9a61415ab13d6386f436cf0c36720cd724be52b1f2f2b469c06877e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd28044b8cd1773a0451d255ad60602daedc7f9b532b287bf45782f128c197571d8ba1a6d80a830265896675cc654548e86625291e3cd3c7ea4e7af413839be64569e39ea7861ea26d7a6184f97555cce36efbc60f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8aae1bec18d58828804ada7b5772d5f34258f527208804abc15e64e51fee3d8dce892fbb2739fd96d8caaed0d1dfe2e4b0f7d6d019038eb0adaafcd3402524ea357b57ddd0add03cab0a272f8cf040da1415d5aba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had42ed68008121edd0ff36bfa1b9163773c5303b81a502f8383630bbf25a40cf8e6726c8e6a0ae1c5ce2ebb66cdad49c78615e9c9b32cc18c4ad31ad53a909f0857b85f6ee66b72157dbfa3a1f7f1f0a7c41a87a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3d6b8f8aa32f0a156f5912e46d235286ed5ddb00665f3c74fd631e13f9990101d5793f0c607007e09f98cfb623a181367e77c127bafcc11474dd65b973e407980e014fd7ff62565264e50d57e414db7cfb2ad58d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3627f5f29169387c1a1c4af9c8369dbccbc6f4420f2a993611b1c3e22d7df7d7839486c08ffe1a74b8f0a32baa786aa2139c59fd48e7f033091520239482a63a80d3d387e9d1befc6d7db883856ce4c270c48908;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h480882c6a75c9d37b92d22c0b54be179175195ce8d99c7f14ea5f0dc1157e727e4687726da76de7ad8c997027a6e61bf10979d333bb04d5c9d133f11d49af566ba02d07819af14ecf1ab3100fecae0ade7924dca7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8427c5b6486d58363e81fc8dfb562e31f2c1c466ebf71749317aa17b6a7900e019f20e0c134d5132e1e9184d7100bddbb47c3d2933556ecc73232b8b06953755f4af7454a2abdf8b37a2f000cc1ec15815624493f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde614df16ea3f3731e2fb5b32b6e8d4382127dd8f251b17eb01b6087813dde1a2083ba5a654bc39f99333b7471ec4950a7e5ffaaae9648ed9fe0daa8fe3a84b12ebca7d09ef54b0b568d0d6d90f8273457ec99192;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b49c334d90e8c08ead0193daf82214db74f4d84be965597e28435a4648234e895fd83171de44bddd6fc419e7fe6d427a35098d0aefb7e7b5db7ab0e89c47630549d6e571f57ab64b9f8bc5ef54f6c49a79de4b0c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3636b9b01ec7355e519ef3e614c40420dfcb6f96b066171669794e206226de7bb2dd77b7d9225efefea007517b29ab5ea9816ec4e3ef96d3899e934494e20fc20a693008ce5fb9f6bca484447893f7271a1585b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c8eeff418602d6e2f7cd6ee00ecb86120bd077fa773b4216024fcbd6de58c048119b859f535f8d6d7b037932ef6225553056c90e4ef5d268d6c3542396fc53904fcce1512a215006974cb7c2b541261acfa29986;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdec664299c78ca9c34ede2356f55391e4a4891a012e5fdd6c326082c218d05b2fc79f5d99d168a100db728a3cc0023fa6a3c33047d116245fceb1ae332836806717cfffd723c4e456d78a16afd2290c4c10346a60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71760969f88d5721ee6a5c4229c713b163b4df80c3f27fd7293b8d36ef27fdab815fad85d926182a69e1ea78b5962de946a1b153afa44c9aa68e404db019dab29ba98e9de219ad0636c427683b9298c707aad158;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75fdc32495faad4ea65fa3319602b19fa3f12aa21d41894d0d9cb76145fa7b615b7157e87c8d52bf24d23ea22b8acab62b7c11e67cd7f5b092c6529d73fdb35b609b53f4cd557c0eb097492871156cbb02d11e553;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha71fec5491b3d99f03126b2e9282ef94830ff5c2870ad923bc581ebeb79787e0bbadca5b884660b6672088e38da0d65660257342a8867a1a986ef975f9f0fea794c76e235c211a229c206987dc87cc6a4bc05f77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h883d5cc0114b7ad411a2694fcce332c6130c260ab7bfea336978495f5d77c2963e3c7d384a052671564108ad054240512b3ddfe5b1d40aa7832258194cf8bd5da796c433d9fcdda169ae69777be1ab7abdb0ece34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81f62e9bd7233d058f40bf061c35380fc6f50287a77fb4228c7e60721268482b471520c534d055260f0c2c0036029a2841872d9b2e5941b5eed7e75b04ba0fce36751d550c1359f261bb684a515b8e0d061496860;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca91c48fa71afe354761b0bf098b04f2df7784361b215b4993f984907b7e173066105b0c608eb7417412d8c89a632428e64df70db8f6412c944b960b6f99cf53f84b953ed30d12c1033758f48e8fda71978b69540;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4af6b8a730712f55ca9f205f8a6550e9a21689b248d5894af56478798f7843c57448ee6b8b1e2653770a5a3fb246a72317a70eb23dd5b292d365b6508378e7a03309496ea4e9835442ffee501ac932b459f0126b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b8f8f0391f0e8483e945749a9a9d911e8cd4ffe6db8f52d248c789ac547a5a96c1aad5b800e65049ea2432c958839d92c8412f8cd08c66020429c0204a72654f3e7a8b69af0cb1a5ffc12c0862f0f86909c23eb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfab512b64703b37d11dab1ebf93892b61dbcc676973754ea2a8ed4a600c5781ed07373ccbcf74128ce177b8bcbe56d1ea12fe8c0a573529cc787594205190c7a6b85bc879c56e38ba15c8b83d9b5b4afb127fa407;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9791b732002a88104ad9dcdf1d4af7c794bae190a0a10cbbec5b02c42f0ec3a5a30d74287ff1e60a83cf1215b8b12e67289015fcbeb3f4e9e029b3203431acd37f2875ba8d40412f7ed8fd28756cf0337b716340e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b1eca6d5d9971403c2769eba5013ada38efa582d8bc4b4e180b42c6b0ed2a07168f98851791d8680128df2a0a1b2693a18021328f916456078e17a48b23f7e0a6dbd24f14a84c70d35f143637401de921cd38bc0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fcb9f74c06b88ae17ac76d2ad07db55a6f3200aa9dcba5302b2e22aa9b0e6c6f2415ee630ef42d3e66849e7795ba49a0ed80eaa7278cfa3a7f370538352bd5de472501bae5ee0edacf989743ce6cfe11023cbe58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d16bcdeb1c25fdc5b9755b2a3f4f5ef0f75a2519435a484703c71395b9b23f8362b1b92d8d962ac134fbf15c3f33b78c7a6686ee465ce772fce4ac8680ae89a519ee6e64639186e9c23c4e3ecd19a1bfa1361f23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ebc3786ffd808a95e19b3cf967b6eaec0116fbeb63b2d4d8df6b8a2d2caf299655cb75758c6eff2211827bd3e0dce5d8bf01932902d6aabe7283d1070b15e62a1dd3178377c52e1e1907600289250db07f7cf411;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a735d6e7fe4a08d9e33f33b7d77261340b34b9211af1824b9dd201daa746488d357f0a51092f02a131f8b3baf37676805a9f13d7efa98dc76e0f78c8e868a3c97896fbca0934830bb1c0a06158ba50f6e460f2fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h498e330c8a871f875874bda1b998729d3e95c3d1afdf21ab65441dab5b0d148c2dfedc100b4952ae5891fee872bbeb4bc35714b51bcb203f2ce16022475b998cbeb2454f0989ab8328400645f4c857b9a2ffd9cea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd18430cc845d3679e846f45eea446a8242a392e0be2776bfad3744192ba3fdea907194fa8af272161f3e8fff26f96de608eeba02836cd9f12f9e4ba5632dd63ea01f355a6c8ac95cd0e75136c9e0f3cedc0b0764d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30c76bdf38c50cf63a7b9fab74ef36176a81f71d6acd83f945b9c34aadcf31bfeec104274eb98cb9c932b08373b6459b213c5441ed2a7ed7d241a81cd82ea3e82e28a79973cb715410f16723b06464d566b65d8ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8eda4dc910d62ff6a46a28a85407105ddafea6a3e75894543f2ded4c642c920c37cdf49a50b0b1deede640e262d965cb350afe384b2f1af20001a8a040ee26dd3d320c8f759ac2885921c5811258a4d8d27433aeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d8b617be342586759561c74e27069ecf26cc02224318b9ab807ab22a9b80c32eb978bad73a7e6811909d6a4a8392aaa3a9525baa6ae1f14491af7958be11c806ef42d9638544f515da626444f1cd16319b2770fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80615a4c53ffcce0bd088ca36b9cbb8935f0b731e62b86958232e53de82be02f9a10772169460e33c9c43ccfe7fdbc280e0a03bb7a6364004fd99d37d0fbd30238fa0d9455bb8faae84773350c0c4b22d72bbbfb4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha541b3e53702a49cdf82f3f46a3798e5a4f10efc797f38624ac26b575b59ed5448664a5753f68d57f84e8e34a43c6f049afe286e8d5a020b12de1b91af47a5720f5091b56669f7db899ddd44214656c5e88e1f0f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd44f9cddad776fc2b7a309962411377ed2dde35380983a63b705e567db34359f733491fced2b2d37b513174e03eafd5422acb0f308d7968f73405f1c949b2783c9ab0df42b543cf671dfcb7e122e8bdc2cb550a06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4f4f0df94b8f11abe882d5d6ca9fff69c97eb7942a8072cbae20316f60388610a023b9516f48bc3865b423d459bcb298f7faf01ba87f04b3aca04487d7f10e21a977aa2e50d6a53c5cab2772074e3de0b37e6a49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7aeec0054b62d8c17a322e7523213d1f38411ec5bd3775ff7265ac444e4bdeb3cc9d33549416c13b24ac665d8c26fc27df13b7c441d1cf2d5efbd4c7fde52dd2c1aa9c4b09ace0777e051a1cca37802fb6774954;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had7283894fcb012d2acfe8260a25059ccd47c1b5ebbe11e2d7be505f145edf323871c6b04d9a1cefc4613f6b04131142fe4bba4196618e602ebedcebaab7f3136beb758cf7475fc894b10a0aac526b22148f94607;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ace906f22d697f41213ada012a51c66c2dc29ee3c663de1c95a064636b1ad3d528dcc80bfca0e3731d43b5d03ff5aa4ef6be04e8f588c199fa2c9e8a2f14fefa13ba5f4ab944757b5ec6584a9bef531bf189c9ab;
        #1
        $finish();
    end
endmodule
