module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [18:0] src20;
    reg [17:0] src21;
    reg [16:0] src22;
    reg [15:0] src23;
    reg [14:0] src24;
    reg [13:0] src25;
    reg [12:0] src26;
    reg [11:0] src27;
    reg [10:0] src28;
    reg [9:0] src29;
    reg [8:0] src30;
    reg [7:0] src31;
    reg [6:0] src32;
    reg [5:0] src33;
    reg [4:0] src34;
    reg [3:0] src35;
    reg [2:0] src36;
    reg [1:0] src37;
    reg [0:0] src38;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3])<<35) + ((src36[0] + src36[1] + src36[2])<<36) + ((src37[0] + src37[1])<<37) + ((src38[0])<<38);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc60839bb673d2fe23b472055dde3d4e66f5380b292b266f6c74a730eb25dcbd5e01cc969deb9179652443ba898e2dcda1e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff6e3c49f8be0e85df555b6a227a4aba7e9715c158d7f0f095704ba16331844f48663bafd9fc8a3d171fec660c2deaa26f6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7017a1030549b6ac0dcdf8f735c38277b6bf21e6f01c4984145a10781420a62972a17a1e63f49db8af1e1fe5bce104c035aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69546cef0d679b66d6dc1c8ab943087be32ae15240a9434635740d6847b6bf4eb37f489c4c2f3a03edbff440e128d6a794f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h989f70a22f771bd433950e9e2408542325fe3fc3f28af6a9a58b5f7075aad3ce2e4aa38c6a799f826c053674800797aa4280;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56d62a9780c69345403ad69b8e9b2895330d4e3324b647a960a92a8562af38ff6e0614e137e229519722567bf6056c546ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e2200b86bc46f3df87d87dfaea0b25667485d038f211008a385b3de6e4f371389caf50001d3dd652ece5dc1a1813e0c07e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h748c0d55694ce49b5cf6673c7b368e14b0c91a4625c639907b21420182aec2bc6d62ebb235766b16e0730bf74a4ae5389d8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11c8a62ee085e0d05a274b4bbc72cbd2cd5dec159058d04bf527d43504e8c204ff841024a502397384f52d7dd97ba74226b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55cdd50d2f9f5516194b9a2359869b4dcc2bcc1ad9f77450f12312ea33673e360096ead7cbfa8a2e9383f94c534bf1a572d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h968578fe29705b876eb6d22af36414d4d7a77806922f547e752c4f93b6e213a03658cb37da03040826c7be21ada219d31a4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h659ef38c5dc5dce85f9dbf133c7ea457f58e9d8177810c91753549d020c7043aa1b080e4fcc16c2e3e18999b0c5c03ceeaf7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b8b95995ed94009cccebccbb6dca22b4ea14c22053f84e9c2f7c46a8263df8ed4a1f7f587ed1a248587ea71dded95113d3f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd43fc018f31d719c9e96ff6713210ff982d6190ec4ef635fc57b5e16f61bdd8928e7648107031373706e7f5357f2b259cf6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5e1954dbeea74100226d6e4e86d045722fbb89114661c5f1086672eedeffeb0d7ade9d2757ff0913ecd10be99a2e0ce908a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd70b716439e977c3e7f259fe2e7a443f4718318b8366159ba0fb6cb68765e39e1f99888657f06e44b001bc1084329d3924d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7289be3e124e035787a1dfd712daa0e79f75cd827310b786f289af5f08ebfea2a6942157a1472ec9cb1a21487d17a30cebf8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27b20c0706ea66ffc21273a702b65ead19a920ffc8929588872f554a83259951e19684ee9d3f010aee615247ac2ff9b27a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h627ab704efbfdc99732b9b874a6fffdcc687b8aefe286b18662ef665fd2c1b2910020185efe4ca395a47b86b417ab440006c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h809984d6ec8d7dc1ecbc00dca718655c4e2e2b7c666e6a4df5cf30ccc506b9a7f92c233a14180ee99c976d89f03a078cea55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b50413de9143298ed9b9df4680dfa14a96ecc07aeebc5ea5e75ac663f76a09c9ce0ac9d716bde6f41f6e9d467b55de6f640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2b0863a517b4be74e050a445334b82d7d179fa4c443b89fafe2ea2eac7ce6322dc422a8b06f8176363dba84f4b9677871b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18835e46cb27c683002f1b961f8c1757f0894439709d09196e2b141e47e294cc2864f1ffcca2c6b3c79b3d439624aa1929b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf750d4d8d0657bad433aecddbd75a61ce1d197ed0dc2e08780a16c03bbf9aa5fd468616a9f3b554edbb3a83d5fe926b71fb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaef2448d32c2ec536ebfaf5fc63abad5cce940d0b365f841ae95c8389b123a66cdebb6ad4d3f3c53ab553d4dd4eb1e93a23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ba9e7f3d7181c39e3ff5166e46167c331788eb4616ed593fa390e945165e4693a20d8829dc22bf192bd91fa515d0a2defe8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18671166fb837a8ea1d14757617dd8a57f983efe72a5bc97695e76e9f6b0ce55cc0910e2718e62ff03f33b2c16b9271ac0f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he390050f140e766f59b64ec702465465815cb967afa438c7313440da4d36c7c090894645130a493418bef4dd986ca7fcd251;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d1ac8ec739d820479bc00e5f0ec04f9707c5c10bdb28043bc0c17e567f74e76e79a68f03886c08db09370c942d2de74b806;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf4bddc273df8596246312cec34b32e156e4b222518d45d4ff62c506ea8ee65389f63d1df9548d6b11b20369031d0aa04899;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h668e92da8ef31f10791431349b093599c005ccc271f1a5882f6806c9398ec1752d5953aa23a7c56bcd3fcd6c0b132f295f02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9715fc70e057a30b0edd4c38c340a6b598013d6d1ed8130413e7ec8766387835fc457c93752fce5eaed3b8823a6e06c2dd0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc410d98a32727bfd787ed61fb5513f4a265d586e4db1f2b19e3e2d5e155e4702c82cd24c1ddfedf47078c6c3ec6e0523380;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc22c2d913d54947d4ea48ec89f79c0a42eca47448f5d0c82fa9f84df291301b297245fe23c5518bc89ae0fd53bf8cb391ece;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e4680afc8d43f8a4e83d36d11b47de4790325968e42ebb2df27df2d3582043e2efe4248a6e3a7bcccc2330658b175992ec0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99d3d737c8cb7d8ec2ca1cecabda225598651d8bb367dec36e60cdcc81ef1b111cfc8bbd047e49ef777478f0fec0287f89b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a5ceabbca789095c9f89f852db6b92d9c225f3bdfc2e5179ffd5c8f36051da0c29add544ab18e5fcc97b2b62264d36d802b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f0795d346279ff645973c111c4114dec7535dfa00c6804fe8a5461cda1a325c6635172fd083a3f3595d50dd6a50d0f08bac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b0b8a9574f922cdc09a28e929b93fabcf08f2a976249d6172b585631ece284753d0a515d3ea54ceb4d293d6168d2d8cbe1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h595b86c4a1166d800f1f046974b160349f2f66a99a6ac5d0914bcbc7f5a5a5ae612b80f93d4fc1ac7032cf2ea9fab98c94bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h405e076805f5f834ba2ec6e60f693c547d4ad1d61124e733a04e25fb4b74dae6bb64102bffa1f0017a4f2cc1c983e37ecc4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59ea1f1e410c5a83198ff254fa8eb5dc2092b334c7fbbcf99c5aaf5eb76778728983ced636afdf1cca8b1b7974da82035abe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0482a4d453c2d0ac14900cd7a41c2c8725556ce5f92abd21b7804d7262a4d49223d66f0aa6541581e942a6489adaf204733;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fd7cf3a3cd7bcdc1faf7f71198d59e45a04c0678196edb7c359ab5f9c6ce6ff8dbd71ec420068ae3697d2a5bd9a5731a47c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ba3fe6cc35cec90071abd3b12a9a2381775f29c1c3ef41c2722c6288d07b63977262a352e227c971772f6a4c9a72d7c0c5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb406863b2c84e31cfdfed68e45510b4d86ce0f618c2fb01f718efc4b9fc5116bc2b184b32ea8009fa04c18679eda770cf7c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1572e71aa523ef34f49e7dbd3cc77497c830425f580827ec488bb97ad61c3c31d0b3ee043e2ba8d8fc4bb0890c62cee95f5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbaa0ed829321ecf0b8c2726ecd64cf8aea34e48e92367a98000174fd417fd42549ed7e38e0217c607c9d1b4f690c16eb5597;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1135fd6a38ea6745f960150b57557be8e6b107011c67c6ce97a1777afd915e6b5603eacbd3d8787e136edb641da374ba8b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9053d79e24633018453119e6c8e03f588615b5f061f3105f113abe9fee4fe0c55a405ed7c76172c7f446d638b5e6f03f20e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1b6d475a54456a23c337823af4237b1a9b8ccba66666cc0f144a0a7ad8678c3afab09b921a1eec70efbf10d74eba0936ad1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d754c6a257fdc81b076a5dce77cf9b6cf295695556638fc781b43c1eeb011b9d7a2b190ecddcf5bd96190288f4d73452242;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a0e7a81c806473ff43a2a84245339d3cdf4555fc9ca1870af6058a0aba5469a913fc8b64bec74f9f1bf60fae4bad9c5c17b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13bb9b1d6c5dd27bd1c4a26460c2172589ce841c7d8c17f8f7393078b4cac4be3582dd2c1dc82677966afc61c31af9e08b03;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc46d69e815f075db99fa0903f09f079c99e4045fc8c89dd55a78b3f3fda81e34bd919c6e5804c9ed6371d510a59fef204fb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70103fcb6b51b4a0ae03d264991e08244aab5031aeae26e2556d69b695c2fb9baca17a4c0e51a2ea45996453ea1f388e88d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa3237ed76cd2c1677be55622cc8ad2198056fc922879c4ef435676e37558e6a41c64d7eaa53b2d50cb78cd2103c0c4e2c78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8b33e8bf519b064e1d63496f9e24bd36bd3b8e9df9416adb1ef9f354e9eb87123e7bd8d2fb2cf6eafdc6b16ddeb75e359c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd62e3d0f0d8becc49231e3e51f8146df652be1835bc0439aef23050a5aed24304633a42e9d727d7846fc584a98b44170f5d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc4a1308da95c005f764da17f7b55af2ff7a9604580f93a8389f4f0ea701e0cd8accfcff6688c1c67fcf32b0fc4990af3c46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadc51c7e1386e0071e823cf9d5ecede14097f7a2b7b8fabdc755d28b3db02f9d6bed1c70942bd4cc014c033e5a9ab9395689;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0bd351e99e6ba469717565226f0012fa4cc4a1e4db80fa6137127c611dab0f61c029b38859bf000643f761de763864459f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4712c42ea9c4545578263a3c64762066a220c7afe5cad6a788fa5f83e65d3ab584a4f26a459a226d5a8f880555ee58191202;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h551faec287cc88c902f38c16d74aff1d7420b7e16ed37608c452fba89bf3b026d33eee4c49b418fe646f84adee5449dbf1ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26611441b2aa21e83a66caaa78bf7ccedac5654593bdf58bf818b51e0e832a1241251e397805b322a0917d548a0ef5c957a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e421b610a523a58f819a9c45f6a0a8122fc3679d005af1e576416df88e0313b1bc363b7cf9d2d9b4564ecc47c0b0e65a8a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc910d3764e0b8605eaf6406d0eddd0c376cec440fb0b4a4da9e18367d3b1ae34def2522f2501521d462b01c3631adc73422b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5f3722d92256ad17d6149fbe3c2909eb94b8308b1be95cca1bb08db5df269442f592436d05124446227353173fe2a214b3d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8965da4d941a7a06f7424457d61871f9c9b8c6872009c00a850808f1fbe30889c00d2f08310414f5ce2512b52e201372dac0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45a7c0f1ee1af6dd595fa1d32395242aae898225a2c05e0f94e593d94869546aae5d137b45655c280f95d25ef1e31cab357a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfda370177fd061ba9934b76d9a3bbe8027d30075af4a4bdde7c839dd251310a1b1f18ba750afccd5870922f586ce1eb90945;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h762f38adbd01fb9701fec17283a89ffd0f78ebf0c33fd1b56ac7d8cd67c95210221663cdd72b5ee52125513998b73a8146a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdba9096b4bf9b23575445fc67e9d699bec8a74ff50d9472fc62c30cc8038728c6d20c0b28d013b6851a4136a0e56e6710904;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha91fb13654df73f54f0ecf6aacc391a4cb3ea97f1e8c762129a7250f452797a051dc6f2f329b984023ac1f61612ceb3d5d56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb432864a1bae089b8f7421a9a36562b5b40cfc6e3418999b4c4e84b8e1c349e13c96370240ed9299eb971bb0902eb351e75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc03def32fcc191d894a059f2b72627031382a3cccc1a55f49bb0669088da26acef3c3349d63d8ee78e05a4e316c541998f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd36bd8843fdb38584a3eea6f7751302043716b185dd3416ba81d87ad6eed249d34ad1b95170e9458648f924c502c1fcca7cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h809c21eac5c7ab66c6a21771ac6e8cca90d255363d7ce7244068433b9c2badd204fc4808cd48042cb4909fbc0f7ef861a9ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2fef5259e66bc83e6fa53c578134f53b310082dcdd34511da1c28fa0caf7385dc3c4e11441333f347afe25c250eedadf860;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6905106eb23c99b173636156da5a527961b9d6043747776088615ba64d1f062d1f5a807ef59a943908cc7716a14d095c714;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf14c187bc496f221cc7e89726391424488150752e23a7916dd4152d9a023b653b5db194bf342913de9cd898b1e6a5c401a72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf422327598f5a0a50788e283f166c5d45a5b5f9d90cc5eef3356b963cd79c937240d211dad511c2872ba2a8b36465d38c29d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c39793c90161b120cae51d5a44cd9efbd2244d133f8aeb63f51d729311016c589447ef0d349aab1f15002faf056eb1ab1f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0d7c380fdf31f40f22919795c6abca3ef309480a417d6d6a9e0c8e61c142cdffeb744cb43ed91a58dcd146761ce81b5930a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h767db1a92befe3a4cd57ff848527bcf7d0d307d4ef5bb003710e0f67b9b855eb6587eb2297b7f64c8fc2500bd1d056075c74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2304044a939296c9666c1f60b242e1cccd60e4931082fc09521276dfa867aa239012e2eb96f6473c233569c60a024ab3b02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cddcf29fc9271881d5afa8b65b5cebfd8dc324068757f76b19acd7babde8bd75d809d5ddcad7f7a36367f07f0983b9662a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcea1744d32a064350c3d7eadd8b8afb42a90d6adcf1a25364b7eda3cdbaded5b3ad2387cfb477275db5795b0524fecb59cd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda98a0c3effbbe67729b6aa7473b97ddaf4b7dd7367c013c76f109bea8f87f226a24d89f167614d85ff5123f58c758f273db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h115d16a03c35bcc845b2c29c26d383170ad74fa16e5864ba2bfcf7aa2ce3da96c52e8d1679e57542b5789a6c8db726be90c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd804d51e7fb1e62e742663c27787666c2ae1dd5cf32633c0980f29be4df5f105b654226e912a01529d33af0ff4fd588528;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3731401df09f522d2f4817f1fdeadc391bf1f969d2f2aab7aa0d60d63d4c04c957e4be7b9127e263f7dfaf019ffdcf36d01f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b2994da1033ad0ab2ba7e8d05224ddd1d7648d89da9050c6096abe3cb5b5aa957b36d62a28c64494295b5609d1767837d01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdca5c3bd8033969f45115432fcfb2a19c2d2710e03cfa7a983217e3d713804ef831480ea8ab31ae30ca30d88f706b626540;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb5b465173695540725bef93d96b96ad5fa7863da0a2e233e8ded9669cd0783ad6972672dec20a161bbffb5901b133a3f176;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7939f9001e081814eb9070cbc087ba0d84ffd863560494be88eedd6a20252fb21ffcbc771ce5dcff26092d0b859b9e64f6f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51d74e85a6335eae6a969e1a1d885a21d06815266dd3cb5c2a6e6f8e88a900c645f9b1f80e54d32be63886a14f0b0d307787;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h212d33516a5de2ab45e2d4b91423be1a8dd10bf497306933c1c66cd3ba37865c34a6352aadca408a31a13f3c5c3188ba83eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h697778b641df087cdd2fdf07eacba362e3ea88e04ed86812592bb9b9b72eee5b094f61fad693d484233c14992df9ef699dfe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f42f9ac51885e8cc0e3cd52e216bf33d85d5649d842c0ee1b48d0c1330dbe78b0daef2c14edf131c1e322e5d094e167f63e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0ff075303327494de6ef15a0e55c6e85641defb08ceff02fef2e6fe7451a476a7f8415e5d7f229a1564c76bdeb43a474983;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6a3a3d3a30b9edc1d56263b18788e0482ab37b36cebc89521e43617d8f1aa0e1b41fc346377a5d5094f8c073e064530b9e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4a948866f7c700a1a6f156e851adaa04e013d25191690097fe67097f5ca5ba77e572e054424371d84897879e25334e5c759;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeb7b145ab7b4c1ddc5f93756a51548a8b594af9c14f27a5715e5aed216813c84b4a08c4d18ab9db2710795c36b150b15df9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b7c675d89ec24577046a4eb3fd936cbdc27d07b058e40dfc035b953d6687fbd8cdb9cc8ee7777a930f70ee5bddf2a137a9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d058d45d3c32b7bc454e57e8e710cf3fcd1b786df86bed008a3f898dd9ddbcc6f20e02aca0febda3fea184699639179648e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d926ac288fd84e3194ac6eb52be83a430779842cfcbfb52e13a4973e35e03e16a95423273401c7b09848cb7e4467385b060;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8847e67eb2f0e4e57e6942fdf6a53830c238e29876d8f0f4200e00a0eeb25bce9a4f52cefee9cc93eb542eb70c7a7b7cbbd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha42ea735447114d90ca98ad71cc665be1ae61fdc17e6cd5d90d3d011177187f82726c64f250bf706b70f82a9166d9b75577d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87b150f1b5059232f8ab61ab2c7e565b1549c63e1130c51ac699aba78e499cd950e826cc89f72879f510361ed0b566cfc330;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a7122e41068be9a21fd71c51f48fd977e606dc06e4441632443a2861568ba6b9c6c032f2d99a34c6d116b940272bf96cd0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6549259fb3fcb02b9dbe384a3541886d72a621584b846fb7c1a0f913561afa597fadbb1ab65adeee28a914d5ef88c7b4375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haae5d9480e6b8388b443d9d223574d76483bfc04bf50096e6fdf931e9f9e3c80a760476878ce46d4ab85af05165953836109;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he727ea0290339e69bf6f165fd08ccc9b918d05391701a7b52bacbecb7f3d2066dd6379d51ed7f02037728c431819a0158785;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12b435ebbd1ec0b5c2114504ae7b2ad313f5ce844b6ffb99861289a6d2a7d9dba59926138de2ad3c12a2654884bc76971fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f438dbfd3aef65281b4ebd06ead6c726dbafeadda4a6ac2eef660b82737d82b9161a6e2266e2e874a3c7932855ccf1ca132;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9aff15d0935c19efcffe2dea754962b90ffdffbaac6a20394bbf685d43dd3ae60930396d8c1c8a4d14655530e2d35df130d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5456835553b9d744c01ad1268d5632832457c6655f01a2c4f120ae16e26d93cbc4b9dfbfb86162dcbd1513159c69ee2a2293;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83415433662e24e82302e2fb4f0418f56fdbd34ea262ca5be864827862676cf613409b093f0f53e7a65a76c7fb6febed63e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e498a768e6fb18759ea291046934440550c91b0bb265ac1fcb50f2c64a1d559139e9ad1b7c18670d7ab8eceb7a99e52fc11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5f093472ddbe49b0f9813e1bd5bd19cd44c3e6e24a95cc580f412f1463e639921d874da68d4a5f066e431d92865f952324f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h929747cc588a84e79f436b0d49bf8971e0e811c431412168b717b1f2d472866f0087fb4bf89762f1c14396b07e7a0eb9e927;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62120cfd0f70b1cd9adc67304e45654d8768402a89aea9e5617bbb06f73ac43bd7361a67d655596b8f7210467cc64362e30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4d63462d0aa3a7a3e9c87464874009b7b35dbf9b69c086732f4fb9aa76429ee4169e903313486efccb6e9b29c439fc8cf72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e01c979fc652c12525d39fc597b1642fab073c14f44f4f2137a5710671a688d226c2448a62cd448b10f5bc947fb8da9f3d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7bdfb791a7ddadafe10706dd94088ae352f5e11e65a73df4a7284c8774394072c0f0af16e2aa30668604eec01038c44b58;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66c39cdbcac12267f61f4d7de7c561f8a86fdbe027bfeb30e136c0d08d3a9c77f51229ae80cab43f9e6c02063322c0884b8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf777dcad8a0fe44f35da544072534fb8e8d6cc4b5f5d6c657009e0e4d5622689095153021bcd8963fa32e3d40c782812af79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d9674f2ecbd8961a030740abee31070bfccf76d43e08d9d54589b1ec6d45436fca11b237dbe102db7bc531733731c62c263;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he53bb756199a253ac847243325d278635456011092e1c7ae0ddc3a0152e867b352adcb46ec8bd73cc4cce3007a1fc300d385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc283e073fb6c4b9960586dd46359b39cc78d76630ad6a2bfe35a124b837c11d2bc13de1c0d6774d58ee21aba37d482ddd334;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40c8d409a1a7865d61beb1f703faa333891ab0f185b3775eed46d596b0f300bcb0d5c71e58fab961d252b4cf20a45dd5d92b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f54ff8cfb85a82411380a57aad567a2884fb5bea09fd104a01ac48e8805c64ff2ef5e715d996e73567f0f011c6065c37d52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17b1c7cde52fd83ced22b909e040e04996c823ab7de3f4e8b40ffade2b41ea51eed068afd3c1ecee61edc7a0f51e4ed58851;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bd9651cc10e2f0045f81c545d2ead774d39172bff70ae570db030134b871582f569a29e91fd354fa06c2a81f0db3ee6bdaf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h237ab841ce01f9f6387e2d0f8665b4459fdd6d143b3d4660e8036a4898ea5ec3cfdd689c09263aa9dcc1ed34d185d9d1b283;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35a8905a963ef1ebfbeb8d7d2c3f3ef770f318859d6b765a917da275c4cf314497ec01549bb584ec7e7a4eb73ae1ee59f4fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a2b78ab67d6371dcc9add9d2bef1aa8bd00c66804d58311a5f4f6082e88588250e935995370f2488fef2552161c3c67a8d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc46cb68512560496005c28b3f5eb052a4ed97650166a0dfe31f0304b44d0aaf58731b9db9826b40955d37213b465a2aa97b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82d32a8005df55205f07af54937d8166a7cffeec5b9d3ffb7edbf5f0ce599e96750aec192fbfd56e26c8b57966ca474b0a6a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c5b0f0c108a832048e8dfd4d814af088a8e8652853b87806fc8e59db519c41fdf1da500e0146f777c2de9f63b616ae54968;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9caeb8daa2f75de5372ac04304a2a4cf2ea5390ebc0b364153e42261941bdf8205ef319a3cb8ee203a48055bcfa09c209da5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2c5add8e9e05963e0dbb91c9b2e2b177e697d385c1ca3480af53eeda8b18d230bc2643ed4e07334448428d6d8d2fde82911;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2004891c436d092db14d877983690e45b5d46878479dd4447e0eecc12ba98a8f8dc927cbd78000ebbd5902d55a7fac72a557;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h637383103c25fab5f42a77a896907c9bdf6637ee566f09e50f396d5e38c25f341323dacfd9e0438fec91727cf59f4ac5a9ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha896993b1e8f473b07c654c94d6f897789a2de0ad294e7207573cbadc5f0aa43b706fcdb39f25a0b49c6bf622c2b4b236adb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd2e6e23fa27eaf9745c35fab314dc629790302a2d738cb0a4abe53d63faaafffd98ff320bac013f7ca96aea57bd9fab1f6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he96090dee7a1399574f946b16a344d191605c99043cceda1898a46f57451e833386ccdad424b86213602a234b36a951881ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7be903168f576b2c37749a8403303453318e1b0f2b67eb089ddd93529196bc42ca552a318fc2fe36d7483abb7af45c737b6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85430814145d65313a12ad29651dff9a3981064d464d80a663c08df9c078903928c108711503c4d9606f2dafa04dd4b48a8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d8d4d1e251dc1aae423da92ef470ad05fb02e5b85b78f4af099a4138997c7c0ba0f78e076f63973fc3e5600a464a1d1b10a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9b07a83a3ba0c295b6115536981040564de7d04be2718c0090e8c6a1de4bceec56f2ccbab16aedff85f4630d305cc4c569f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7778b36d41cdad7b47c1853a9341573527d2deb5063aba69268480d83d77a24292067b88a9684fb3958fc6d9e0313b7efd81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcba0fdf5a9ef0f17e9f82ccf2bcca6e8648d16c92306015d0da5f3be027fcafd7d63d0837c12404ec8595243cd929c7fdaf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b58939ac200e71645dcc372c4afcc6592e8fa7dd6563852c47b5623b5fac8c53631918af2bc73794e8fb23f94803e586eb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cb687ca98f888e59def69046fb7fec676413cc1ba4b65c42e9a511c56c8b9c7acc7a0b68e9fa9f55750e4cfdbaeb69b8c8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bd5ba798a504897bfe804ee861d45ef4f4ad8e1de60147fe1282104162ed88b646d08d2f1c3981e12b851403546f10bdb26;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h516a9532a8de1ef222ff36a52963b0e01fe363e840054e8f459eaa14a15cf7570c41d300ffe89eb905e89fdbdc303310be67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc00f163781f0f2108b84535151ef5a9c7fd34032ab42f2d20b7e327f3e49b92e5d05d4642bf62cc57d5fc22cc22ebc601af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf85744019d92406ef86e6b338380ab00420b60af6a9661acc1ca58c8423dba2ff88916344f24398d113f7359e48034ffad31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf191d4b8e12aa57f73c3cefacb13386f0c53dcfd4f00fedf007afbf34edf8ac46e04104038fe0c65339aba32e38dc340f22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb7e4c43eb740af2b8b5aed5bc1d193e13657a7bed86218d1e62ee09aaa11501ed802913c4e96d8321edf98175ca630aab8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61de6881d288870dfced2d89fae7d11c66b1acc6cd55050c4a19813b06c81b48d7ceada469f56d0d75c5b2c59cdee2f4dbb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae2ada6a47c344d8e9ff166db7ce89dafe4643a1d43efa23717950f5e51caa4d29f247959c19a96f088abe86f1e3715ec3e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9f6d20a9379898adc802cc7119fc1ee2b7425ed29cb437c7965d916ab0704f4b6c1498b8b703a2c9f9e3cd1893cc42814b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36206ebffaccc47ca2dfab12181c7e2c1a2ace28257f0df410f6e2f8c28a1f21c71e8e3f25e3cb0752bd4481453f3245d791;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72a776a8a247f9752c382e3a78d80628a378563855c1b53353c046d70538828f89c59c777d3af317ac33d85130f46d9d490c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f98196c9aa0f226835975beb7eed3a93adf0046fab148a8a43b9612ff3019ae0c1c3b9b9d9596aceac2a40c3f270797b2ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he981bba0a4722a0cb59e8d48f659fdb08c9dd7f3b3111e49f585eab450f9179e483591b07464b5fbad018a27ee98e733c780;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde86bd8ccaa397f5c25c5aa5c4c1f6ab0c1188b06b0b773cfd785a622753265c58164776794df599607269914bbb1a13bc74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbabcd5a1ebd97fb2bb2dc2ecf51c6f46fd095dd87d5dbcd845aa10dad2dc36914bf0132b97cc9d057b3ce44eccfffffce66a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fd45d3bebdf05da4c398d140805b970635b774e1c0f1ac58dccb2a67e3f2bc784b8f6ad6fe3e65c1a86b241fd9a420a7f8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c054c45c959206ac1874e73faaffb017548c6bd3c3c5e755a1db0903445d7906e655aef29f064c1935d2e1acddf7d4edd50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h110d4609c2fd361531af914bb504a5e84df877bcbe98e0b6f5c0d657acb5585b01dc9360a811cf7afa4674a6706b9ab2fdc5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47c32f3628debd5139fe6da8ed50849d9d09e117f011125071567b99ac6e2eedd7b58455d062f2be60f2c29afebd2b8be7cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbd1c6ecdaed68232600f0dc12c9901da528c4c70fc59a725b300bc65d5053f90fec42c2208c29a31ae77b06ee7e1a9f25be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c8fc3a3eec6c2897ce5bb23591232d691bb8fbb5891638171092d12d732b3dd5a0db8e0c88614b0bd325c0af58f3cbd7f44;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a98fd3251fea286ef144a891ffb42684512c5f7bea852d6123a7f57231c510202a5f3a4d2490b817ec886537443b4ae54cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb5b7d3cf79389fb8c4bfae73c5ef8f2611912c19eb0cd752d3da21eba5d44bdbb233935fc33f99d65944743087a6c3c61ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd20c209b8800c49d526ba3571d1b6e19a90334dadd77bf7dd71b18ff39b51484629f1bc33634017795be0aaba84d2459746b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c5037c36ebb5f13640cb8d724c4442c3bb3ae1ae23d379086ab64580f96be6513e2b6ba9d57366e2d7dfec0fcdc8dcea33d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a61e38339e152fa60bb4833e5bfc400734a4d0db5be1ab51d567214b4b34e8032168ca44292a1a52e9a759f69d3a4007104;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf16e09a05fc98396f211b392197629aae7521ba9515d11c970e691b9919db76b520d9498f85d6747913011c62ff4696d3563;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1b90f2ccee74d1160b57a8f64a9bbd39c4e01632bad4afa76c31ded1ce95365652e7958cf169a00d9af8decdb95e0e0d957;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h550a2a24e2e763be24f5e5956449562e699850532a195658ae684b87ed0accaaeccdbecd86ab8c0a057e0313d3e85ff3d5c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a6b4c342a3d4a1f73f0fffd05b93500d4d5f59d61918914e6f577745e9cf860c07a0ab03ce9d45483b229e40f90bad90b8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c594364bdfede7c92ae3a3abb0110922e49acf88b9a75fedbc5a4d3b8835c0cd09046c6213dd8958734bf688a022c8986fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ba5ba426f57b492e195e07180774fcac5109413d888a65b2e72359ed27ebca0ad68a0951d0e514ee25e01c896010c212ef4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc31908a18a9a5732e8dcf0deb9cf59b1571eafa2c7d5f041604d64c163bb055faf79f13b08b6a5dc82c45d57052124c303a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6436728706f0ad6ff4b5b534c19addf56122e8de4b2f67a7e6b5f1a21a3eb58aacc2c812a9530cec875053f2c4b3f593118d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb221b2117caf404b4f495c14db2be7ad3b1869c625f5cbc45fc2e6ea30ea7512174e76c77247a3e68fe9998cf879ddea707;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5632fe90b502d3066a20d0484a1a09f01209174d216dfadd8e720befdb8c65c6f61b23986d4128d2dfd71177bda920f44dff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5471bc806716bd928864ea32508265685aa01499e4e152a03f7ba04d8374a74ee79d45e9465ad679c3606182da288c55d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5da6820f6bef3080861c46418a60d6e13925738c73e352ce02d2a266ec2ad86dfd8557b6a2461aa874d55601a04446723f61;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf3312f8460150115b233cf95feeb527cf5f4c90bb5612329ed28b77cf6540b23e4677ad2f66eaccc36f0ac779e8689eb6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79feac2b9f372a9391049fcf4f2d78f9dea3d64e8b8b0ce21cd9961e932f3d77c9de24496f93f9060d0958e74b59295b7f68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17ccef43b94c20ff07532b1ba12d4ab2b8d11671503dd58140c284281a24853e9e2c1a243d41be199ce9c7d3d5a260fa64b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd848711bba44881312f98913d5d227fdb705b44f7b0cc8c22a2e345b130bfa3ef8b96ff701d2d424cf53814ab5feaa2e21d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0c3ac41b47bb847d1d8c2708a0fe3e234d4693674bb3f45ab240aa3201fc7b6b96046610f6328acca4f30319e61804c72db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7381ec397c84914a971447ce3a62856389b8c90ad701b4c76a5b8d1515d14a6c6fadba1cb2b527a416d57c73666a8112650;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a8ef4714b07f8896501b1d96655dc7b88e0db41bb02c31687cb7d1d036913ad9aebd4eb237e5d7bbc97bf6ee697b5546555;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52f96630fe7385308f10cb4f14a8a00db582dde39c4d82c09c404cce923a04a894b8b5d15fe4d07b0af817d62c5f3282fc30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h742d919949bdb27fdf51469d7c65b57635b693d3bce8b82f5592545146dee0db9e9d410ba124750fe6306b2811d1a2ee4fc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3aeacff24849bb623d5dd7d6b94684ed7aada24723b759b17d043b62c04f1eed1e5390a0383077cc4f0ea41bacb16101a82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha232dc090e3b0e00deda54975d3eb05cedb348f30598a52fcedf92e47026c9263446e5293b8a001fc65a4c1f367b358a1187;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h134175d313cf6d6762788fe52d722d4214a4d9b6eab3089c269a2ff7c3df27d2294b817f025a7a32009b6ee540af9ee34410;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he631a2ceb3e5d59a43968e7bf8f08d4b7b5ae8d60661f63f1964501395300d8af78e9f9c12db8ba4185df822554921c6c71f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h649db25d7a94f2d3ac24fb06774e6f2f02ae2371658fff92ad11785d152e5957bf8996045d5925cae6a59074a793fcbf8771;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heec0da6484ad55f8e6c10a0b03ef9ae96bf9ba1a8a8fdaa5f3c59369ede395bf529c1e93867daee30739ac88f30862a08b4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb7d8a2a5c35f6929c4f0516faed56a78ec18ebb89e7fd142724f97b8f7a27ba2908ae7061b107c3b12d781ff71d311141f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1ba141b553af7be06a8a52cb72939116d34467b83be3cdb10702bdef1b8c30ad7b49c189fe2e9f891a2882816866063554d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e6c89dced7cda4a12ddbe73a1199c9ac82f54137507c9486a5d57b5b7ac428c37a6fe22610a04a6c49e63fbd3c39f180f8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4d34d99bb04091857267d8cdd66fa3ac97e5f908d761a35728411a3b2838efd3be4a87d22d075fa71145eae945cb0d14578;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebca0064bd488f9937411703f6089a946d0bdb68e7740eee41934189fc27fd667451a843aec6aa70f72c175fa50947c1d43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc16e3b5d45506180c30774cda5afb17e0ae2d59db29583531954c84189f8fafb371c3ea172a8cfedf4d2d45091f744656bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90a36ee537773f8fb3dc9c11a43c960ad0ec9f9a4e0725a2546724edc8bc714b338533b14f8d61e93edb34ca2483eada8eb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e8a4e01fd2ac4614d238aa8ed546f47fd381560857505614cbdd0187f6a9a4142b7d535f1109400d375cb821403852c7b56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f129a3bb781bc9e751c26a3b3fd65e097e2da4e42f13ca7a7eaf5bec1b6447c86db6bd3cf5a1b33757cd5a852eed97e43ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f4bfbb5d37023bb0dfcdef9ccec2031991d340df6792b9979a6c04d225f439d058c87760240b415b19355bdcdef9334475a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d74e14827f68ab76d8678129417dcd567344e4c7f71e0bb9f28b4025bf867d12f858ce0dad1f80c2410127afaa159112176;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h887f0024d8e28be2be06f778df25b17f61f82093aa5755e31afd2256e1331b592fea6975684cc7ac9e0a38d08cfa80138874;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h855cd7d1142215202d08e62b920d069bea9178c33f4746191c25456424a494778b8f0ea6121085f078512de91aae73df362a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64bae0141a212db434b873cca5c6c89e2e794b20e28ac4fa579a37f4a3e58686aa6f36133c4564fe9cff217fad026b4e2994;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f14c101e000f3f3eac94e1265d7f8123b260116501ed72f4b76cd6912de6f1a7ef8a0112b7e334e8d4bfc492217ce8c5dde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b488fdfa43597f2b82daf6f1423902111de909283a5897bb5bb73894f59615a102c1fb05a8ab6555391ff9161bb76d70a04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86bc1898751471ed40a2828cbb91acffe62a9619689e4f9fbde2d2db009ca9458867c33aee6a33ad8bb6ae1a53e313e62706;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3392404c73220187e5d64697dd5c4d980f3df892ef7653fc95ba1a0428f5b9a345a1e2439525b090f25807d58c485accad6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3747e45aaa195dd6aa99ac46d361be9cb23155fb4cf2b80542dcbecf05f7219ab86e6ba4e329e40b8bd92fa7a114f482bda4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96108ffa77518c1906557353e125e717d0a6f4edd91dbbb61310e17be7d6b58bc91c7e49f7cb795cf4c0564d7a1f8cf0a108;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3eb290028e195e31f3bb63ef945205a491048d7746ffc352370db72bcd9822f2e5114fd9a84e342760f6d6483cc51d44b4a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h481151971f699627ca255739409d59547d8543ff0e5d3330fe19691a3f5a3d829bfbca40181fa5b68621c4e92c7f3a703b83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81f9fd1a912c4672af3cb79dfba90403db593139bdbc06352c5eb6dc7769fab6d9fe7ca3f7e1d95445f0d010d7bea67a9ea5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h607b8764d90fd7583fbab2d22cb6d18d533c1f2b4371d821444b1b36ac181f10b9355ce47fc6cea322bd545a7dd6ab3d7da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb256039d6732aa18b1cc383ccfd29c612373c4e1d2b7fc67109ab02c2933192b1719c7571ebb4fc2065d9f00aa486dea8372;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha890f91dbccb9d91aa8c827ab324ba9d556cfb32b4056f485b40a981cc1d18ffbdbb9af7b66f5bf89fb204f2121bb313c329;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52cfc866f0eabba9d7000f952140d1439dc6a08f8a732806020c519a81e12eeaec3b64a7534643a247d35f6bd034422411e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbcceac5ffee32a761aa0de266d68e88647eb441ec326c16d471d77ac63e0b2553785037c1f6109a782a96e9a14e38bf1074;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6daa397503ad7826201da4f65c1be04eefa9b7402d53edb3538cd3450b8436142cfbe18bd0202efe86dc9b9468f3819d093;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd47243e421abf4341c62b05f8a4e47ca9be5e4682cb0b51fa1233e986e94d8f8c793755f1f6569ca5de98913fc0971d766c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d76468f759a97c55a145b8e299d1aaa0a0a890cde68e73d5d685dfc76d6ce40c03643df72a704103058cd9efbc81c25dd3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16bc1959e07515625bb72ffa4a4569b9d268bc58a46abbaf2c7d54e8f74bfa619ebe706735fa5c3fa34a5e4b09efce3b084d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62e6be4bcb323d5ab4e19929dd2d368873a58e444f89d4c4c01f7a8473dedc07db85cf4a488d526e0461193f4269495f7043;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62d21e3167dcc76e61a46411d7cd3590100c32223ff6a84b8892b1d884ed40e32309f3f9ba0b76d1e22cac78a644512f8c90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87e6d117a92e787d8d9bf72cc01b6682de5d63a685f171e7b347b847db5e67f934f627342f52822601f15f4cb58b51ab36fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7babd3ffd9027db6dfb9589bcaf1322be483c5caf5965fd717e86da1d1e7955bafe9d369bb7a919b663c5a46c6b4adcc311;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5831a52355d1c4d5ead92a90db92fe670eed1f3d5728ea55a38a89a3fdb2529cf9a1f5687b6bdbcdb6f3a71844c7e7d00f13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40d76af511c08fe2dd50d8fed526a8609eeec88fbd65339d87e4692b47b6ae730101bbac088965a227771ef5b80270ad6cf4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8b4652992d14fa53c62ca811e99600337d5f2285c443ab05f38650989cb82710bd1afd96e51a132cdffe5b43bde796c641;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a77aad87b2cb2bdff8a0d366f85e51c8fd653e021e5d0627745287bad03f570be33aad5aff2ae59f1d1078b6bf861a01506;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h985de54ae87f164554c4fe4933e7eb4e688e9d96dba9b0b9dd5d3d1c3a9a7532d79a996ce75bf9c1ccbc11f8e6293c34ad37;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c60759051910e7b491097ef6465872aedf3c6fc062fc07acc008c100ed96f894b2f0c5542b1f770f16109866047dc7d6213;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc6ca0043d0aadd18892272d99454825a52b494f111b281a80d739770672f7a0d67db71ba7f22f947b31d94bd09cb48091b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heca71334df754e80df97bc5dc119d5a13ed9cf9536af551300d5999f1f16a14732adb4507a9c62b4f9045d5caacf4065ccb8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdba8de0499487d4e1188b2e147c37189fa55013cb0375a660ec8d58c98d5be91cc6554585abf21607828ff0bb78a68b51e7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27f3ed2ee80a78b9c539562224f96cc1b5734d2c00b87dff84c130031564711fef3a6b9f0056a5cdf11bbb399ddab97f515f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ce5bfe76b75bee9262843ac36c2f74a8ccd834d49e2d4c04dcdc2e9775531f479acb409566cd79b679cb6413ad51d5c9bc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5f3b6540eac039c7ebf4fd2226afbe99356fc36a247de42afbf881912fffee001509afa2a5f81628ae9188109cc9a0351bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ce0001e2481c28a3ec7ece1659f48d44d328c702963b29dae9746f14ddfb3dd8306a0c150ed13c8212134cf6c8c2a96a7b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c3536edfa6e4750dc438626c22c189577d63bb08ff72190d3023b6dd14d5d9ef613d1d48ffbe3edc46c722e1dcec5fbca65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda59ffeb640dad63f11dea0fb073a5ce2a496c6313adc521d52ad73becc672551f81622f0603680d0119d6849e38dcb73f8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb784e774aca879b58b909f2c3bf8afb5939684eaf36d73351a38af7d3941612b8074da393adb6ddfb7204d0a89fcd06a8c7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f3b78878c15b85f2c701bca24b3e0ba52f06de21b9f679d9e7a7df7e3a4c7fd77ca53c1e8c38d67321d3e796878c33a462d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h167023103689ebde6ed16c092448368d97a671dc900d79b04ab09a6d12c4622d3ae811f0bdf71a0f4987ed96c85b12853a77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93457bb18d7e5a58473bff0c729da657a63f6aa005b79aece0371941afb8ca2c48d8ab58ccf81348dd38254c62cb0c062aaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h916cc5e806216bf8d276bf2440407d4e9d8603dd852b2b59b6fff3e1b99dea5e8227fb1ac4812010fdd29af1b0007ee22082;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a818db61709835204566054fa3debb05fba3759eea9d5cec18ef8411c50d2ca9054526def1d0ee9293e0147122c3667057f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c3b5772a617649f26f3c7ae0d7622e8c76283f39751ff4bdffde710a1d2c51cdf8cec42be345af5ec379af92c2e7da70d67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h110171da464bc32be4b94ad14b7a2ee6a18ae080fd964087d78fe9e6946ae32b680974120ddf15ce9a169f834f76478df6f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfae0b19cb60dfe492a45062b202a106e4772b599ce92e0570c6f4fa937c379b5abd5d83bd184b6b21802101d15dd6cba7954;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha912e9ea3bc690265282077ffd8b1de63c0d342c4145a743a2e78157f6a3f63f395cc2a28be9aec9c0214b1d130732f034c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36991d99384f16d56e9276dd22033f03b2a20eea64c0844cf37fc35de96ce1be1765377f1524040aa2dc973bab28962e26bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98b9b5a0b4d976b0eb08e933effca5228ad953bb6df767c753b41693e4b32db9dccdca7b9f21162c21c6a60493c038fa6467;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7576adf88bc992bd0005b1ca57edd8ff051f3d7543b27fa1104056391a0e3be954f6612dbde7d98789b73f36c5ee2a637970;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81d6c5ae44da83ab63f0af8a4e4353a2f27249e84665d2fa6d415f052bfc2bde992f6e57d17cbc7b21dc22f4c24a91256771;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h905a958dbc22c6654e9a6b8e1833d2e421bdd820cb78a0c0d2484fc3097a69121682c0f6af6007fdedc3dd134c1638bffb53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffcdd6562c30b9cf31b13b697e7c4acf5b25810e99391587e3b29242802b31e890cf37c689c4916e29b850f96e5b62c255ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a2a9f6262149a1b069564a03ce578aece1ad424d6f3f55a71f56d2ad21607f3196f7f9490887ca82738b17aa209dd496c39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6948490eb9417e90b3f3c213f42e204af3c631fbb722031be2386d2864d9798d728c3300953445a93080971a84f9049373f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dc31af5d8eec9b27c6b4395ee482e81ca7702d8e50b3f9f053735063ddb6b165e59ab322f409c0413fa7ffabea1a236c5f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd63125cc99bb7ed7a67963c96dc8cd719f16253e76ee90f25b3dda7122d73716ef6271bc0168757b803d868fbe9106d70994;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed746119cc78dbf49aca575ad8d965c99977156b40c7d2dbec7a85267571893c5ede2d3debd0f682ab3aa81c0405d4e77a15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h652f32fcbe930ed8cb1b39957e33582093d9cf1eff70e8abdea9ac7a4585f2e4d01bed53d9daf5518a26370a2b2a33f11fd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa96033faf92e927257d0f470ef5a74cca96d89707e4d3aada93d0c2b4ab7c3e6bf614ffd28642c5019d960f35996932392a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h860315b60629291d2ba8f1d2bad331058b0514002b1a2a58887a1b783b5ce0cefe806bcac1ec941519bb4e8b4bb87ba2c35a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha47e4845e5a930759e4df9a05b047cb2f965a95bb277fe31784406572023053774a3d97183de028ecbe99d642ce22e992991;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb342f2dca6b699cea936a8c39c96cd286f62b1935f84fae6a7aae62c641061b68738653e102dc3dad63186c15cf064bc25fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e44c0c48c226f4f7435ac3e9642e17e43992d4133dc306d27ea8136085a985a562d63da937d77a6a71342b0aaebfba23991;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e4c631d8cb5c3a82e24bf781883c3f856a801783ab005bbd3eecf2a9aff4fcd734c84ec9da1a965ad1d7086ef117909884a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h165232a7d582328b9d5a2a6975b39cc9efbb1466041ec00aaa1aee177d744709026da6f5ba122209df6194261745f3322e02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hace92a479ef436feff3463dd2a1082da2d5bfab503579f66f9e2eb03429386be223be498077a701510e2b4ee9cb88781a599;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ce88655f7a4b6c83a88fb4a6ac664c5145df5b47644d519ad661cbed24cb400ea496e3db4a9c5eb60b39213c96b137b727e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47e9fc9f2a50777285f5c93175bca36429b48315cbe0414626140b3fc23eb1984801b6eaeb353b9a95bce1ecc7003e9b1a15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d7935be6bcee62e7a598980d27b98b89ae28ce71779cbf12d6641767b468d992980b5ba4dbf6bdfa930829874e785bbbd6d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6e0615e7a73162a74c2120833d8d67e6a5ff04882070646e66bac7af7cbd6efa8b0805d327ef000d93f26205f8e682b41eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9f9c4899e004b1bb72c2a1c0617db2cdfa0aea58466e8f1e589bd28629deb36a9b1ac109be93baee4664925d031b499ef27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4f71b87efacb0e4873befef73a11ffb0e07a8f22c302bd3d63c5f4a760794a0df442297c71ea478fc2e09618d9f18f377ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94f0bebc8264adb3a413018ba7b2a3b41b33cb0f47c1cbfb80cfbdee28b908b083b2121644adfefd35604e8155cf74425641;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb78492e2836b59edef8a0ccee7b65a904a832a198ac5beecbb8fa8fabf13c10505954bdb4b33e56c67f572a7b061888eeda7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b93195a384977f3ce1b5ac2e6f47a57d6ea091beda9d960ac3873f9211344682b28408a741299ef20dc6ac341da5b9fc41f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ffed8fca35d170e4b4070484833194044c647ef03974e907ea5ce8375322c49d7b19e85a013d356150e8d35b8fbb5e7e088;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1466b29071d391f904a8612f19ff72329f4b76ce111e16ec41dcd52a2dfa07b3eeb7f723b00b0fb103d2b671f7dc4ef05851;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h282dd7cb45466b27029dd3224bb7399f46f3b0346ca3f3ecd9c8103145777b7d4bf33b89c6a8e6e01964eee3d504f845f46c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5cd8915dcf28f1e12558093871a4a8e37bc3da2cdf26f72117de40b5e997064eff96c894c56967c60103982457fbd831df8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66436cabbfb1ffb8349fd6473f465e995bae4cc1503f1ee9b42308c990415ed8139c96373ab7f9061ade8a51782025a1db63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f8e8ad64cedcd75910cd99e45a43a51cac5db50ae4eea38bf844274582c772b9383426021f19f4deb347dd7583e525555ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2d59658457802a16f63af14423287fce8babbd176d05e1d33fae9312ba53856e4858e6c4f88d5217f454dbe5083dd6ea215;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcadc5b13e4b33fc3c7fdffe65704aabe476b9f13e95b5432380b36d08bf783c44870500ee8fce266d4ddaba8ae541cdd92d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f0cf68072ad21ed213ea23c85853b497936c7dd4a5862cc3beaef3233b18d1a68b417449978aa7b45a9cbce8736f4a985e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb05e4ab5fdab19d7f032904676db22f0f4d828d4e05855636b35d8ca29e3c755680f4baeecffde5a160069eef463108ed379;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha86d01470f6629c2c47f5895b8cdad208e0c6dd76990301bb8e8c1a7beba02b101d6e7fff7eb428305575dc059fba9974407;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d16367ba324a278a346905ae06162f6a4786bdb9cb0cabbb6059fcae72aeba7a0179fb0e611964e53af065df291c2555ece;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf07dd865409eebc461959bcb0a862cf7574ad0e994d8fb1adadb9e6fc6fa60238a325c0d592f6af0f434d2532c3e22f8c021;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e94f534f37bb3f6970d367ec0d09944bdeb7d9eb352719bc17f742b9606b8d442895410210f320008315a37f4b754ed7575;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb850a8f32aa3fce33955f890e840b8873c61ecc6ffc92fee87b1a6b08cabffef206acbd1d1e64b7ef9c13ebad61c978f0614;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4baad86ac874fca07e05bbae7fe33bcb0dfd8638030f7e9133b0ae11364400a4c857918f055921af5f5dd817361803cb6bae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2728804ec39051fba2635d3176d67482b040415ae6d64024259655553ddb9a736aed1a6f3e5220726cddf6a73f12df69dbfc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he53bc484234696056d585f3d7d4c997c1cfa3416e622314522d91b0d4f6546f4463f0a79c819ee21e7cfad5da8ed18a7ab2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h444500ca8f77f3e9a54fd62775de0ec61d991be85a977e36fc8cfd572b3ff510a05ded320cd51bb6a2e241a190ebd700f48e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedfed8002094a2cce43900c30bb9316b0db4ed7e03bf81cdb1bb3da5d26330be6bc8d125b7facd8c53963868441df80e9e0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b2751668d04bf3f5de612af416ab21800409a3a06ad674dfae13144dec692cfe357299892a068e06855a3b715f3cefd8558;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a4af9bf9487c095168c7b64b9baf425d665a737bd6a64948f18e19a411903992a5839c7395a4a3bf2d10847e3be88086b6d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93d334bce3fde78a468326802f2800b8a18bff59add5fb7c59430fe6b271531ba3e29b77afe0b248062459afa13552caac26;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38c2c9b6a3fb19aa30aa3e1122754391ae4c43050a2b6e317062e5270c8b1afa9c3f8c084ee7ff79a6504cc583fdf9d2d9b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9423471d04bc0cdaa4a620e18a93a8e60803acd0567be496a41abdbe8276fb26f1855281fa06e647f89dfc06c49d9395d7f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81cfc78bcd01cb51acc5428788d00713c34e0eac06c3fa8af72ce438686404d628d230ededb2a589061c7df358cec4e23d9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94dc463a7965d9fd44e0d08566c20ef11bd80ffa8fcb89c19840030fc96d5b53c305e97f631f65ec4de0eaf55fc269ad0479;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h373f123a36e5fa8639d29f2bb55e12c688a96e8a785efeb8fb32ac7d477405257b923b9a8bb5732843b9dfe6422a8f5a4da4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd60df8b2bcbccf20c1f139ff112fa402dcd53ef20c43c3f7b91e51a07083a013b1eab8a3e63aeef55293236eb23e37ceb64d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6368dd9b0061a9326b4eb58e93328eb9936aeb1acb59c198eb1199dea060aadc76430e02fa9910e6168567db3e35839e6fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0580b931cc29010b713b50544aaa507be964570b6d17538f74b6fe350a9bda952a31e54e6452e276af659f03a6d9575f7b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h966c8eab509de48c1e7dacb8cbd616816ddc14f0f28430650d9db705558eae2c4c841bbbdff1cf8798aabfa171175d2a145c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a439c6fa36e963fdd614a68b0af0fd36f40f3ac388179074ed1f71a620cabf17d6b9f7efd4dd99a14f7b0d9815bc290ba0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ceb7e0f73c2ebf25911b290c7c10653fa4f4783f69416361f77113b493f889d6176c20498920264390c61ac5deeb021551f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52466ded233d55ff05efa684f78f96ba3074a8593667f2a0ae2ea0e0cf2121c7052d8488340972e5f46053d2e54f71d01f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d0a0933898e4d10da6c19437434ca8429bdf4ad1eee1d29e288978acef51384d08023dfc40cae28d95eda8e8ab4501977a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37df0812a2ff98bae345d26bb8732f02e5cb6a5c34d2af62a16861d6c53cd0804850a89a74e99bfce5b24508028ceaf34944;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ccf2994be48e46ad793508fcde27d0dfffd58add8994701345b6006efdc4a2c444865a2ae81db4bc65ed806f8cdf3b086e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90e5a309992aecf8521d09a6dccaca02e5c8e0e9de43794b251bfca187a493ce3adff505d8559c2a100f026b66aea9768717;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc58ecec0ce6e8cdc7d9829baf5a38738460f0fb56a81298406f8ffcd96bfd9bcd20e5b9bcef7bff6990493de3a05d7eeaf5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd73155a0164629bc231d5c171befc894946c9787b167e88d681431d5c86af011e38f2a16a511ff56d4fcefd068b5202f0681;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8826d75a0744e64009d0f445477be061a047f06849153690ffd0261239f3cf3a8d8e0fe31da389a1a2e507683bcc7fb9835;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h206138aa898e03e20e7cf5a15739edaf2c5599c7c0d3e75237e7bc9eeafbb01b6fae793ce3ee26ff31eff63720faedfc464;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28bdb1fe0118caa837f5f9c72151f51bdad94d8533462a042518f5c3d2424926114a38f3f78ba42e144916ce915c73e5f246;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab8edaf3557a2029275bafb499db719419edd6dac478d101021ada4313c11aa7eb356e27c8d438d95fb1d35981b995f23cbf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he131e9a3867089460f857f0cc4d6f3dffb8abeb55d15c628c674364d6fea97e0576a42668b0c7fb7260dc6eaafc1093a3f77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b16ac35cd169b126d3e8515f80913f28c396ed7214f38f14750e2e80f4d8bb9f047a550e1eb00454586df212cdbde23ac52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4596b814f8d75c72a4407c88aab0402d0994db814573268612a63909e0456e8c6b2aa37e1d91b19f2f0a992dba4e9e8281b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h604e8eec54ff1cab79abd216d8f32b4645916662724b9e46f95916a3bf20758ae3f9f767cd8a005907ec68c743f6c01d0077;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c8305ffa1b1878b61f6b363b374c72dab4a9cf9a11a732cdc3e74a06be0c814c504df0f2e059158a58654c73c5b0a2b600d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f94200023a40b7ebb8ad2318e6e94c1b185eb575b340f42b23466e241eb4ae813f0b8fea623fde1b25dae713d49e2c0736f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he62b0ddd69f2e6f082c275d83a1c3bb8642388ae07970248d7fbbd446cde146f7924f235dfaef70e8963256e0eedb13f24f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e6c096bc1437681e7ed03862fee9834c25a57561d540e604ab9be403e1239c28d23dd00652950923b987e11ae6a8c749348;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c116ae0b7276296d4d8f0473e7f2e81fbaa53940b37f868cbfa5e8bb4ac33c1d5116e17100824d7252b4ecd50ae484380a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc25660f142948bbcc5308aacc5b96dcd24ff782e894cd21c8df472f6dc0171bf49ac8a38bdc394dc478b9d4e34abcb82d4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61b273218b78d47e2c063458e3bc69b37366878d68728d1de645f242dbf67a44f146f2fa5ba4c2fcbd14d10026155a81c25f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf999527c9d46127cce845418e06329cb2019c71be0e3301625f008b917d3fdbd6ac72f9661ab944b95dbd705e6bfdfc25e09;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h725a88ecbcc66a02c4fb6509b5713e9a5f71e09ebb743cb373dd814e184872969fcb412c66d1db5aaf5aedfdb123749e70e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e72dfe70d2d61f193bcdfbe2755b821d3ab68df8a1f9c537671620fc2270d864a7602dfebe9ad984cee18dc78ed36d18e5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9133193d375edb0546db42ded22a4efdfe32dab25100a43e0354b4956e06b296007483bde1c20aa1aea58f76db09916295d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86c64ff792ffd633d611f41f166ec610f94a24626f5d324e42668e1ea2816018629c00358119e0270b2d408b28dbacdb2b4c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd527ab38daa3874c8b7e576cf8bc0cc26061505632cb8123c339cb500e57472dd52034f76c9a944fbd135dd90d6817690415;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a9f2d5e607206ac6f87baf7b73b0ad665202cd6c3fa83cd4d183d32d3ce88316c232cf9829fe948abac2f3d3bdac54fe5a4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd05fe8046a711d07b9127605d9003f3ff4a2bc6f77c395491a9ba8b1021b8634c8e1b68c91c9c96938776b4443722f0af385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd558fcbff04f225d0eeb6a042a492fa44fb09aab35e8259a23bf570811277cde54b0206dd83035fc62172094aa8c64b7c4a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62ff1a6a68c6b9de035f82b11e6ef2b9fa1ff6edcbfc0b0a39272989f8a94de849a4b10f208e58caa2bcea17f70dc7c38b4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcf4f33de35fde53d12895e0bdb1939b200ad02476123b2de59390a1107c35f52eac92013d6391dc4523ee2eb1b3107bf204;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h537a056ad20e2fc83ae8706e56e34b9082abd36de1f9cd8010a753ff88cd46c5a619b26dba921e0a1fb2b34035832dc33dec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2b2753e0c8964368270d76d11c56392585f4d8833d208111d25acca5420ef79f0c80f9b0d432b142d8dc2403e7617bbcc3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h541005cdb3c2ac1e933e3d60925c280d77f2eb233285efe507cfa05b79428fdf6f55f2985a57fdcf55147144ae0441e03d5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68959e9f60181ac45e23764cd0424db26572c49c8a0b8a03e5a9f5a87ec8ec760196e05c9bf4b133196c37f006e109fd7b84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe7192fb9646be7851bdf62026441570a43ca64edd54007dc409d11906d011666c8d2493b1b2b8e2e570b5274bf9219d47bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h378021b75dd992a3cea0651db7a9686594e55a4d2a2902b786b59a697ed68e65182ab7773a3a974ad79d89906320249d4894;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf28995deca6361d96f6d21984f5f8d7be9166beabcb270687315baab90c4144665c43a6900ac6421d9c873e818b15dce43ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b36ef5c7413d871af46f1e42d831fedd8febb3f7e2514dec94b89d425816bbc6ffedafc34bf70a966ec7c240d73e9fd3d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8eed20b531a7dbde9f00369b184f11b7c5763355bbff0fd33331a4b9b28838c8c3f49db75e4c92e13dc4abdda2da33202bfc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd02c95d2bcd22a83de7e18a677b4aac044e808920ec548815c615b505b31fb981292542e009c2aa63657cf5e56ba2831dc57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h738f832faf6a5d6fc45cd30e03c856aa602b17e898f6edd88b8f8278adef693943d2dfdc25ba52d527a23a13d391ba1e7296;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf84246770227f758b54ba9f1e963d700d46ad19dd37214c53633a12f629afd054675e68150ddc7c087c677b4a27003fadc3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3310e6d773ed42a6c78349d56c02b73ce9cbb2684cc0b2f000e6a83c5a025dab1fbf85c5a1e2b9653b81d535f0096e1005a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7946a13dc5bebb70fabbe8439e51c28464e2b636711777298cd3949ed3d7f905bd25c064f0fe6a9aabeca2e5be0e53fdf8ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h116eddbf571ca7b372f52e6050a1c2f72e65b6dd53d1b27b03f9491a1886636491bca8113fab234c51ed1fe31f66b10922c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h476053dd3a037d18b3886e9b757133022c2d2dad20fc784694acbd3255d74b6c9dfb6842a8ace1c25f4b4d71cc39ab1cac2c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h209da4821ff106d7d763665acc52f188b8bace4e95f923ed652aaf21c1c510ba81724e5c1b09a61bda5ce6e434b6b3e4766d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba21071fc2aaac61d38e81ef7401e9bc77c2b6c2f675529ce96cf491a576d68fcb5ab0f6adf4ff36e682fad02274fa164500;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36ca78a6b5d824937296beb9637740f78ccb41532259400186f2c17f353758b76fa3a679fe7d3e1e48fb61a7227a533ad5f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha70917ba8d9db7fed89a6d0aa20de05b33e1ca48bfb2184fc5cdbede99cf0c02e5563199cc3042e259ea0a8b9c13542b4fba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4af9f43703fcbcb9c2e37dab42ba918cc1be6e9b79aa3935adefa34c227f97602fa0a9848b3d35c9d14001cc3540f08822f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe467f07307e6b9a706196536c37339c719836c337a9e7a4a2e537420e827960b746d0c4c175590c8a49a6e2ff329c24a835;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fd0964619743ee14e8bf4cc789f2868e02cdec0c65e487995933ed3d17e59c86d8e33216db7f99d71695a444920f53c7133;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47ebfd773b62f6951eaf71e69e3becae1ed63d44fca9697b75a4ada5ea42a004337bb178d74c869121c6b37d71a3a619bc5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ccbe64cca0da5cfac7ed5ed4db9cf80cfb8a84b10ec4aeefd49ca0dd8abd7f233eb5082e37651eb5595f3b145bb803a67f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec11e2b6eab8f1be8054b00463ab4582a0bb3b7014374fd4ac665870f85204a1abe1bf0ee4908dab2ad6c191662c1d3e14a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdab736e2fc48370b42c5ea5d2bf011a878d9569e976568ee55d1cb5b3108f15f203c2b31df7bf9d952e6a114e209974de68e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbb65f05dc1c7e16f464249c058651c64266e288c2911ceb2b2baf17f2b1cbb987681f5fa04ebb505b67079b9844cc40dc3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a94d0bb0b5438aac25e6252f6a650b3288069da2476e135be890749b0d0a5e03e6c3c30a7110b0c5c03ef7197fdd6bb5795;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e7f1f68eff451f9db8a263780b80004ec7559733a89063f1aac8d9c11675516384a1fb81a40f7d8eabd550bf5b60c3f53e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe290ca3286aad5bed9958e6ca8559fda22441741cec1dd5840662162462750651b97052fbfa58b9d1d23ac586b82910fe31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h433df0cde18e3ae1dab7127e04620b7823c565ef3377c54590e3ff1590bb9d47904bb7872c73a63e4d7aab7efc3f15e0a5c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a1b3b77ad32b8dad464dba2c885f10eaf18b71905951f67067818228fcd5c70b7702b2debebc7bf677d9fd1d3b7c706fa26;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h599a8b11240891047e921915c7b0a9455e6392e751ddfc4ae786eb27204530df801be593621a4c1f24cecd2cececab6d5bd3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6ac0c0eeb97b998adb68a1404a6fef3e530b356d9f0c9b0981c2d2e2ee81caae4294b8a1629289da13d8ce1c64ec12a4650;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91e8dd345bb75ca3f43f28d0702896d81151127d28da73073fbd2dd8a6932a188bab5b767667d42c5478fb311b0f21558d86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1595c71ac85e1b724d4b9533a92c0d1296012568562b07c24e8a47750db861efb530ef016f0667ae5b23401e248e05722c8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha83736a9bef0368a18ea530d3ae1131057ad2c9fed0bb02d7ecd9d4e9762a45ff459e4e71e7643565af734f5805668e24a6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38f89e7e7edbc16e414efa769682f2f3413b0cabd15c02cbe91e9afbdc4803e2860f72a9b03cca67c7f8539760f7ac4e2941;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19fb2fa1cad76ad8d13d5b8606c51e4da831c92eb25b53f51bb6945cd7940da2d88fcb2b8de1a34aa43088fba47efa63f8a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6491f5d203a0f8ae5fa16d962e7383c60f07e91f6eba8e947aef467731b59c65e8e0c7d277ea8d6f6cbfd4ce54e6a8222e3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d3797673e9497102071939934956990277767b3b9360fd8a066d30200f6f27a6f527a6b770fc9f33fcc386993ebcdff6ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0a14643de3bd91c945aeba88fe61f7da906a8975dd3bc126ed3e29a848706ceed29da7cc4879914a2b285ab8e41d2cc5333;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1313449bd1ec189217459c07be65f1dac50c3d498074233e43e11805a9c9a9f08fac8d3493615af7430812b400d04f1dbc43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd148e703382ace3d5bd66bc502ab78d6323fc02294b098de6cc1acd7edc7ac84c567b351bde864c70e1ade18fc5e9c3e329d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65ebc445a1584a89881ad2ff3bef4a64be50def6fcca060b7666fe8d9b27f3f3b7c38858e2027f7021d4f948f501b0ce13dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he065b30c070f00d71da63dfeb17eccafcfaa0d2ef769d433987713d84742b23d136c6da37a10991f9f318699b5fff773548e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0ed537aea1903373170c3339e34d206f130aa0a8c6a35ed408283b8b3e0018786febd09195009bd14657eb8823739ae2b59;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55b1ec30ac818468327d616d89d95c875663e8cd478a22bb85f527dcc54e5b0d365e24c8dacc135a2e220eb4dd4bd26ac0f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3392379254bd237c03ab7ea1389228abcdc7eff1b9d8a3703402a0276053b37cf2104b3d6e71f8f60fb89a3f0852fefc929;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4a9acc87cccbf8916a4090820c0968979779af252574897d6f2dc57d3be936cc8a205d36eec08ca0541efc6d5b55e20225a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a64d17637f2b616fbc457cbbc4f420268fed1a4171e2a1c9580fa28418e680edb028db3d74ac7639112267a7f14cda25d31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefc5e410da2f6cec87fd258c6779b67e65bdffd976fcf143373b1fa96a775fb5ebbc442e1e4c317c2e9219f632c3e1990ce5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fa0756ca653604bbfc1bd3008a2de44861d9f8ede47ee61f3819472195dad566c2c196db36d0ab128e04e7a1acfd30a7c67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1abe71ab5f0e512921521ae4e0dda392fcf5c8e23b60d583c21396cdc8b19438464ba62539496c375bbaeb94393753049534;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f85ac2b223061d7a564bb4d418315fbb6bed56604d289bdcce9108f4b8cdb90150e68aad5c000160a51215081cc6ab63d99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23df3c1938f490c3ef21ae98bd6f83f87fe8fa313a9b4e55a36cf3de6d1d9bdfbec84ecafc4a14328853ff4ae7a0a13597d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6551131947b5c84a69090b438b14b358cd28b100240fd0e31c786abc5fa6247573f6ba59d72f0944cfca56a590942500eb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a0c511ccfe54da37c4803f109d7b59a96dbe4c74414e76fe4563c2fd5e2ea6605b02d12d943eeae2b5b01dbd1aa158e9006;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d9e7e807726c473781f05ee2576b0a5a65f249cb1c6325fe733bbc93d04d7847d06d92248f9408481f11693aefcb43258c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h295f075ec46230c89de94ae120ea5491b6d1ad443a164088d14bcc905de50cc63591508993039713384f7579a1c9ca31eea0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e22336e3f6a29c73453a193594e1865f9d8bdf1e6c47598c401a99620852e9715f3c2c76eaa1d492080d32197da7ffba814;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4011efa592bcf582e43e6a5bac52e3a266f4929f55baf92f9b9b2237207d4ef9fafda3de9464665c234d2593046ca530e098;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2a789a18fe5b094edd2c5f307363b95b5dbc7f02fff47916c54b46af52e14180c90e1e8ecc37a0330e470eb761888c1afd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb837534566e75ae3bb9df1730cb2c04b23970d01e40cba5791f46e9800b7faf9ee667d65d8599c07d24464417033f0e430ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a6b55d2c963b3bccc5475893bfe2c696045abda99890f610ecc211beb80c6e6701bf0f570a8b305124dd237342090169f47;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96af016ae5e2b97414d877546a6b36915daf99c0d7917e4904e492a107320af7a0a8cef5de024699333db038627f6b922c5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6a80da634b165627c832f32f511e8283377373ab0137728c31a262dcea4bd5a6c9e0cf39fb4be28f03bc446164c6ac0e339;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9ce288cfcef74d4d3f1a1db4e0b46eadf995141eee3b73a3cd0c9fc0b366040569df7ea09ef7f608b96d11fa135cbc14e31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67e22297a06cfdd453a2bb546e9bd2a1ba04dca9ec5c5667ce241a4850967897974ae12bbbe9c9acec85c66ec61c1bab3c88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d1410648becdea552f89297991da29b17fb771010c7cbf4a87e880505ca215f83ea313a25a1dc4f0736b198b12bf381f9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5ccc187a9025512836fa425e7ab2334d203b4e15194c8fb73a910359717a735fc5760e6e701299e2d0c63bcc905cee34b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf47fef97d527e883e03c872e02e90abfda7b6443348d9ce9f500d5ba0d9d0f8840fcbc07bae007da0c1714f9acaedbdfb7dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50f86752c22e69179b5648e5e3ffbe1e49c5dd5849b920a3c99240bde3a46dd570e9ffec57f28d792e9f49b43a603ec8df66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h464fd5dc7e59a3436eabb2f4f0102fe7812c17841ea5e5562b4f3b19fc0f7218a58dd72308bff128f95a04c744c3847d7cff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59665b067c7fd2495915ec751ab3d810b29fb7bad7361c14a02b8d2c9a7e345f196cef15cd6cb4fb75a339f15914209ede8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521a53af2a8d25fefd154eede66ee2fafead8ad402a7498cd32104ad647b2f95f28df9834bacf61685d55555f8c6afbd0c94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heffd62b972a82d87f72344cffc125f76c8f6f8eb5e33d9040603f7f488f1a53a25e724e393629f82e32eda398a97e0398aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94ee3fe733e4d08de7f08dde994bba0a235298564791b8d9ebc582215651373e91dc5c52a746f11a31088a41cb08bdef8963;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9b5c5cc07b60165e1c0142eef817b5e4155e5f581f6233f0d8a4b1550823fe381f6c628973573902ac9f6a1666b1eafeb02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd070a9f38841e581f45f0965daa7cab27a906e22b39a1e74221bb7105384d5b97c710695825fffa31c9cc724cd4200231e81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd5e679f253fb69cdfd33211f6cd66bfe9edb12db5cc577624e3a55af19d6412f7fa8f60d026fb940817e9c7101fc350bc24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0a3822ecae98315b34fff26352eb3e6b20ad8f16cfecae0e1a0b95300b15686256975d7fbef801d5c18e931b9839df8d774;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd915e95305d81b6f77f5a957eb35099654a0f25aff0d9a05d528aca54a658b7341f32967dd0a74cf0f66d35c9523c45bbc86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68442e83db2ee7906c17952737ceffe03917ac9c4450bb703001a6e243c95f4826651d9de54a0ff93e8a315d9948a2c4cd89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd0b69727eb5f9ba22ac147b22dd1c0bfa5930614a202d8ef0ee82d0e87b5c5288c423c318d66e76b7cbcf27b152ac721015;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb60279d1bf31ff436b73c10368ca28ee1a321ed9aece05b7f6dba40d5aa85e20529f00bbd7d244b6e6c4758585a2fe9360;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a7c96b32e2a1b67fe586dcc6065aa7c97fed802f6e1f5121271b3008a69411b9e0a49d0453dcdaee5a86290760b548ba2d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98cb4f756827ac10af2337b91f485d1e59f00787e96c314d33559293e2b43ce00ccef0af4e4a36a4efc98972e6232dfa170b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3855e206d310e0936c1f0b5ea807498522f0d8be5031caf8a2014014b90628f6525af288826ef46908a3922092cf2f6985b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf81ee27cbf9f1d527750c2f02b1ebdd91c5c23c95a5d4aa4acd0f8764268fb9e2e8fa752b1e66fb556e70ea5d08393dcdc87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ba7b96aca53519e38e94eef6df1f952009fb03217e91fc649e01260e1b202e0eec1dab8e9d1b13b33603d9ce6a4f03fe360;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4ad0f11dce88f1cb9e497868b99033110c12972780fd804c199f34c560103dd0426476e3ac0144a883a206f8a3babe39a50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20be7cf51cbc573be4b06bef1d68f0caf8dcc8fe23d8eeb4493615cee8fc4e2ff129ce19f742258a910f22dc935ea7853779;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96ba2c678aad751035586c8aea6e84994dc691354b9feaa1e67a13d3e4a7b837b35ff47fc8c5124e089a982cf5ddd7736f58;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8634875e752a39030964c491fff8ab075712451debae9c758f91d50deecef49d25fe4ed9f26da61de12e8ab122d1aae783dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd99d00d50300df7f7413b459783f1bc55ea0d88080dc4b58f9c92585e4d8315cd127f7f2e06f5462f622e2a79083b169e53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35f1403608872e4ea8f5bc257a3266523740b015a36ef1d53fa907512ad306c842d8a13858edd3bf518a554bd1962467715b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41a79f9a20905afb090c15993886e6251f5cba3f2cc59dab01918db7377e113c375e64a4a0d400f4b33b48b93b1051ab569;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h792cc3012f5f1355b306862f80b2018d8b80d1cd94d188c8271fba4f62ed9112476ecc9ee521e7895c02115289b374ee15c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fdf94548c165f97e8d916cd96e5db37435d4c93fadc7b267353be7145bf0e036969f59b2ec30b614cb51e6d5f1bf1d5ee5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40acdbbc0245255afdebf25ccfd5f64e30b59091fbcfc0614d1a6718305d1fdee1d82bbc00919f0ebbbb5c84ac3e1de1bc8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6043b34374cf100f3c28617a9ea273332501189d0e15a21656272e1b39183a2f4619d403ebb9c320a38215d2a122ecc25be9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd87b14eed36324096405c717e2961207283748382ac42a2e4d8088a2eb83f123b634bcde0b5d0fcd1e23d16ebc03564c5be9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6e92f0c3ca8f7f94d88270791f7030922485f816e180371008debca344f9cb44e1fb99b043b0b473fdca69821ad346b3fa9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd84e13ec228c33a072fb708e69c12e674ba6464b51dcc0dad43f13c609dfb348120c9aff1532b6a596da0593c8003ecb9678;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64236d9e76e9bb5959c82270600054b3055647bd63da402138bc62e0da8ca20473feb7aae06a9419d2e1e6001add06f79e66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9b46b6abf93ad312cc420cedb649167d38a6bb4c36d4cc14813cc830ee396cc734105ea71098274e3c445c1aa36a0bebb53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e6b17afc1ec45ecd4b0263bfbf024376b76590b2b9cedb7409388ac4938b11e47564fc2c2e72b66a22acaf3d5480cda3d34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56cc94f534b3bad42c5bf2a6654360a03071216a2f4da963a7214d2fa1a01d434785170097f758dcc096bcc156b8069b64cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a136270dd1e38debc22b0487c8b48ab2a0acf065418873aec8df5819d6b2d4d2f7b9dc12eb5be4c0354fc90abd5d99be958;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bd55bffb1b682aebef02aac3859b9bd0d3d8ae182b210c811359c10ce98244b02feab72febc8af467ef6f9354e103c68b4c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c9ff47a3f6df83a60a101a8101988c2a3572daa0cf104c283c97ae5bd741edfc9a9e1677f70615bea7a20fe9090f9097f8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h113df4222da6d5902f893c6f40973fb5ac955a8662a5a416165f52ac771447b91316d65c1bf163e96fad6c8039027730395f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ceac15eee7ea4e787fa228f2bd049ed2fc27ec0a23403a96f3992ad0f327d68b18e5eed0e4b6b653eee5da12e749daaea4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bb28de354c8025b052616c2b7f17af22231d378c7210a3f57326871e6ef5d7b6568fa651cd36ed896c90a8d7d1c22a2b6ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h548b1177521fd381de394f3300c458d5fdad4625db5d3cadbb91edc33009c63cd69d273bdc6f54c9cc055fc4021e09b0aff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he64609d2173c60bd9ca748e7a5debaed7c35a68587f3463942880a0f4207669bb0c1713324322a83ec517091ff531a71bd8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb043d01a3bd9fc44b69ec67491c5adda3170dd01fb0a2ba2d2139606bbb2963453f0e2d3889c3668f0b79d32608cc0fec42b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc261c38dac777ee7c7a209ee57c4324afcb245b40c805eecc6589dff00c28d9ae5a8e59e3af9d5a79d28e36b26d8c4baa251;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he64503a4977337ebf0c517db072188c0ab0172a9eecbdaaae8ba7fcf822dc2baa5360986c785dd9f9a480f0c14188fd2879b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78438240cc62490669cab1001561f80b30ed0e20002330caf8ae8a3d5bcb94cfee43f5a145665e10d9a66316ce16e85ac0c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0a71662289e08ee7c4a1bb0561cc19d210d196b94e59c7588ece70c1a036fdd72be1723fc0d3937efe38161f0953f2cfc87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h742511836126b29d80b37154cd811ccbb0c5c714357b688340118c985ed2c4516de4bcc986fd832392a548511f61692e5e72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a12b44d04805a38f5ea6d198b3eff1ac1dda32216981d9840d27b3260bfd422f6f3f33a1c6d86b5a015bc982196254c9448;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd4cf2386a941f0d9622977c37a014a1046dd2d63c66de7ba1f6fc418c1878af8e2727b3d7b3ece9412bc253e56f21b89e73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2eb2be54e56d8028fc7fd0abd95cfeb3fce4726de3d3d79d9f290b6664f049039fe7fdbb714ae913a994ff0e234264012b2a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aa1f9e0b508f2d8bf57f8f8981ddc3cc824103c6b14bc6c93a646b6a3e48803e3feaec9542914de26af9287954878b7e057;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6854b4cb01347186b14121dc84481197c8437c5c3475ae38df0b574b953f09d65297402f7f2d819d4174533d11180d1b444;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e9b11ff10766fb0aa33f38435128695381e8ba39d7f4fb80678000d7055b675cdec8e87958eb6e4d4e74cb4d7c4ae354451;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88ff5f4ccd3ac7e91d640a901056a12cfe9aefe4f28ad8dc77deb73b1dcc4d9a875c728b1568b8092e660355bce005ea1af3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h598c6a3b94da4e8a21735bd0ea6420b185db450ba7ff19eee5df4f1fddf39c2e161ac439f91754a98e27c2c912d9f40e7c87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0e6a6266683e8701fd05ff8dd5ded17c63bb9a25d769cd3d8cf5354a161d831f9b9ca62504d1a3060cac0c2fcdad8decfec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee483f789c2382129650c904dca0d81d530aea26ef8652fb2f8fa37f22a3d29b56ca11a75b40d98b9630f011224213e90c60;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87f6eda9af1aaa8c775ba0bb2e35bb66eaeb3fa25ad576b578e2bddd6b41d27b10b76cd09c3c1b33937bb597f10f7782c29d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe3f98a61c48507c70e8747304306a0e19223fa3f6c6a3e8fb87d05fb88d31e7aaa9add25bf2b942512018a9ab15ded79bdb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he66571dea7a09e19dbc9a4772a8aa049b06124d91aeb732e37369218597b086fdcc4056713bea970e82c16a897034fcdc4d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2821362939dd48e24dc0f96eee310b5cc587c3302d7e687d478078df41160d59f33a938dc35bd6e59f65c53d3173e38a73e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5b6e123bdb068b5cf6bca4907f980131d2798ab90a71b16d4973f8ba02f120adedd9c34b8af9f198fa0b16c4e9437b9e261;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53c8140a20cfb64c6540110b639015b1f24f87ece192d4b3ef1b37be862b926ef7fdcb25117249759e2e21155c7e8f2ff072;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2f2beb1f0e214a8174d5ad77c6d71e27c31d13bc5bf287b6c40ec2dda6fceb7be7dbeb9498a75d5272437609c35dddebe8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcba7b7d815f28b0330e27936db5ca3e448f17532a89f281429e1d5bfd22560826bac1edd294384d62841c361ea88bd322665;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc888696a0f0cf319bf23accdd3d04529555e71b5035e530dfa85ad7f91ba759457fd146eb978d8cfcf48049f66e2fc9ed5b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f6bae9baf188050e8fcc6d8c0ae8660244f059fa9dd41d9434d1171fe769b3918579b99346f40da0cbf673b864cd2562fb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb43a72fff0003d3803629432237e122e0ed7791596eebd78d23142edebef49f94fef211fd94bcbf968f31c56bb920d8339d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc435cf53644bd087a02eaa419682ed4f77ec90cebd1a93f9f26dd310df2dfd674955f55fff969d49c1f8dfdf9b6140ffdda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96ac7742c2533ff16bbd8be3b779c7e89b710e423e122935b7d3d3c0c4238bb4eb696dbec776dccabad12227948e91e3761c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8a05f35bcb99fe10e0dd81e97d510eee7825d4ff4ad828470c29d29e2a7d6d5b2699fa98999799d853a9c64c866845e9851;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba8584a4829733f0763342f117fc2b86af62da0bb53ed6434219e78546d44dd8afa77a9fa1f567936f431c557abc135372bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8a783dcca4e39640c9c5cb2c607f70a7ff3e1fdc39bc54e97b7392483a65d3ae933c04aa570de0b308138725a0149350821;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he99d015f6ce8cb749a1db9318cf78701aaba11f99b9142ed10492bfaaaf412781408e034a4999719f43b68bb0f79b499463a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h965dabe0d0689662478fc0a3cd6eccce069eeada6d52e3a7e982a3b7e9f33d88efb4bd5e4f0358cfeb9abe5d3071f1798b20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e9c53fe9d30dd6c8101a4788af41d46e865d973c2bcddfdda705e8db5b8ea1264a095678f23678349332041409c0045aad7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73e051f418449a077806dc1a5860e3a94253b2750e97e832b221b1cd89dfbb87cb643c0b10fb92dfc19e272a7f7e3de117d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b354519686c986a3ebe0f5b53f3e8b85bb72ad975a6eb925016ca62eb2f636318c6e72f9b47412ed251ee74afb200a08d8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9b3e8d5cb18b7db7e813e33512b5f0e56730d194e33474ce6c51143711826173905fd027f1abaede8c2ec2c548671de3e29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he04ce3145e45ce9f094bafce857748819ebca0b4f6e5eadcd78517079ee06432a617cabc02f1629a76f259e59ddbfeec79b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a6c0fcd93a4b727db3dc6532006a9681a6c77a2c21fb2af82f25ca45e31baf9f9d44b0aed924ab3f5a860700a497b86869;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5cc2be01afd65268c11633da21f82c2d45eab2d4bd2c6c45bff99792315b9eb0c51b2ef73197c213daa8f32d00dab1d7927;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2a6173197e0b9f3fefa8718210c649555b8020fa6c5231864c81c86eabcec14f8dc0f9be5ab86602209f61121f289450fa6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2dbba12b71d88fdadc800ce61a7f2dcb6a86ba9d025878891433bf9a90824e6604da419b7e87a26cef261f31a86961e5911;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcdcf05b87d1d75a9c08f0219b61c964ca9cca4f721d26331b057c4c6dab00d65e9949e220f7ac47370af34398648eaca3c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2073ec2705edccfa62415b71af5994c7a6023a8bc0112e87af02b5b706877c2e570e8d9bd048f6f61cd11878e5904ce7cebf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2fee4a6eaba5b3225b70351ad96988ef03c6abffaeaba6b5ab2afce3479ee45017ce89259075887a7e2a4b77453591fbe7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd086d35e6b8e996ed04dfbff9048db6185ef0877fa1f3aceeebc93b391b1cce5689664124179446350dc3abd085dec3c1b7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb31414a7a974bd8e62c43f6888e11fc32452bf5669bd5e8999aadefc0981097bd7c2143578d064c34a5e0469a804a4faee1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h674aa1bddbeea5581ef911190fa376578f1766f6491efef22a1d4b5d3131ff32ebc9e7a79cbbdeab3b03d7ac1b12e29c358e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83d4f83cb754e6231a2dbabfd7875a620efd94f67a3516fbd963de6639ae5b89923073f26441d6a94b79673e1730130e2916;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6927247e999c98772c35fb0b7cd05fbed788a72d441448c904bc15ab354e8b845354b0f2614585c0365108911e87718534;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h428d15de1260195c5363518b70ba33169d9fbc2c520486364b5b278984929e2ec6643a25c3624d67955cf664927ea7ae1eaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h387ac90f4fbafad15a8ee95f81e5de88c27ce0891ef413bd7c5bac1fb541bdd23cb80f8ec721a39129e4598a10b68f2d12b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bf7c933550c390211604e98cfd52bc65953b59e00898e3f45a31e2f9fa0be1b949b624d3498380bf9ca4811eb30f5026f4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7239198f015b02bfa1b4e060a02dcfdc75ca0871bfa5fdfb7831b3bf1f319a9a3fd9b60973dc6ffefb4e49ba641d6e5b9ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a31d8f6a841d1d433d7e858684a7511ef7497d4409dcecdba4be7bfbf94c3e2d94248d00681ab29c27a66c78f59a3bdd644;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h930fb1f5501709e33ef21bbe5795c32c654cec6a800584f59f8e024548b75e939a277c8ca31d9ac9d665e45138b0ff6f314d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0bd838b22c1db2c96cc59a4cb755211241515bcec460f2a6d30b24f8da83dcb9b554778236b7b33e720ab38bca32d94312a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h937859b5240120626782bc903b5f9f7ff6ebc6dd533ac02bab1410eba54f2da3aa141b40c80dc5915c725c8396547765920b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd54dc299c37391f6805fea5198e4079c9d48452560cfc76aa8011f3fc7a8eeb80daa9a073dcab8454fd5b8cb08ce9f215ae7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33598a1fd4243d230da5d3e962357eff028cabf508c0bca63a0794bcf2b1291f0b24a9b69eff7df710212424291bc76400bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d96b44210b461999a7cf8a62e9007ec7321eb36a588b6a6c728e3325032a6edce61a0f5e4e0ae1a348c59546d675a360519;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e24b8f2f6311e488b47c55f9e1e657f2e3cb033f09c85e8acb95fc28db87edf8a92fc2799fc5f9ad98db5391274909f2069;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68f3a6fb99d65816ea8005c3da9fae324d4f3a191c2867a2a9282ed17fbbcad30000e83dd9b2e0fd3693c776517fae575ebc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he383131e4866c0dff609f8a1e7f8794e779bc630453c415856a2c3d557475358d7b78079997007cd3cd3c232e6f05f2035b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb551b3eefa364d04c0ca7930a6a4d2a8e453d63146cbb64621947618b7b7b8453c8f76092959856391bd2a901f394c24b22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcd6217803db0f65d3f16ffc43babcc9fb491b9efba2e71fd2b7566f1b98fdf0d4f7317c4e9bf98b3da55c59ae33e6660f90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25d898e4538187812b5366beaa66cf04cc6e6946bc8639878ead2aa9ca73612b8b547086edab415cf74f0d6e30d4a705acfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50e3f053bff7756ad789502f68e2ded8ae9d7d69ffee0257072a319ed828c29d7c080b228413a3f7f22aa174bd4fb8ee2a70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf27d3f9b21f97595aca884745e58c871e87f5c77458ce80b6131da251a8dfab4eeeda822b489c94824b207355d8aecf4d9f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd105f2e0644b14c5d85352c8b6df80329d63d4b485efe01e5618b21fe7a2fd31c038aa70201855c5172c7785b24573f885de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2edb5308552844ca94f2a258d8816a7d4a7d6d36be45c13b5900dc5e81b0dd4391cd8f1e5fc86b445223fa2841c7a4123c03;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h542b6413a78f4c39fdf94ef126e55ce28aed48db4a1f1e0b3ba4d62aeff9409b46f3233bef1b255fcd04816b30708eec03f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha762425e1ff8a8a2e537fb0ca2194c8950bdc86267fb5841df769d4bd35199d58775eb3a234bb5c2d3de8e5b42885535cf21;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1820977c90525f0833d557dbab25dd86a81234ea2212eca27ea5e026a26a4cbd87e83e488a8158c83f84078520bdcebfac66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5de46b4f998bef5435d66549b3c65db7c3598bbbfda0ce90f77d0bd1cb7e7c271ba2d63d495618aeab3d52eb1681a78c8806;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62ab70cfff4a936b48fd5de47fee25eeece840b76933fc3d9f964187b1e081f5695a227d40570c4c88f2890c0e5132ed6e08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he30ebdb10e5275ed54221b7983d590b630fe6e1452c86370423a16f8042a910bacbded8f71682cf9d43c43f7f4a4bfc0811f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h990f1eb103f5bd78b4c8a2fc0b16d3c65a6c66bc58cb3b25e36fa9f986f99133c0e298d9188787c642cf59202ed1f4862adc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb8c55e0275e655f7f4e5042e127caa02494a61930b2cec244e69dd274794a1e1aabf2ad19c499312aba98e80ea264d93100;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ceab3ad460d22c48725b027dfca5a9de4d5f9a765ebf7e42facf5d9b249a8e991f43b8aed5b6a72b3ea09ad836da9844135;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb5facc2f95c18a8d8d53a3b1136be94897a6f2da6fe7376ee7b49eed2c7751c6e0919a9b35cb7b8b85c297a484e6c8b2ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h128d45b79070727cf40fec08f71731b58b9fdb266e9941e85f2339975688a740947bb848a2fce31b0089dcfa5c3aa08217d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h920f2b36bbc0d354948ebb7f37957869972fd1865dca2503975c7b79b111514d0deddff3fd7d5164f8c4412fd239a79941d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3fd3bc4e86fd70a2116cac2ff4a80f8edbb8518210138862004c34e98c4ef8d76171b8093c8fede7125802755e9d4b45577;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66dca7d0a059305aa1b192a79bd6ab23191e9f094f4201804057bbebea69d2e610b08395f7b6e281779390732174ebbd53b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcff9c089ae5db6579feb3e787c80591a054fbc9e9298a14e89f1e508a875c226c4b671d2591ef77e640e1a723a2dbc84adc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5cf02fc9b28961ef9084c6922e945330831614f601deed61a988ae560db513d36bfb775794495ee6919107a56eb696e4efb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d25f8905eda2a79a197a1e00cc4a1d19c1a0b089245b00be97184f63b25fa234de8881ec8b72dd3926f1fc328a0d6a70951;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee79e53ae86b54b48a9f391fbf07a5f8dab3c65c7fa487f3c567483f97ffb1a186a8597884d62889938a9888561b1d83fe09;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f9b9401c7c73620e33553f2de85c4564334baf2d01fd54f32b7470b53e4e51eb3a19ef80ad93014222b4438f17e08d1aec6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68e787df983e8b32645c74a5bfb78e9d356f6275a8d1800aa3b884a309802d6df9d29c781d5ddc81b1f87d31f0f4f983209;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e302181c1e3d3b5a887898a50e8456bef566a62ac74328a5a5d617aea67b0e117028d6987b7655862df899417f846fa20b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf924f6136a5bc59777b9471cd81c8c7f1033ff8bbedb69fb0ca3c540f9b99eda3862c94525db9da58e7849a235848cc37695;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3f3ae6ca1ed90cebbec25cdd6b8850b71138d88a088659805b7793071e9793dbebb29bb5708abb5c55b920324b1e7a88641;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haab5cd50c9e55360f5572ec646e01c762743a6f97cca615a68dc4d75b04f0385957764151e2282dd44e63dbd0cc8847c8a7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf68187ff994ac2587676ec157e8c8df84b3417d452e2e237dc0563f70e202f98263cbac3ced9eed1fd3aa0e139318144df2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81facc7ca1ae911747d55f386d6bd12d3e551bc1ce31cab6011754ea0d82983bb6f9cac0e45249bb68d4c70e714076bde8c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4915d2c3403d0be94765ae7a4934790d1fcc29954e092ce94fe4e02c0c98ccd4dfa12d4021da29dcc5d9c701d2570faeafaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd83d81eec935b69503de4a6e126ebb5d3454d431e3230f5ce357835f4e1fe3feea8557f7196763a8a04da205368f453ca707;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa6debf843c634c621edeaf8ace46422db8f0a9377f1ac117fe338f83e6a5f7be20a298a806037c9f6bcd65d9ed47711f366;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6c5728615259d6d83d68e60b399148de4763ba095be62393ce6c014f08a7a3823d367ee405bf9ebcc98045c4fe5e6407ed2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacc7a77360277565dcc06f4d7cc69a7038f505d3cf60dd16b522fffb98d9e915071ecffceb3ab40755981eec5d7640cc56ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7221003ef9fd4fa343a41e3697e64019630cdfe8324308e8bd8b46ed87582efe1f85844dc8c2bb20a5e5b41d897cf82abc5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda4031ef0ac05b4c18fd864ed816652688001634d924c22db63d33b5a0b17b549b721dd09fd5189776e8d8a81f4f4546c526;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h860804890ade4fe159a3ad24f51f1bc3455b8d3defd67f174234d1afd6556851f9b16cb5b9f1d0adac783a3dbbd0c0476fe9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbee45f1cb815675aa7cd6d0c2c7047f248dc41e8cbdd343256b52ef3b8f7d2c0bb934035e8a0492c9308c538f7c2c733bf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6287ed6d096c60599ca39850c0ad049876b5d5620cd473764e3f2bea46c0acbf1ceb9e16a55ac310c905c647820096b9833b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7c0088076bf0511fd2bd3791039d583be5ce69dc4dd113ceeb311ee882d4792f577dde40fc38c748dd0a166bae048680b12;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69e185fedb608fb8ddb75f8b35dab16d72966b2527bb19e139cfa2b4c28dbcdd578970ce5aeaf3c3355a478371978d20d117;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he31792a24a1ad8bd88e6eb0dcf30ac94fcd08968ba6f2234aba2c244bd1c7f2646cc7d5b92a1b8cec22ccf0431b6e149b300;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8543926a68fc5f76041c1dc8b8fe1b8c00385daf5fc9eb92d491fa2e145a522bb0b0669b4b67792e4cb624fcf4d7037d8a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce5a7c4cdf47e195857a77a0a8284e38f953a6fb1217ff508394899d8855075f33f23c714e6bd431a1f8915aeb6cad08a89d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16c6d51c351cb219d7fe7648301b85f9e88fb784ac171ff05c6cf6c47fd0f8a5b36e13b21068fcf1cd397362de29842e532;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfaa8f689d6eaf8cf1e45eee648e21400cd0f040f4116e3fcbf3158d8cdf4e006c2c6383395122c5722c62dc49b00e5475c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7672b00a80a3ddca81b69bbf376d72dd9ff8535fa19ae0472561a25366fdb25a6b48b80563c229a6cd71b57e3fd28dfe2101;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc400165e58947a7ff821b34bb48e100ddb149403e947cc025b8dcf6a9f2199f96939b935954d314da374b91367831abcdfba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7881a1b5f1a7e572fca82718009b4197edf6747830f6b6bbfca48af1e28835f87c6d684df90e3a5ba83f5810a7001e213958;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f0ff9b457036e633fd07b6bb8f504c8bf34be4b8abf67d3152ceee0fc63d47bee20a3eb6dc9d3f289202cc21774e73bbc54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9501f4e7d6bee786f851e265a6fdd2eacba7a3ceeb1ee323618134c9c21f488227b8f2e966d5761e3f17a9b4911c6d91fe5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1224cd5406c3c02230b8c536e63c5f570f4d4761ea88f26f1e8d63d0f86500b41cceb54c12f3626462e213002620dd3a644e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha066017e444634b1108151879e258f4442ff5ed687c748b57a23a9e3f50866824078955510bf2fbc466e0192ff367e2ba2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb0e65695aeec7f02b929da30096b3cd3e2e2328096e84749a29ae5be0d8722f54afe214d157f70a49a57f17de3dfecbe2dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19534655757f5ab79f83de7ca547e4f0495ff3a56fd09f7ffb05b9e5966f1152e304efab3739cca6d657392fbc19c64ec1f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76e4e46eed917f1e39cb031d75d1540629e29d3219e3eacb559d6a1b230b19dee00abe19955df24c14f8b844b419f6ba6a19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6725e8ef751bda5c32bb695d7c4ca2c9e340637f1c045698405d876a87e57e4dfc3ed721c7cc78d0e445b354180f9828701f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e80e7354d354510a3437660159ae15781023cfa6417496a8a382f5be9b2f1d64511747f24d095304d33f6b9d0ad8a6a8b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1ffbd96105ee4387f394da9225dddd0708d75b4d2202da5eb3410740d0e3f246316ce0cb9c255cc0c8597d41722b77bb012;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92c0214a6eeabd6f65098747d3023473de676f99a403e0ed40bed7be497abae287558555606f22dce4bc552a520af66a4b1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd259b7901b5ce09c431a65e68bd58382f0766063242ff29fb16540fec14cf32dcc6cbc01bfc7ed88a6d2bd2ea26c1efb435a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd84e8aa9fc16b8e831883c6532eff520f139eff532b5c9df8aac4cde17205d06eeb7701003b84f0188a696267130fc2be7e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8cf620e706ac1cce2dd8d815efb2227cb770dbe5a14dad1d020d077579ab4d5e7376321070e97564e16e50125750fb89a77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a92359326134df9a3c29efbe391bd3acba2859f28ee7fb0ebcf44850c4da0f0740e3894b5af3d12527136a74d0b3aef2c18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6ee8b89534c61c36b3688e5cbda06e5b304130430034353ebe4401a1090f1187ca03719da48a858c9b1f1c393d17b7cc890;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82d96e80cab7e7094b9152b0759dc371002f58efea598825dfd7824aee8b257855488a8cd9cc56d966f3f5d4573e9fb3d0b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1bdf9defe78943a89f44c7e85c45d5a5d0675e576c120f604aec05128671ae1af3bc3146175d9f394bd405ef2cecd50101f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6937382f7ccfcc298a5e92d7d65cc268d1d7602ca001e092e0b32d8522e498a965a9ab698772d80f537fba899bab8553e568;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6eeac3e4b241ee6cc30163883d325a9475e0f8a9b29784ead2ad439898d37328dae35055e79e5c7c24fc91636aea7d9bbc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18e25ade5ef184a6d26b58f48208247ad6712fbfda927740bbe4c78df59e73706bbe77cb54963108ed2cfd7d4b20fbd27eff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h993d4f1d1bbe2e52ff4249c9d205abae4a9f3a95a5a83db032accf5565d3c4bf58af9989ded63c60b3a1e402553324332c85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30843e29956ff2ac6a1ae9cebabb6d05df768a95ca9c698c0fd2f44a266d837502895cecc6bf05a6343bfc6597fdc6534885;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69d74b02a7f72f067c4970525d163c74bb68a0c36cb10e2ae121c7b3bb7b9a7f941e4fa2380a2cf4b1d68a7a065e4dcf96de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha946e1cc3c2f8d9eb4d4b17833e4bd3d76b9d641540f304a6f30f020a4a253fb65aeb2ad00ee1c0ab75dbc599ee312b7ccc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff1bdd8b971dc82ffee71ac15b8b23219198f186354e120498ca1b1ff3580561207d12057b8099e8c8e1c46cfe73ed74fd83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha441f436ea1489e6ba7abafcdb1d7529397cdd5a99ecfed0bd7ee2f73c97036825ee567597a4ed66df42e60287f3f8290225;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ebb42e2c8bb6b8d14e742e22662fe38641da88990c05071e83ffb150ebf89482c53ad008e8c66f8924cdc81d8cb4c8355c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4868aa5b0d1fbe00a26308a58aa599a054466d3856879aec29c495316b7e517c916b8cb41d10161eaa3acc36647839ccb371;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb05861d9d3a215eb8f10f2e4f4595ac2148e358b2e9c55d1ea6ac100e997838121ffe0e5f11e6ceadee8378f71f789e71b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb42eb984507bc02c4a835a73c39decdc4386ab8b266cc5bc70ab931f124b4dd02f7cb8e4b1c35f3461f859140bcb4d9a7b07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb350103fc1cb8ccd9811e83a4e69f6c196a7000df5699bde173f254ddc9dbe7e97e15ee408986af4f8fc121bd54fa2f6606e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9f435066ab7bd63534b517787cd97be2e98dae3309927caadb38919c2293ae18f68ee40c3fefa8427c93cd5f270dc8aacca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a0624243a4b9b524cf250e978f0b9e31d7890f4da5d63355975638206d33a02a26f865660c986a2dfed3bf51387f82f0df5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab158842db5eaf3d13bb7f856c5dcdd6f4f2b8420a217c8e8a1b32ac027dbebc6cc12226acd9bd62e870fba3d5e055ee30eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4d7f0338a8144b1dd56c67d2e19bdb6ed09cc72a830d82232e6754dcc5ba685b908bf152e1212bc3ae9c9c9ab041595351c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66d31491c0b06f90e4b7895f67fe88f0352e903d76f6d98724dedc72e9beee71c8765323af27d5a91a4e4343e2067288cf99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e26d75e5a1c64120cd3b611abd8a1091962d5471c336db18a536a04c0add8260aa48fc165239297a99e3192beaf886f43d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e88c7a54202c25bde9277472d9dd0acc020b8e3617b29e7037da7a9fbd723c83b028cc75f41c8ec63141a72566a9354464f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98d024ecb32af11258a4c402ed8c53aab84a22563143e3603de801592fb731bf1aaf587aa7b7b40ffcb01004a16396266890;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5f31cceb41024e461941b30a865a705911137fc5f52a0bb72b13b0599b06cf284d8a762cc4946957d1d8a37883e54e7c12d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h498bcced33c78181459afe135ed22c4cdf6477dc01ce8146cf6570d713eaf35e539cfade2d480da874a1c6b33ec9797deac2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb761c42eab6c0950ac956c87fc2d76cd06ea415ee367f16b66adfd627b9aa04d9e556a9537de454c6548672c34110291f405;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51ca909113ada06a2c87a1250f327b7ab39ecd9835037d639b9007eee25adecd6be4cc1b2eb954033c24c1dae2c233d518a4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f88b17cbad3d6e959dd6a27aeea0ee5e259c7b316d85baf596de659e552a44d3e505b4ad4ec6e5de6959678a1027e981371;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58d55ad91b8fc1fe9dee63c4b5d550f457931d413c48142231d256b859fd97403f4fe53c88a09a88f164702125fb00908f4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7508514488c13cbb0a203d7b85903f525602050c219918e8c7eaa18a35d97e80da7b3defbf5b05c90ca4c394ce590d992069;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44620d3a257212a4a3c71d4e5ec0703204cd8c49bac4960d5e7cc7a07529f16265c68d58e44434fbfe5dcbfd62da46c315a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf58b7ce20ce0525d07ba18a5f8f938e4e54c1b9e5d4ca316ac6d042868d98c6b67fbf1ee78a638ca3aa1a31405ecd95eddbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef7dd13352aebb2a589f2fb62a549f14014e711d3e0ba9e117b7468726c247847659e6362495200c79401f0e8f29da63bc0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98b490863d4ee9509a73bce426c68d093c601511d43b9debf1b6a68dce644fb4386603ede0ed7ea8cb7db17bf7cbbf46d0e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b96f96d5db7e457899eb048ca11900db55eb2ad31e620a85f66ad1fbac8ce8da5423d8f04deea9363d04ac769c40df32891;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28541d7af559db4ecf547276c3e7e5cc4eb1fc288b8e79aeb57b5b85b7967b38464818801cb9a89eeb683172620fd2615dba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b3e76e5f125d3621e32f87ce0d699e24a5a36d49c59399750d76ac7d25d337ee4469299fc2fbb0d8be1a6de0409b01e5f58;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e28cb55ed914745c556648d3598f0419261286f4f4ebcd0e0f8e8a609282a4a0871b0b1c48950552d25d2af228fbdf5adf9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbed33c4b6e453f7951379407daa188ee822562949e62f678b5c1098cb7b70c7cfb4f21679fd2de82ca9fa59f1e73909b18d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c67ed559c109e56efec6c39edd12ab3009e034a7f7eb2fc4e2144eb32b1f98ebf23d02da6537b68b174c1acd0c5aaf2bdfc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7915039ed76a0c91a110f39d40ba7f25a29fdf8ff71d22fedcbc2ac357773bb620e1171c2545d9226744ea222ff3b75c7c2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h195e4b490af9949e199b19d81b8ebb0149655817d099cb1c00779e07256d9294df5f0494f95c13d11e3b05f4895f2398ea3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd98cab52bb77941c41bb5448b97dd76e2d548578711b7dbecd6caa3c5e62bde14dc72a3d077ce22cbbe48484e45f0381e3c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb52b3fbe926a0b6be18a37109a7c44a1324ae9fbd7b52024f0ee88be2eb41bc5940bad8dd444088f9330c364c46d4de34a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1e0094de302cefb3447aa33db9f38e8bf4b108802ba5040ff58176167f9e58a4c8315b76b50acd7257eb62bec017b3b86c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fc76bebea80a2f12441ba6aa9b9e280a573447bbf38e60d231d1a3776642576d92454670cf318d7b7d443cfb999d152c089;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc941884bc0888d6d7bd7c13edc1d37b5fe664350ad6271eb70039121ccc6dad50f781e8a6a1044ce19ad1ae3682332a373c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47b04a1a9702ce33a2301034a6ce59a53b1ef1863cb328c4367133be42245726c86fe3ef61aee352fd5f24790a4911aea3db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbe13aff0f8fe9c56ada1be8705a0fa5f9d42038fa3696626ac71738eef4efe2e698dbf93dd87c635f161cfd116fcb1b41d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb89c2a11131e759cdea9105fd56fbe24b058d7f9a058832eb125306fd5559daee1bdd769495ad7b197e97b84d466448902b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a6e0394aaba0c7af73a9beda52503525cd8d9df2e2ec3815d8cbc9608b93d9ec0c7ecb299e76256452422d78cbf06dfa35d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3270d15bff36d8c7132d2bdbfeb148c7adc5a9415bcc3c38a56605778575d3f7fe76ebe9173181bffeae0fcef03b7f06667f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a646970dfbcca0e43a31f2e01d1f68df08688768940d280261acd476fe4981bd1fe127f0eacbb3efdf43cd7ac72cc602496;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h354d632c9253580816163cde97bffb21bae2efd7b436a8d1b6770d706f2e57efd3b95388928ad6602d7e3d590fad562ec758;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h398a058bb91d8344e00006b585913695d08438affa3d77fa3f9ebe67e1b5f027d121a0cf15516a3fe4394b9ad35e0e2635c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7af0eed0d9d11632ae49e26bc5756b7529590751c739af6b316c4b2d0d74f45a6c2d6c63a87798be741a8006549f92f29ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41849ccfc8a6e0407ce3f7a4c0ccb89798c3ac9c263786a167c96d1d639516146dab904a83014357389099fd6ca3812bda85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6176c777866f2f247addd150b5027d33fd5ffe56475a88626511e6de74374eb11ee1e35e05cad09ffee212d86e773e5d82ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c6bd539c0e7dc1bf68a2ff9f0cfc2fabc5933142253a6e42748dffccb295cbb3280e12020e56cb248eb4ff33dc1a6e1b91e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8244d82df645b6b2fdde895ede0957e9f1e4bb964e0c68b0a1671c833cb34801f5a7f60c3cea29bad29afca227a5ff47fc83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f0f7f498c521064a6da17a44f9a7c9dbd52eb05508e3d3f68db85caa65f4bdfd324fe22ee4122fcfc20b9edc379cf41ecb3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9e62231a5b64af322b896811880bf308135010b8a9d2e00614d5ae4683c1297e2e33b1ce4be59efd98a658a9063adbb3a18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h699fcfbed382fe3a30b5b1719ee923c1a9ef0ea48db4ed3790b7928fce72ad322966056fd7256e8a88ea525ee6b2c028c511;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6307670353d32d53f13f40d35e78df136fa63f517fb49470d8462be3f677953df698ccfca6a70ceb5e41023ef8be6240ff2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h841b232f3d963bd136841e73f0e9aeff6fb7a5c6e54ec49b1e0fd222e01c9e22172f702911126b663ddf7d855d01e663d042;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haacb1f35d8b797994e48505cee7829b8001d679d7658f99212bf79ef80fa261a1fabb782562e051c1593fafcbd1a119d96ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e72958ab610b451237f1a507ea6fffc265834e8f41d88279202a835fd6a08a5256284fe42d4370693664fdd4407afac44e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf71f63a95d35606aa284a2c372de2f2495766bb161c87a91dc3f47cdfa6505b39322c4e1c93b675793ad90e4c7e6329a8c17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8b4b92fb8e802f1cb27e01b9a3395aefc2e0419db1c18b638adbaa02480803bfe556cf4aa672a6a43ddd5c74ad0017af1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha35267390d7f7ecd41512c73b6165bf87617ac61ff9ca7a4254f88d0ff82c557912997b94e499536904446976659d6329247;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d0ced329461478fcf2149dee98a7ac1fbcb8b279f298535a26751435829fb5d90176edbff4ef9f4f0c207925f1a4ad33fb1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h814cf37a39e14edee2bac6b8a4e0915b01d3a90ac6d70398e8feee0ffed55c74b14ff4e1790f557024287df23aedc74d7f69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53fc53c362ab20a77eeb8599fcf320bfa894fdce93d01873f9906b41d4983d46998b419c27c7f9e288a82d6a2dcaded2ec47;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e99ecc0b2de13d007b793c239764b681156dd1e82bfe0bf1c903cf8fc638b437086a1dabca41ff247d271e53ddc41f11410;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he64f3605a8cdaff7a8ebae668c981b7902d9e7bc85fba995cf6172c0922acc7cf0cc9ebf3dfe5ae5ebaee18e394d4f1eff92;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5450f6828174eb3fdf8eab45bde1de814e35c88488ebab09d517d68731f8d5070a692aad864054c8dcd4fb55626c65cbeed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf188c5c600600fde682d890e30daf7e4507fc5ab96d468e5f3f8f0c0f9362eb19efb64a661207a6a749036bfc29765aec933;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h674383613cb055cfe49117571712d9ff8f484d2e1e6905a7c5f7d144bbe7ebfad1d7b7e0b728a41d7a78e88bcd7c55d42075;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9a82f7712cc2d8f1e1682518c07f7723fbcfe85f8ffdb003f3e87c0a436194c199aa9ecd4afec277410114c891531361a96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dccc217e802c00af32b033fe1e7df627cd9b237154d91f085f23511b647e2e586cabe66ffdb3b414d773a6da55d0291ceb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca9d667942f68bbe06bf535fc8873e1bae845a6f07b1d60d79b120eb80df14fa4d4b1829ed63da97e88afd229acf85d47d66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12050ebed7bc6ed752a1b515708fef00063797c96f0a81a6816f9272a528e2a2246c68a7b637a32d7298c43b637c1ab1d19e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86ab3f449ef872f383bd44e8cc091a414a3e165578369f26b5d9be3ed5bcc7c0653bc6ac9b1feb49f5a038922474bfbf3956;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4475fa305778e55d123daee71ce9868e3561a87f35384837cd7f2505dd727f3db6c3a5ae106e87e72b45422345f575d9792d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec37d593c51e5d01947727e13b9af0159a862671662cf93c887e70de297e699f868b56c1c492a8f38413083ca12848ff840b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h893be5a82413673ea05e3026a29eba3012c585631bacb4d302ec9b1ab1b1be05d59e2312bc2b3e8da1fa1cddee77c9d443af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2d27943093f84b9eee34b61854b6d6e96962120f8cc0631ecb818361ee6753ec02dc1502f1c9f3cd45c8b7bca00c9500550;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbec23d1f776a6667c8177d0605a98981f7e5c7fbb1ed3c47a487721bf5e652c5bfa3dc264d40ab832fbc4101fa8ce4792790;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h771ab1d718c38c5b9c4c9c5461fa47257b518768138b33807128e8faaba92321954d8d3a38c094b2cd8cf567af64b68fe505;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h719fcbdcab805ee97ad5b56df4a4701dd9a80c90c71f0ada8069c42116c60d62638bea2b61b1348ea7db8f23cdb7e3cfd37c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52cd288ed8fb42836ddca1df023fd7cfd4c09e61467dcd5779efa914f30901b7ac559dc53a4c3922375dd97382c130778ff2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7877fde35c6851abb9af734d36b8bf6e6abc2689f951e801bd0394cf8070e31787c404a73419e78d8b0a945227743972fde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2949dbc782642157210814da7fe6b783bc919a48f23779175395de6e64b1fa580caad5a4a0cccc4c5711e1c409aca82f4a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha847f742c086545bee9092aa5c39579a0f6c7ff7a623d09c014e53d63c6800fa81b4253757a1c74b5cea6ef4683b24dff7f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a84a108b2f8d55c2bb29b3eb72ec7885dba7ea0caeacd9cdaab9d49f27c0bc1f9d500e62e40f78b3fd338c66eafc513b2c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h224f7d8fe87555ee06cb1f5446587464019ef1a1270b35af7498ed2c5536e99f9b261413d10686952948398bbdc9a82c0467;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51e1051b6b01f9d605609c2344137a5b36f902d1bce7ac28a1576d357c52f7ceef17659383b734c028d96903b073769ebf31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h314ab1d2a50b1739594b56e04ded35392d2df040b399dde3b910134c4ad6008d8f2a7418b3651c67bb68f1e4869499f29127;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2db2da43554aa1e6a613792aa49a693c0dd493df85766d3fcbae089aebb1ba77251831545e2dfe17aae48d6c237c4244472;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60fc1f62756680fa1aaa5c0ab774545e4958848092c00775ac4316381c2ac98d300ba752addb7ffc4c5e1768f5f895bb3043;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5cd3dca926989cb1ad874383e8b8d12b39a00c2594c0d7facb0bc02f27516b710356ca95537919ba8a2ac12ae2bfa85512b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15d36abadafca8bfb03328a4ecbe9e80c4f105e52d367895b71c009d025de9275e15a37eb5c3e416aa25ec459420ce6f1b69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54e277649e5411391f81031c7e99460fe99269ede98cb5938a19a3bcb2d4924c3e7e10ca364414fc9e20e10c9b31ff20b24e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0a25d2fee5e7dbcecbe3cf278c8a2393c51a8e4f4defcadd61f8f8c1eb970def743f1b177d7568d7994bd89c0c9aeddd013;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f401030f40fae7ab2b51ac20834325e61168e2006e92a58fa467a7ea55e706233652c97a5da9f3c10bbaafc86b3305d47ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80fe4a42231217f5ab7eb99b7be39500cc885aa049085b611cce7b67049f785cc7f62897b929956b23190d0dd7b4ffa4368;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48a5ac7411f2071cba76867d8eced02948d66a9ad6510d9c7e1444b564a70eb1aa7570d85d7763501616821d8f13086dc07a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a7b50deda3f99ab5cd7b04b8459fb76788484010bec3c92ad23ef3fdeb05ce5a04c02bbf788a015c6ea06fbef0684898e72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd24f9eaaf8a036052f1f4ab6500d0cb9eaece15b91d9248b3489cea9bfaed09529406803fd95b5e94d3eac581d163ac6c277;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1cff245b2093c9b813ef95591c220735abdd66226c5d1d017cbfe1331d1eb7e22c92f67410039a16241cfeff8b84d2b5408;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9481490a986059e0051dfbf80735eeb92ad3bce1b11ca1012667400419d8b519dac324767b16b3ae2a28bd0de808a89329e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa246dc27055b51af04cfe47f281645f742333c0b75a5453d2e4cc64739ebdd07b5e88cd81c9a8b0b54a3e508ed7db2675d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12dca0e073e7fe04e751e227eeda00f591bd48d0898e18a2ad0acbec7e198aa2de2046c34b62a56623d10952403eeef83b06;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7885c49eb279f44ddbd14e63760eb406670bccbc7a28fd547fe260d3669a638b0a77b1c570d49491405b32d11176f73e0080;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46232e6beb6c049eceb2b5609949a1130c4ab241a3ec5ac6538581a9e381e342741e8a6194a508ebd2a022b08afb596eaa7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b568562045024551de305bf9a7dc27e2225d556a9cccd587872b0490895d0b608047c9ee3b6f40fd23a89f480d2fd9b1127;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6e087023323b5c3bb2844f3750585b9371d70402c3ee9bb038e7b6b688316d3e1e741c7fcf16e07fe98b652ac2b3719be41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h815e883c16cd0f984165cd880c682062b65f350b40abff72ca1551a462724c5b724d9cfa8f9de2b61f3cc2a915e194c50f8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8212f5b929359cfa18417a3b5876daeae54df65ca826051b6f56c46c4bf7098f5fb0a63909677cfd230724b99736bdbac55c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12a824dec96153441a56bed40ef09482f6d68ee8dc5137fbfbd4766d770e24697451e698511dd3708b4376b83830c6cad05f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7cec8377ff8716bac66b7265f23b3eb400067a5f0bcc70da799be0d38650ef3c7426e40c72d914c2ab07979b77f77771e20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h708013d822d23c51beb5e7ce347e464a0da06a61ceb7260c987b5c893f553fc839c279ac593596f7a992004f303c5339f04b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6976ed5c5694a4c82b4f04444844db34cbe377d713e859e2165e96d00ae9101a6cdc894d7ea3cae75433ade3bfb9c5ca75c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1cfbe1cf25f03d036f68b55d6ff48417e934a7e46791965e4efb0d98c6c98fbaa613012d6767a5d20c878efa436eb225ef5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a0c760bedf0c14e1488d2f0b59102fbbb6b9357f88a12869fb7284f25a94d601e954cff84d22738d4aab5fbe540c8a4e225;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3aad0d8a624208bfa5b01dd94619e499d90701af1a12e3d447c05fa36c50d201a64e0da87ad5d0a8cdc2039501a5a6d05d7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa0a4c84e08ebc0132fadcd41613da96be42d13d72b19596752eeafaf9be37c8f33d72bf3655f4130b1f5a85dafb024e317d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5c00d3bb50df81d2ef23a410a08988f4a098e891fa33d6bbff9656c97ecd4dbd8aaf782d20567d658d86fd4f7ca5f8f2f30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h756f9c8bb1521ee0077b50612517fcb8c22c332ee7dd79681686a5c114cb7cbe8c698051fe06efd5f1224db445c57b3a276f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2b29ba8cb2af0e5b19e16bc3245fee2600fefffdee79517bdab65d3c1a62ba0e4727c506d4ef9fe406cbc6f25e483f4ecc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbea4efef5516d6f9ecb4dc81de0f9ed9304b03f45ff3a8029e2af9e97bbb098cf21924da78078185402f10d00c2d0855b640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha36cb8f406817b169edf11758467a1f1db4400f41c3e7ecd1acb0e5a9197a237222ec1f7da10298b8a7cb5ff650950ae9b15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h760aaed0aca09f5990d002112303ac1c67cb8737b3bc024a3a8164bfc63914d309bce7e5e4fc7c6bdc36e6387bf5b696bb96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f691d1874104b7c0019ae8b9c8c186e50d92702824a8718fe35be540b50744291822242033e5128199bace4ba61351bbf67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb37594ff76966ca1f456cb6512469be68ebe2e92a54e5db8e25e0451baddc42945722eb6899646c2aa1eb0fa05f31de0dd67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddcfd1891785bb223cfc3636c3e957cfde9252894337972f36e5a0fa6a777d56719a5bdc6d312afbea3d859d5848646ce582;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3554d22b09405b0cb2419348bc890fbfb6ad2831dc5bc9f65ac1790f21208148cefe3e0c568ae31968c1d195fbce5833f1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he99b1b77b79e0add22e260f5d3e635b1eb88ad4882d7591fe3409b3f81858f2f715eff20278831b886747c1211155fea9cde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7eb21aff41c9029b9b7824e7cf3e89a308133befe790ece05cbcb0d54fb8902218f7644bbbd594809afe199acbcdc112cb19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb915571664c8235a7c5499aee9d901bdd16b4d9a37a915961e0c9c73c443eb55c6c299aeaa303a47b6e431108bc1d641d94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52b59bcc0a8652c8259d507888a646aa0df29cea1421dfd604e10916194904a18a8b5968e13aade7d55d32e0b460c23adb84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a3161cef0053738f4536e5892afd2fb40b45a20b28721fe806419d3461935fcb287865b828d5324e72b80ca527d29bb9375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce5a72ad8ea811fcdc7142412371a7b5de25e89cb64b44d751f8fd7109b4fe48154ad2345b0d9a5e6dd6e29e45432646858;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda622e4c140ab49ec794ef330c1c479a9894829253a2e3f0fdda54203b37e242f1802d2c63102024278f603dee2b96cd7f50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3d3bac4470afee49f57fef84d71fa3ced7dc0e2c8c500ab8b247e3731d44fc6390f27bf09c1965ef492d0ed75ba1847dc99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c3f51b532b577a0bdfcc141da57b4e648cebfca934b9b04711213fa39f36e768b1adb732c8c8a118730aa2ab803f844fc5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h411765f898b2a7f4ef0dcd103fc73257a608969e2e80c534935cfd9805b25ce850f9988f11daa34dfae7477cd82689a122c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a7ddc2ec84c2877353649621b8acf47993996d368141cb38f996a8f39133a5d6db98a15545e5dc7e49666036c3504941eb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b6b8ea3ec0e95b10dc03ae5f6c3ebabdfee34d342f4ee7d4c1161a1e1292506595c1c0d6818d0f1962226979424345733e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67f6b271fd69c4b34164a6e8051e776997e7207be9536e80d7fb02e018b676a63aa50d3d60e8d31c8e65196a3134e923ee51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85e501f7d31b1eb8f0168c07de603e308646cb3faf379c9bc3856898c5ca97d39e4fe962915fb6e9c17f8b19306c5e9345f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15e17fd6729e74cab61eb0b635cd9cd5eb537960ad7a02b4e721366dff83832806a375dd78090f60c766005df9f92963f647;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h805f5f4f0bbf0d27fe8f5e38d248013f280dad54819c47b82e24aaab28d2ff47a4a9ed6969c24a09be23be7a083be980d78a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e849f707e11c3327c7c1faf4595ffdc4908a00cd1941ea47cab706128fd0ce2fefc14b38d2d5f75be79634de9da46f45d0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd926f51b0a42b90b3b038edd1a9f48b23efefef51b003cd9519cdef8d70686261e04020868fec9c1f86efa362e25739c2cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cfae8cb936983de62ef955d397f5a161d00c503230333221168e1f0142baa3f334212d19b9833a04d8cc48e53c6e01abe23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1958b39627798ec40bd34437f94195b9456c782eb02f1310e8da10c8dbc6edecb56e1854f21208855a0e22cf9a95db632415;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98f117163a9df1525c59dd06e1bc49fb93836652519a48ec58d725d0fcd512e504ed81e8a8377a6e2c7bbc95ed2689d52f70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeda775fae3e94968f1d309f683c535827d3963358fc038ffa4cfabe91b5ea33675757236ba291ba587a415f624a5587bda0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cb1b0d625ab5db0735dc804be6ec324710e47254b19da937ea804aca690ea3e88c60c158a10f31836573bf2508302c07c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h193a75ff16c1d6486689c6e518d9e7137d8eb2a828b3d8e0f525698b88e6919302ba7350a9c449fb31222eead40ff51d81a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a66133094ff95cf0a3af8e53c8b27a6cbac0ad1df9fdc909df46a30888eb6ce1f0ca015c9094cf63a562ec3e36fcc1ee469;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4843a34e0a928d0e9a166725174fad49c14e234ff4e00c24dcdc384e7b707f019f1d3faadf6602a6c429a55a4a740bffdea5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43435bc7c46589909ae852c82baa95686d3aec9e54e2ef186ee21f81e0f98e19822e1521673c0c0cd40b7bedeaa927a03d53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc105169117ade51f03d1fa66fd0f0ff5e85190dba19c83beb7d359dc59675ab4a607bc7f66ee367993cd6f9d5442bf5ae84e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2392bc12545e1ae9d97cb4f1b266ababe46e41423ad8b1d6111ecca854d6014c08e6dbc53423033d0a2bd5cc9fb50a567861;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7ae5eabb0ce477e0734ff5ce9444a5bc7a291f3381c0064134c83b164bce45750056163912a345e489510df83e034364715;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7e3cc74a706d9bec70c3d37d42ba6690357441593f622dccfa0f68accdf8e53a2eeb546d4a4b27d75a2346cc09b7e0c3d8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he243f9fb64a7f32393976ea2a418beb1baf2b7dd7e4bb1a4f8a12ee3947a5a99fe91de1d15d5f6dec856cdb518eb1dbeb367;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28b4c7a035871d79288b39c3ebe2185d272fc8cd550b2a217f3b9f97044f6bcf776819b7f25875f34283a3397d61762b33ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf535ad44f1ced2495895f9b6c6f93b9505d6887e5cb1802601e6bd64a5f6bdb3cf29e1a48501bbc216d02411c85c1b6b5c99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd09b321cf0f159cb1d025d3c252f9613b4ec123ed6192e01fe315132adf95d4bbf9b1fccb0e07ab8c35c98acd8c141d63d7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffe2080a8c97a6bbc980ca634a30627e3604724642a47c6342a4dca842d6d0bf290b9f893a1fb7c31931898ebd06f414cce2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ce9b701bbfbb9a968bcece76eebbbe38b6c6baf9601b8d299eb62bc7673fd090bf5a8290242d4f8dab2612e15754b2c9a64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h284fb4742d8a6e12629b180db0cb6b647bc1c2589c2cdde01dc833c9020203f1888a3003fe143acea207b62e671c44643b97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6aad64a6682fe3d0911b571c04b37c61cd3072fa47134087c9dc75d7d780cb2f82e4355ef3778143667bced9ba3dd5bf8d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cfa7687b9731fe2324d5e1b2d10d23e9530ce1509139d43e62c82f7fc92618a9480b3fb32572608bed13c3ea383ac197016;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf84bffe332c74c768223ffa0774d63783d680c879020a9094122f157f9c941f6175ae72cba175853ab7b4cbae0549550f3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3711da7a25e5e38b171e6b8875b21e6e44c4de2608ce4224117bed051b8d3238e67187a5e20bd91e903603368f5fbba6448d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haaaa58c43aec48dd1af57f363adbe6d23e89681d9ce8f0ae4e8f5869847ddb39bb263b768c838905be51e535f6696e6f3eb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89040bb1d4aeddf221e0ad152e8c12f1219e06d10a53c29f3f265faf0b3524c04784fa927bfa82f14e21ca74f6f8809e3a73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bfdb9e1a4ec91adc63ff3a822e2bdadcdb51e0346491daf8e3bc6f985d17da7547c8eb20d1fae29af2f89e12882c48220f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h792261658caa31be358c4ac86fdb514c9428376d983e7b518fee68aafe7c15e0ca0a45483dbeceda43c871e0618a6c27e2a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he51ded201ea5634fc53ea4286e5ce7146223bb9341c5531855651e0658816bcf1cdc96e0364f34133d33567cda29f7d0677f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6579090f4e554a618752d53e44c30ce30b33b72c6eaa8f1cf7e88f45fe882d043be9f36db8fd3cf0106aa95e3f8b76e4c936;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5efca644787da3184a13aa32f0c4ec5300dd878c88ec1b4436b0e3529f10f69e961d081433b9014d8a6b89e470b1b70aa60c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58b05ec183cdb53cb4501d40b92068e398ef8375043324f17fbdab9aeeeeccb557d835556803021c219fc1519559151137a4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcb7154c0abf15bbfa4a3d7878adfffffcbbfa997fe81b0b4f8a2c0b03f3ebb45fb165c8d066d705a151c9e48c78a9ab4d2a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h681bcc835ef18c7ec536322119f82c92ff5684b3d5f23caeff0bdfc72711075ddc3a72a6b05006b0091724158b3b089c059d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he895e76623e340e47ccd1290862520855f5953175b3e877f00014d831414635ed5f6331470651c0ed065ffaacbf324b46fd7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fd0cf1cf9be17dfebe561701d5a6933ccf1ef7bb6224bf1ecc4816463cec20ef866b5281a30d36bb6ddc7e1442f1ae9eb2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfc583ba26e99162d8ba2dbef20f2b924e3eaef80252588f71477352e93e0de58fa24cd886a4580b98a4f218dc05e237d389;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb36ee4e44518001e34947394ca618ed2492a723dd95edcd2af2eac65e581c7d2ddb5d2bed49f1ed6045193da9aa7b38ec51d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cafc6bddc23c051e7a36064916e8fbbad9d4b8a09b59ab7073693f8322c109cb5ce58f6a532a1aa3380200dfc292eab3211;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdd866a0c32794e02228f15b0de7b19974a59b976683edca671105b5e9d6063a00f365988c89729dd2f91ef305ee5dcac002;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b41b36f52be4c3f2427c9155d414e4ec6e1ed2d38f98338b54facc2838be95c131b5613f6b16a19f12e79435119f6868b29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf00ebabb0b9bd1e515b82e2cdc55eda17742c89f986d3251ba035cdbb73b7f6dd7cc753664c48df17717c7d324c682b43307;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24f1b106f2b4cc1706a274f70d2539f4a5f6c7b0bc2896939140724e70632009eda6cc39ada9c4375f20b3b190bdf117dad5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93890f56d8f4fecb0ba8572cebdfd74bfd7666a46c72a1eba86a2e369888707df45910315e6b70098f7793cd61a3d6d96972;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86af59ec82406b0ff476cb8015b00b229950ef4a43e0291a96218f4c533cd7755b02c9b8c04108a04961dbccd54d9170922a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h332b10291c3d6977180eb513d90362c381e55c077b8d318d01a41e375289f28e757a7b6c2c0cb6822d082a7a30e1359db9e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ee2c2fa7220e248d57b98384f10b5669a990c8c8442ccf853d882ff5b779db5147b6d85b7f14e1c1813833045c9f424dd3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h834ad1b41cc84d1105c042966450aa4431b1a2ae222d44fb378ae2dc0e13c0e3fc1b8fcf1519e13849efbb7e13f34171d034;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfebee381015d60b3fa986e658e2228f2562e6769aba2adec478052fc2f8211e146b91b1e5db27dcbfb75f8c4d041360c8aad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60e6fcb4dc2eec7e67c567b374ff17bd583fb8580dd0045516ee8898b2953b6a6b4dcd67042800cb47d364593351e967596b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee083fc6fcdc0f0ab79099809ced3103ca00233a793b99aaf5bd4f2e04214f3efa790bb2e5411858e25d6682503d10228d51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h640bfb180c62dc317b73e9e4bf68c6eb56d4b3aa25c92c0b256b67a5c13f03e3b364c10839d011bb99d5eb59a7fd158d0dbc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc126f71106537617eb3fa98bb2c0e4f7fc866250b4410573fc5f8f94cc9f4932d8d1fbe80de88712c5c04d06e99a192bb8dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cccc1197376b9dded33cf665d4c1ff714647f3e7f292f5608e71774c78c4841d70541784a0c40fa1023f633f688903e2e1d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f15c1a5e08409c851b6d2014fcc59fc842ef7e29716134156ff07b309d5170b00b0148ae475c5325f9984282e429373a71d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha791e6f89d7a46d3af13c68d2a3b2f0c4853aa59110bf25e23e3de00adab293c89123accf03cb7adaa00a43f20ec11acca65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9728b17a70f258db1aafb5b807d5834ad19b2cdf09b8a1228a3cbecf4e9be086f67f030d0dc1d280853ea7cf4dc9ee4c28ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc16b4c91a66e3cb68de2bad207b773363d0317ea5f6f0cfaa23511b86a90169a60cc95c0d462c92b4dd2a90103e4ea0bc765;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6920d6667d383635ea8e750ad2b2a8a02dbaaa198ccda38c7bc9ddf0c1ac46b2a93a82c004e56035cc066126a0c0a61125b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc82fa7cf7bb8d049f368911c56d21d6aaf1eaf4ca48efff014d0396b3eb195305d22bf35ca72d3a8bf0943f47c64e3969344;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6035c6f7396487d55d2e079bc9752e640a55191aa4aa0224b328a32b9631460207c32408570fe00eb396ba59cccb897ace6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha21aba56cb51f51b9c2b8f16341a3a7b57b5d78f7b2e4fba5c8c3ffa59611fbe1c423a70887ee6551e93c6f1bff19182462b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccff84c4e1385c9f559eec7bb133d8ac9f314e85a3a1826c99674a85eab6084f0b9f6de66b979034400c9e505674bce213ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6efe11830a04474098bbf49997e8aafac253702dd05f994007b38c7d32d8c42966d4f90dbf9e6760757694ee502523c8c090;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84f4ccc1054b8b4195488f6fc83f96f9b081cc18bdf82ed270c7218f15fb6e4872a579dbe51b03bc518737a3509fdb8d33d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53fcad2fb4ec6dfcd592c88a881a4ea54cec216eb6b8db5d80a96372350e892215ece2597231f282cc198e386db9e6db49a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70e90017bc8c6926394526d82224cae62a651ede59aa158a7de994bf30747bdff9c0fd6d02ec44fa44f83d0410346309254d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6a643983c2e640b7a473bc50b190a8e20886243c9651bec2aa070815a55b4606e7dfac102444f7b308199f15cde56889c75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb362c4603966a65ce36fc6a0e0b3abf67f9caec0568fbe70385cb00767e2b70d67da7f3f9bbbe55fb994f79e6297bcc071b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9959b41fcbe74338a1b617e62819cca6f56680fabfb8ac0c7ece92d24d5811d9c801bf1c98882d003f6d76448f1b85d8a954;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ded0bcde3e56f453723361b5ff896673924088b1ef1032ba614ac9a98e07ccdec5380b0bf34a026a42232e077917d7f5b66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he47b8ea55a65aad045f65bed87c7d9623808d14f4f3db64cbe6c12d5070773207c87d64d21ed807a22b1cf26ed15b35ef860;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a6f1c4e94d524f8383158b2e56a8bd0a7cc67065f6f63f3386a6808bc6cec323d22d01e90f1c00ce43e034fee92166d4e2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee1efc265cb529762da1b81db6a793cf82eeabdc5e5ed635cf51c5f1fa4d4ea4a5dfd3bb7dd7bedbed6480d5e325f5659e96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c4654ec4fde3830989da39b24415fc2323a8735332c7b7f8481504e93edca12530c05fe29aae75b99df948bf380abf68a53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f4dee929081ed5e638bf9101908e7253bfce8455d1da9b1b4ddf63b0aa1c67b24e9e2949664a9c00bfaa68a2a60c07d6d67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aaa9ea93fbea71580873f18e5de5b9718234492bdd0773358e23b0c2195838419eb48efb065cd241ffbc2f0ad33ef55f0c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h858fd5ade8ca65c25f32b0f31187269cde4c98d816f4b5079fe8c606f5d99c550116418c0bd4a2ec3f1950e436b8a8b7ce89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46c4859f0829fe43948379246e04369ade3140712ca37ca152d3ccf75f81e6289719954cfbafbd59c88fe592e0bd8825a1f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37c28a6715c8b1df1b14b764ab47146eafab264d3d4b3d20be6da71f4bcfc660c6373f42f1c79d163e5b0256a5f9e659e446;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5da52b0794d2a43b2e17d29437c41d6694562154c1273ab0b87864631940a6d6669e6af2f734182c1e122e3b6a77d8192919;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3a8b1b1d364dc03a9ec2abb6e722231070844db490d457a0fbd5db59375379412d6e90b985360320c6bd2c08ed8204c3998;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b087ee455ce02eba46a3f529592e29055bcc632c4ee7d8c534e01880c84ce54f49d3d0bd82fd77d9dd0065e50fec836c8f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aeac685ffac107f47d6a57d665fe16447292f83345d5adce067459e77bad04859a9cd00bf3b61844a8eb80c783565ab7a06;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfba3e6e90709c16a665131c86f91d8d5cbe2d3880b6ec0e220fba0d436cde2813b5a2ab7e08bf23ff956463ce49c7aad8dde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3142fb9af1cceb6a1b3cd7de062458279ead9ae948fd7cfee6757f96e59a31724ed33cc535ae7d80441b57e6c3b9c36991e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he11229222e097a89f81baea1c1ab7bb17a643b6860fc605c21e8d72e268670e2ba81d8cc0dcbf6e3782e55b980ec9b3841dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h289870d1ee418df9dc3652315faeef0b78ee84686e4bdb2664e52d6f0e08b7a58dc8cbe991a6739d9143bf5222f2f2ddb302;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5734f5e5e899f7474bab03d43ea5953607c751247388e4b3f7e1d3f3cd513b521f5d0544453af6572df12fb4ae809a1cedf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f57ae31340fad1c1a20c3a7fe1ff1a4b58c965f3507f8e6a2d79f4509fe2168f2ef91f5f111242882fa74a2cbb6d76f45ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc08fd348038a6f1ce15dd6112246ede4c87d100a3ba9a03eeaf57791417d63713e8a919e21d25938d0eca9025f85c91d1ab6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd40a2681dfa995fa9dfe58742959a53dd760159c174bc401ad1923b55c362eec37f673a280448c1d0f14e484b7b464d4d214;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4a0c44305a158692e4ce331ea6ccf12a7e6625ca143d8dd2955b7d091f7ef5ef964f872aa0dfcfbdd78a2e00b1caf5ed8ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e2a4150bfc61f076b08a3377da532f177fe7f5e06f17df13571814d1b1f2de623b3508e16a05d3df7dac6df7de85ac9f1ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88a16c62c19b5d360b985e80e38aacfe5a115979c739c648b257ddef33fe9a40d5f619b87d0ae678f75d3eefe89bd13a62d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7777dad02eac6346065461029c9b69afb2e0c6c0ce2194f70337751ac4b6adf0958df9df463dd52072347b6d6204673e7945;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf27323661312b9bddc40b86011a4ea782ee81617ba49101c6eeec54422ef351479b396d19b81614fa6c2c62a6c20f28feae4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94054d4ee92483450154735dc2eeddd3f30228f3c8de4e7896d56625c7f2d919d2eda4502f9490282d34c047e43895962ed2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76391bd8d3928f588c172198632d1324263bf858bd9d3c5cc0bb8e5f81c6672f65b8a3ff2a226dbb6ebc1f086e32e1a1c577;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb8ccea10d462125e3ebc51ce2c00308f982a9d1590b9fb9feebf5211a7b881598515f82d9cc88c707e26a70844ab2eade66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c5b087c412cc8f153164964f67263222ab4f7101b10b961b12bfe5e49a94a0d40e7011490b39f60b54a0dfac47735f77161;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fa8f1c9b682c8662ca1aba904036f2a4268297219a386bcedec0b4346ae8149b2931ea49beb7713838a79d0c17459778e55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf76b2000e8393dca762fdb27d389d16cdf9ad346933927b0f28b9d08de896f282c5325639156401793b0160866b96ef6a89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf03c67feb5aaf6316a6f9991501165a759dac1d1a1b1bbc03fb62444be85737310e06e487ed640acd6052c386b8228031de9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h562147c5723f3e0b2ed4fcc85d948935d5f04c54f1288b906efd378224173f4894345708930b29ec3ddca3fe719d29d837ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha45d65d6103bd0ba8db6e3344624c8fc766f620f1df8f68c341b1743795484a22ca59674873e2d86e8df31215f21a872b77a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a78c9aaa12a14bb2c3765b9f986506a4187318e7f8f0277291b52fc973e3ed12b8c043805eca3db50f520223cf03fb0e0d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5c740401c1f51a5492e2a2e4d159f30030e3d9eb3af626fcae52317ebf9a26ec7409bbb291afc09fe399838c3b2460d69c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ada8c923f136bd77f1d28f46963bd2164c7b7bfb5e2899884fdc36cbb1071e5f2e5039beb99beab7f342ab6ff9a97037c1c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a25ceba8b978f7dd85c68dea845ad41746b8334a973153a365dd29e5d52d8ce63e2f42d82914281d32c3e9f08e2303bdaef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0d59c07bc50fd4be98f30355107119d2d3078c2262cc7684f7dfeb91e609d63f332f9a190e417fc164c54c3505e855e2c3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72006973913df481a3ec69a80dda5148d95440cc9433e5a14d219758719bfaea77caa7d71c917e0cb92d15cf5608a59ffaf8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95524f663099d0f120299cec1aae2b7a6c121e2ff16169354f15f9cb00fd922706c118cd021cf50ebf138b3b0d8a8c92f3fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a06b482e23bc689f99bf31d4aec53ba717ea98bfc0403065d6170157c405d911628667d6f4fd20e883c12413a2b40eca3fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38afcbba226650e902355af63b9ea499cdd6aef2e7318de014b370c7c58b1ce60647087e0f2b27980bcc27bba02ba2190f15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b066eea749df79a2d0aab66cc740256e04da8df91a5d7ad287bb91838e2dae8bb9e664afa04d1d141fa659bef61e3f5eaea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75ef5ffd91e1783b6f7622670bacaf71a1d2794aacba12cf3b62107d08e21b4090e63da624bb84b2e9b2c704892ade79928;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58160befe7e564958e4d6ebce0c18661ec0e527daa3d2402163a4f54385ac2ac2c2023697a6e43a23dd4df7e5efabe64a606;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66f69e0359fe98e3e609d7aff4158de765b77d5622ed154fa98c289a8095b51bb32d5fc03511c8a9da997f004f65933813e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95c4eac839603ddf003f0569326aa78cfd05750571fc92820e14b7ad0189bce27976a0a154e29ab0893fd73b7d0ba8e60d67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h231e8937a544e002e2d5b45b90cc459c3e58cc3bc1a59152618515fa9f4463b43bc4b1569933f7856f5a8c5a9b449a5d548b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h372593c27345e534de3bcd726a051b602aa4d54e4d4453dfaa7547edbc4b86efb9ca34638dcdc8a3572de676fd78bfdbf893;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31e2642cd9fab26d7db0b1266a161afcf79b6d99d8782e21af2ecffb41400a57ce5b859ee03189e0fd3c431c7fb12447ba1b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fb29a5ad9fea58020123b7e0de948d546b23239a487b86732028127002a6781c60353779fdc0e28d90400371b23434a6d1b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae2d625408d3a0b9f82f1a6ae0921941d44932753868df6d4b2aebfc34144f6d670cb399e85b7036163ddeb008546f0d911b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdda6fa72040bc1f249da71d7075d6790c9d91287685f4bf4f34d84d295b65879f8a251f5c654426fb110f751933fae9df1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71f758e55dabaed924ae684c596048ec1afd9c2ddb081b9ef58dcdd66614a56f390057c5c5edc84fcc7d2d3fd673e9374287;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he58cc71bbdd3e92046b1a6177893acef7a14e17aa4e5711cf79d0dd23dbc7acaad751ec7f29846c8d6a8d04f52b858ff8b4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87109b21a7679adcad8a5a340bcf99f2469cc9f2c3c3c8b45fb7e327ab1df1d08bf4375eea323fca867cb091691f9eed1769;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4d59ab9fdf34061a2aaf0a4485ed47adfddcbd41a201299ff500387a88dd851296cf3e4f0aada3c7a732b28bb4e8f91fb02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf96535f422bce90c742e26754686cebd3358ad0e354cfabc986e4a77454626d3010e09d9bf255b814d29acedbb47f4c2ebe8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c3e70f0f6a782a9974568ab1936bb9b39694e4edec70cc96d75a15146ac7804561e911a3d0b5ce164e801fb30038323e5e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h439942374e518a20abdabe498d0114a4fca5063703b66b4c3887840b358fd5ff43c56bfa39ebc27b29893c4c3d2dc50410c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h786bd6f9bf00cae397c2f0852694b03df4df738ddaaa08adee520041a0d856bdd12018429d447a911714fbf9a56fcf47f411;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a40173abdf6f656cf377c598beb750f7e46873acfe718712da7982afe9590a08353f1d7f2c81cebb0801a8b26154cc4c524;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f73eb554efdc40a35b6681880e2d22d1b47b151f6b713190731468955320ad537ce5ce0d5e949242cae8ecbeee392b96a94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92369bf4328764f12abc908e3ecbc4f77e356d4bf720735b895a700df60168817678585a125c574b91f9519a2c84756be8bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he97e00fa27605129d7d1e123706019dc519d9a3656322c32bf21262d0f432d8afc030395a41ce904c27ff23261c5526ccf33;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dc767e240d2a604295072710ac886b46238d34e9d3934d84e8f58fe9efd0df06357bdeeba1182bfebb29c999a12b80535f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52f22fa07917f54b3350eb6edc9d65d646461f3fedef07dd5a6e2f303324e8a50f16d4cc99c30363860c0cfa09704c113176;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbe6c737ec00c6f2b21c173a5ca2ee3ccf19bb42fac0b0ec96e3fd8eb9c400ad670be891f8e5041ad2ebd7cfd83476f4454d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he968ca0e8ccf435b92b9ccb14363313c6746d4ad6c4fba88f39d3fa44bfcd43b32212c19e853cf2f4cceeba76f534e5f4ddf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8124277a2029fc32f1138c16ac792e4a1155a73e4f22d7a47fa7c047ff573e31b11048027e23613a8f084c5a8a4e33ed4934;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d3a62221e5b1a16ba18de6a4df383aaf54d4dd666b133d2dd796bde44188d584e8f38d67304d2e35b0c11820143287bd343;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8896aabd9f39cbad830d392742b9babe27ced9e92b514265b90ed2ea9ec43120065d7395ff9e79de22bb9dc3aaa84ad216fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4ab0e256f3d946166eedfe958488f406213875296da3f74b07281aaaf948d29daef97037bff2f8c496488b9e4b612f9a23e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d5d9d2ceca9cdd9f3553503d3a236272982401e7a29cf1bf4fbedd7c43647a9168fab05838e4dae63f3940cd203471be382;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3eac3789cf8a3e88494067087b82937d2da55cdeb9890b04c8ee0676b99fb2cb93d560e17d744d4c9d899ebbc4e4fd6965b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h145c5ad4b50738453d118405194394600eb6f67285816235d37a993f3cfe30e4c9d12c0804df1f984d8c5d92de0f20460544;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe43c93031447abdc757950accd92ee13e9531c565cc8958e82d50698979b046bd23f08a82e5133d8b2535a0ec56069633c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33a9311e11c2425a580ae2b7d099571f487912b07f5850bda3d9cc65f029d348437b706ff556a128ed13b48d374ab8e4e5ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55d3099da0900dd64fc47fd50468b0f2aeac5bf529855109ee8101d96c76fac8d9d5577ab388c4376facc90a1157fd7d0b0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6db830c18213ec24a50857fed7d1512d49c3d0e41e294bf207227d90cff71772cbbc70fc465ca634e9cd7039fcb9f14c8ac0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c000e1dc1597490b26ec943108fd34a38803ee3ef42aacee365a14300317c62d581a74e69372ea9446760656d70ed31c679;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57ca25d2b4a769a2f7cdb069b1a974ee02c5dc23113a808d58629eea44735f88fc4de0a9c2e3645c69de3eae05e58a9d2b2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a6e74f0ca8f7a10e6776965cca920ed7fb780d4c825571723c03f9d9f8fb4e1bba1f352a248782ae36c77cfae740d1ada94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a515aa020ec14672164948e0896bb72c5945b33926b7b01efc53b74c7f7aa61ecc49ec94a34f831b6842d706ccddc84abba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d8fbefb3fbdc0043b792bed775dcb0ad96e0e8e8ec99e476c446a55100e1dbebeb1bff1560f8006742941e1a729304a264;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heff51b6238e204fc4b005a6da4a2b1dabc7ca29deaa66595d49f6b46f25f307acf757d5e571a23fccf9df47ea06704b1a82f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6dfcf4d446c13ded8f4119555a106f2831191327c13ab887efc5e9bac1fe52d8c380317a7a1aebb897943db561127f92c171;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea27db270b9c624b73547db21052282ba9adbf8dec61954f57aa2899863e70be57148b61a03bb0661ba8a3487e0b74cd8bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47f72d34e8432f97753080c1733e7f7664f53b88e1217610f3476940557a058a04cd88a5161e6b10f603481ce3994b760ebf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdcfa9d65d5c506bef51253ebeb559c1bd861c4e1c4ed7384ebe7dee70df0429a874a5dd72bdd0a0ee84a0b8a6964c2cff2c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb35f3793d5795bc76c56ccc187389af2cb6471644b43b86b7c234029e58f6ae2c4b8bed62122d7c4321967223d87a45c8540;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h764f8e5bcf9b24e6a050954e192477c140ea81bbc1e62488933d832a28a22394cc95d1b436e697933fcbae527db025f64f1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5dc9141bc67215ed5321f864a12902e23e60e95837a40c9493bebf3d6756673c7eea7f3b63434f6f5f5e5ca3ac402ad964e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99f4f2c9b98a08c3fca5475a8ebd2e4a42001f8a1680f5a243f9934065fefd7c4fe1c5ff0aa4e2dd1e4589899095cf987380;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f4e5237e8d9f7026b73d8f66bb31fe0d5f2e9c1d60cea3e6dbcc5c0aa288df64e258b133a983e23e93bd24d686e56e3ba28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4a59b2799ac9f59dd2fca9f72b629cd86895a172ac4ba98a0b141bfa3cf17f1830a1445fda6d520c07726f83bbd01406602;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc9c115509602f96a5a20e3f7d34baece3fe6f91b8325c02fe9b7319dfb4cbcc6ff35117e8ba281f8d0f131f394bf0740f88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a2819ea5fec8fda8cb7b472444d0a406ecbc40f70f0667e1ea1ba3bc10aca0292ccf3cce0896dc2ffd789dd0c0a6430fb62;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521103f0db187f61d22d953b38a91fdb2c9b3df866cc4dee189e6e6bfc79b2508312f5497fe5cce3d5dc610dc5d5c743dfc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h526e5d9399541211fa6c659474aec60a967367e681195382438f9cce2affc7c069cb6ecc768631d7d34e907c4f882fa6bf8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1874c749175c97affa3fc74e7c77e925936751a105770c18591e6c1843c5b7f7b8c98841ea755f4032d5343173f95189371e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h200c4e9d95238af8610f98a5bac2062eb23727379d37a4c90b8666aa997a131b281c9c56132e955750cb08a7f8a9609e5916;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h597afae6c3ec2001a3147b04bfdeb1fb23880b3aeb11ce0a36530d9cb3c43e478df7fc066928048e141b74c44c21104b824f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84f169bf048abb28b282f36908136f8771bcbce581fafcad248d5fdef4d1fac7cb59cc86f8a934ef265381b3b2fcdda7ce2d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha32a83ccdddb6809f199b03f094e012fc03f96a531023c95c00eb1c1dd610fbca1d24d58ac1e8459cb9d0b292fdce24886cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3e1bb122c05d2d3c22c882df45db57255c24fbe592ed550c27e383239bcdb8e5042d89d362af7da80a18c5b3cb96e34db90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc734c898c9508181f81ae4a12dad4afb4b93133ff12393e7f8050d1e1873f43db2f3ce371d76aafc2c057e9d0421c5131f36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee401557a71fc09befc844a66cf6371d5a4bada9e023049c879a1dc244771dc809f7d2ee70dd2abdf35c062f5d7d0d5a6628;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cda66a2ea5236efb98eb7239a04e7880013f83b1eed317a6e348aaaef91899228822414f4a75d2da2ad43ee19372e9d7f5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef9ad31d9d1a1163dc97779fc1b89efabe47fcf8d5ba42ab5a0e6ac0812d0d7e805fa7952f62b902ea25740c46b8e44c6d34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf8758de17b9287023ba874c9d4523c1958f38551af6315d8ff000684f1518288e0eb666b0bac29fc71f54a00d645eacd4bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a0f8ba707b0874a4b46e5ceeb1da53723fce7c0a35faa8769d3c21d46db662f50d2d28372ea66a1704b95ada7fe2c204399;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb3c47d30cb44b7ee544a0dbf2d427969e8d3e1c417d808e4b2119182907e20b9039449b3cde120c5572b3d4f2f318a2fa89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e72410dfd299760aff15d18dadda8301d79324066a19f1e0b6353f995f32ab5d7bae1ba7806cf9e58a6efa6b33fea57e57f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h348ecbd7649151276bcc4f0e92525be80ca9f64c40bff5600b17237eb51d874668f96f8294997bb178f636166a87d6b678ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha58040e5ba1e879937137c22c713f02e428cb1dfff7f14c06d2daa860cc216c4b10bb611f6520f8d66e05ed89e8ded86c119;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6cd772847bbd330a35734c0efb50124547d176dc9c137d9761202c045f6a6dd42ac0d225cff277b27350005b8e3554a8656;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc37e3145ed4d8169b365524c908f8e569c93559e6259a9fe99d20562f7c4c97760169044d702be028e3dd433cbff2b51217c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18f5cc4179ae93105fd97b13fac4df660e536984cb2c6bb4dcd1c93444df0d91bef6ad51f7d3ac1944209f5af93bf96d1450;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2add2a5546c8297029a01409da53207318222fab6fe59143cb9a6fc5971f892ff8a170e0dcb8beed7137929f61ab8599c72d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb85ab202821d9b1390a34f1ba97ca798445026b7ad2d6a7b32b0dac90624399c9dc62ef6876b8e20a243d65f8c1e49dea7dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5537715fb5c462214f8dea1c10c9a02512491d94f96c8e48df5fb5ed2b289edab64888f1ceaea97141e63f429a6753046a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6062425931a753d9a9f3728f2b1e1d78a7cb962ef997863d35557d6b139842381714e8a8ab9f510d150553101a00a20b3b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5451d5a91b22ea05a6f79201c32e348188a9e84d73b0a2c6eab0ee90eb863a1b648f94fd248ac8eba53825cfbeb87e9ddc04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1f1df8be27989865c42225d3f3f103e61e9370b8b57e16656fa9768dfd1d45b795d4a1b3a4209e7f93f1a76eea7bc999857;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc90317c3d665b58f477ab7a1b3fde6e5bcbc134da2dab25b2288c1ee0215d65933632b7a78a1db1a614a7923428713adc006;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e139101fc13acf82921907d4f42ad349cab0bd48056a577e8d5c80d81fd8d79f71d75300de0e5bf460442f2f9eeb3994c35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc147dfc9e7b2c311816077d926791756d3cedad01f16c042bf3aa15a418efc8de955606cca11a99dc1c3c710fdcb3bc8d9fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dc65ff15b59aeca32bc9419ad28ed38be85720f7b2a04ef75ecb0e4aff73f39a59d19eebcdccb153e64d006dbe0affa3dd4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5df7696a48fb1b1c85d540bad403b740f0d4d4a438551d34d0fcea7ba1a0ccacf96da2e4799676501f412d69d894b81cbfc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e074028eeabe4ff8daa840c2e6f882b707850091f6166d63d6dbb45820e083c8e90c6e439f24110327ad3cf417399034409;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1677b5ff45c39b61c17e74d2485fff8c645f0b53b085b42f553b32c4e0da5ee388366c93eb9d2b2e489f3b9a2263394b7259;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d303f799763704f4e017918919ebb32a2af1ed04bc74c4556f7840e6d708ee4feac820e8a69e4fe8c142881e1fdd2e40678;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e3bdd81a114d0f051707a9030fcfb68ce6776a7d3f34ccbd5ab20e192e860b6bc1f5ab8fa3640ff0fc38b48ccb9c17be949;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57e637df389dbfc2dfbee6182a4b865e77f28a9a2862ec709f565febeef6d80f682e72770a9670ba5236ef337af21cfbf14b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb03669a188de956b1e50237cc40a9d7ce46637356c58c81707b0e60e7949d34807565c03790dc0d4c55b282acee7986325b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h789a814324c3a9e118deb377de83e71cf722886447c9491a87c139ac75e985aff549a5cc90f4656bb35ddbe89b6c26795ad9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha380610abc7e628c152c6ade2c08c2b6899fd9aa2e139a56b35435c35843ddfba17a9e5fb6ec069dcca77d9543d16cde5472;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97d6c93c0f46488ae4a36dd5c6c07ce45cf1311285c3f1fcffa90c197d32f21b996fa232f9ccca189f46322a9e277fd68e13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he71eb37fbe642dff6cca7816be120e3cc689c871a97d50cfcd3dc090ae2e53517f840b120a07227b2d2acbd1a2ce4dad1154;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e967157b650404e314ef35bbabf5d5b961362bb33737f892672fa3af4312ed23a0e5950dd364ca19ffa157930ad2042831;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he771a352a380e9999347f9ea76c96d74525e300ccaa6dba2d8247d539f9746e338c4484c0b14a62cca37f0d95db8b10d54aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h814703afa07e6e829808472f8911465571e5e0d0e7a0ba55a13beffceb5b89a2217db2a0484604e5390587291701b7e01ddb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd470f4a2cfb8ff24967bbdf9b8069b3a1da89f5a14ef56c1220504a2876bc3c67259ba465644ecd3382706578182e2e5dff8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9738bac97dd6e39e1dae9cbe81a673e5fcdfc790785033eda2ce8648674cd49e8d4ffeb8b49c39f16cbafd277efd4ab32a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58882cda2f36447f1ebd58b1381ea4b79c642ba82e87a2e0d1a830092f6657e0631a566efeb7cda6484c2eca9d24e62fb660;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h343b3157cdb209b2edce7125456985296a4c9d9c753ccf5d89be77ee1b5c43009a1b8220b6c95d15d81acbaef449e0e52024;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4da98fbaa074e1a55bfa814465d35f4f4ce009edfd07128b76df1593dbab9a950f3a50f5f7b795050bcf90ae5bb25bc0c79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29e33e614595aa26a2800233793d503a0c1d6883b35a47bbf6ca1c9257ec435cb20bf715bb993e22fb0cc303ae9f3c776e85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88940d8ec62b930f0c74b46488c529d19a8a4c0b142a8717fd15009e8eca606cb1acd02bc530d405001101d6044e36ebc109;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf973834cf2d1e79dabbe4a62527a94f57f04c425d1c48cfe42d2bec71d38e754848b24a41625b84f25831eaa481c93e0400;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29ee26aab5f0cb66cc1de6541e12e5f88482bdc395116598632535a1d9bda17e2597f49961b363a856367da9b532f9fadeee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedd2ded97d9178324f11545b160c38d25f2e3218b49aa5f54f9b44e79b2ec4134c0ee5acd786f6227f9ac9bc9b409d55309e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedd8393107424bbf0d0e6dfc2b436aac8b653c1b02a4eed090b0562e5c24143d6c234c11c1b8442c726f53301b8027abf898;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafe6c9edb1e72fc31ea064090f96c7c3c56d5a5a019b14089c02f3612f5db9766be75c035b96c86eff9f4dc20f35101e6b4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h364b67e015569c2e9e7be162d315ac427133353c7ff11f3dba3fe0f12ad5c5bca8899e99e5a54eef821017a72075b730e085;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1a7c302854f1c19ec8f690286cfb30f93b6c191e89f29e5ab1c29ff01a0bb6ce3d14d492426b42ee2dfae9017ed22e0eaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h365e1af557edae1142618388ea3477750b93f5a4f4e2ff4a0ea647d27231b21150e5b23645799ec6d554177db89c5bd8a9b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c52f81131c2d8d6d27f11a9e60427affef444b6ae1dcbaeb3e209eb7cff8b752e0bdaa456279dcc2b8f823695abe11ebd88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h911a5a25d69a29f3b613e52cc9471ff0e3b820e67538ed2b612df7e3f2df8a02c60f3815b7a73f979df0e4ab24d0427568d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha09b949917a79165e3bd7d428842a60d1d80e8afe4e135e2f9fcd22104f6490b4ba53e9b0dee4f6ea4ebbd50a38a675167ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6610c6792f9731996719260ff346fe234af4e33fc1038ded3f56ad8ba8f411cdf100f7c03755e2793c8a547cb5604f68fc5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcafc4213c13c107872f3821d4eb358f66f10c2aa36c18cf2293dacb2c3e350b22bf235eeb1ec6bfdb8a69cb26ee5dfc7ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48032e6351ad265080a68d44ca81c38601c8e3c83e6d50adb9db8169835353bd87be73a28628300006ae7f4e0c6855eea30d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf7a8a9b350a2ba3435decdacecc9457afd6c1688a1b39edeb4ed9c13c7d1decdc6a1ead10f8f20574294f3d14fd52c8b15d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h533f33c5e55589728001ad661eac04e735371a989c6f65eb92a3fb2a0411abee9c3ae5078b409e7c6a6c4a1d86998469077b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec4c0d09a698e9f288e1e9714262c01fcb043e87a4833216728a6bc2d6f1a4bd383e7a978653d14fb73606bed1108fee2230;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6c8cd71494ca5875436f2b17d9e3de243ba1bdc46ffe91952e6cd4ed5177e53b83499306a9c521b1a8f24face5b0a99eb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf105314217d10149d1b4bd5715441629f04fed9926c211680fbdfb04839e7d3891cf8a4e56e5b67c4eeeb8af66bd6254c589;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c9a585711dd1c245551da4f33156c94056619f3cece81be735a08b9947d9567c6890a3fe1bd795ce6afb5a3404190b50d6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83c0d645637cef31c4cf7afb1d8e2269123a4888d3d2ba856e7bacad1ce3002b9f824cb2647947d80e4a9f65de0e178502d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c43f021f02a798e0388363d47d086b3ee4e7c070a24bf422dcc4cd28d4d7724d5cd5543b0d6f2025c4676d4e637ec6dfb04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99295af0e8904aeb31579ebcd46febee462826257de25de2bbbb56a6960feb85e680e3bf13f57b109501dbea9f68a43d7d0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb1f18760d92383c4016fb866d8c8c906fb7ba9d59a2f75728c79b7efeacf462644a08898b6454ecf20135ba76eb5f8b96b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a54a1e29a1188a140b0e07becc03585e56f91e0841f5d65c2cb0be603d43cc3fc3b7941edc206358e0ae6b5717b0a4a320c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce685d6d5ea46593f0d1335a57578e224cced480c7ed15456b2a0fd59f7151028163176758facb9956c3c6164ac05087ba41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bfcbe5c25e184c208156ca83200baa8e413e2695a33b5ad3b33fb06f71fee53639cdd85f8076c2cb06c8c36eb1f3b7736f3;
        #1
        $finish();
    end
endmodule
