module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    compressor_CLA162_12 compressor_CLA162_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA162_12(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [0:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], 1'h0, comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [0:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [30:0] stage1_0;
   wire [52:0] stage1_1;
   wire [65:0] stage1_2;
   wire [57:0] stage1_3;
   wire [138:0] stage1_4;
   wire [67:0] stage1_5;
   wire [111:0] stage1_6;
   wire [47:0] stage1_7;
   wire [72:0] stage1_8;
   wire [78:0] stage1_9;
   wire [58:0] stage1_10;
   wire [52:0] stage1_11;
   wire [52:0] stage1_12;
   wire [26:0] stage1_13;
   wire [18:0] stage2_0;
   wire [22:0] stage2_1;
   wire [26:0] stage2_2;
   wire [32:0] stage2_3;
   wire [44:0] stage2_4;
   wire [37:0] stage2_5;
   wire [49:0] stage2_6;
   wire [33:0] stage2_7;
   wire [41:0] stage2_8;
   wire [29:0] stage2_9;
   wire [29:0] stage2_10;
   wire [24:0] stage2_11;
   wire [27:0] stage2_12;
   wire [28:0] stage2_13;
   wire [8:0] stage2_14;
   wire [2:0] stage2_15;
   wire [11:0] stage3_0;
   wire [13:0] stage3_1;
   wire [18:0] stage3_2;
   wire [14:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [17:0] stage3_6;
   wire [18:0] stage3_7;
   wire [16:0] stage3_8;
   wire [11:0] stage3_9;
   wire [13:0] stage3_10;
   wire [17:0] stage3_11;
   wire [9:0] stage3_12;
   wire [12:0] stage3_13;
   wire [10:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [15:0] stage4_2;
   wire [5:0] stage4_3;
   wire [6:0] stage4_4;
   wire [7:0] stage4_5;
   wire [5:0] stage4_6;
   wire [6:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [5:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [8:0] stage4_14;
   wire [4:0] stage4_15;
   wire [2:0] stage4_16;
   wire [0:0] stage4_17;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [5:0] stage5_8;
   wire [3:0] stage5_9;
   wire [2:0] stage5_10;
   wire [1:0] stage5_11;
   wire [2:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [4:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [0:0] stage5_18;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [0:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [0:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[12]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc615_5 gpc24 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_1[13]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc615_5 gpc25 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[14]},
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc615_5 gpc26 (
      {stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[15]},
      {stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc615_5 gpc27 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_1[16]},
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[12],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[13],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[14],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[15],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[16],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[17],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[18],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[19],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[20],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[21],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[22],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[23],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc615_5 gpc52 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[24],stage1_4[52],stage1_3[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[25],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[26],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[27],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[28],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[29],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[30],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[31],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[32],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[33],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[34],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[35],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[36],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[37],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[38],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[39],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[16],stage1_6[16],stage1_5[40]}
   );
   gpc606_5 gpc69 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[17],stage1_6[17],stage1_5[41]}
   );
   gpc606_5 gpc70 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[18],stage1_6[18],stage1_5[42]}
   );
   gpc606_5 gpc71 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[19],stage1_6[19],stage1_5[43]}
   );
   gpc606_5 gpc72 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[20],stage1_6[20],stage1_5[44]}
   );
   gpc606_5 gpc73 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[21],stage1_6[21],stage1_5[45]}
   );
   gpc606_5 gpc74 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[22],stage1_6[22],stage1_5[46]}
   );
   gpc606_5 gpc75 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[23],stage1_6[23],stage1_5[47]}
   );
   gpc606_5 gpc76 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[24],stage1_6[24],stage1_5[48]}
   );
   gpc606_5 gpc77 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[25],stage1_6[25],stage1_5[49]}
   );
   gpc606_5 gpc78 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[26],stage1_6[26],stage1_5[50]}
   );
   gpc606_5 gpc79 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[27],stage1_6[27],stage1_5[51]}
   );
   gpc606_5 gpc80 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[28],stage1_6[28],stage1_5[52]}
   );
   gpc606_5 gpc81 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[29],stage1_6[29],stage1_5[53]}
   );
   gpc606_5 gpc82 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[30],stage1_6[30],stage1_5[54]}
   );
   gpc606_5 gpc83 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[31],stage1_6[31],stage1_5[55]}
   );
   gpc606_5 gpc84 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[31],stage1_7[32],stage1_6[32],stage1_5[56]}
   );
   gpc606_5 gpc85 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[32],stage1_7[33],stage1_6[33],stage1_5[57]}
   );
   gpc606_5 gpc86 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[33],stage1_7[34],stage1_6[34],stage1_5[58]}
   );
   gpc606_5 gpc87 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[34],stage1_7[35],stage1_6[35],stage1_5[59]}
   );
   gpc606_5 gpc88 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[35],stage1_7[36],stage1_6[36],stage1_5[60]}
   );
   gpc606_5 gpc89 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[36],stage1_7[37],stage1_6[37],stage1_5[61]}
   );
   gpc606_5 gpc90 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[37],stage1_7[38],stage1_6[38],stage1_5[62]}
   );
   gpc606_5 gpc91 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[38],stage1_7[39],stage1_6[39],stage1_5[63]}
   );
   gpc615_5 gpc92 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154]},
      {stage0_6[90]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[39],stage1_7[40],stage1_6[40],stage1_5[64]}
   );
   gpc615_5 gpc93 (
      {stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159]},
      {stage0_6[91]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[40],stage1_7[41],stage1_6[41],stage1_5[65]}
   );
   gpc606_5 gpc94 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc95 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[1],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc96 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[2],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc97 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[3],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc98 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[4],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc99 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[5],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc100 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[6],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc101 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[7],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc102 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[8],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc103 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[9],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc104 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[10],stage1_9[36],stage1_8[51]}
   );
   gpc606_5 gpc105 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[11],stage1_9[37],stage1_8[52]}
   );
   gpc606_5 gpc106 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[12],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc107 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[13],stage1_9[39],stage1_8[54]}
   );
   gpc606_5 gpc108 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[14],stage1_9[40],stage1_8[55]}
   );
   gpc606_5 gpc109 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[15],stage1_9[41],stage1_8[56]}
   );
   gpc606_5 gpc110 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[16],stage1_9[42],stage1_8[57]}
   );
   gpc606_5 gpc111 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[17],stage1_9[43],stage1_8[58]}
   );
   gpc606_5 gpc112 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[18],stage1_9[44],stage1_8[59]}
   );
   gpc606_5 gpc113 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[19],stage1_9[45],stage1_8[60]}
   );
   gpc606_5 gpc114 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[20],stage1_9[46],stage1_8[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[21],stage1_10[21],stage1_9[47],stage1_8[62]}
   );
   gpc606_5 gpc116 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[22],stage1_10[22],stage1_9[48],stage1_8[63]}
   );
   gpc606_5 gpc117 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[23],stage1_10[23],stage1_9[49],stage1_8[64]}
   );
   gpc606_5 gpc118 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[24],stage1_10[24],stage1_9[50],stage1_8[65]}
   );
   gpc606_5 gpc119 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[25],stage1_10[25],stage1_9[51],stage1_8[66]}
   );
   gpc606_5 gpc120 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[26],stage1_11[26],stage1_10[26],stage1_9[52]}
   );
   gpc606_5 gpc121 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[27],stage1_11[27],stage1_10[27],stage1_9[53]}
   );
   gpc606_5 gpc122 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[28],stage1_11[28],stage1_10[28],stage1_9[54]}
   );
   gpc606_5 gpc123 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[29],stage1_11[29],stage1_10[29],stage1_9[55]}
   );
   gpc606_5 gpc124 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[30],stage1_11[30],stage1_10[30],stage1_9[56]}
   );
   gpc606_5 gpc125 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[31],stage1_11[31],stage1_10[31],stage1_9[57]}
   );
   gpc606_5 gpc126 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[32],stage1_11[32],stage1_10[32],stage1_9[58]}
   );
   gpc606_5 gpc127 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[33],stage1_11[33],stage1_10[33],stage1_9[59]}
   );
   gpc606_5 gpc128 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[34],stage1_11[34],stage1_10[34],stage1_9[60]}
   );
   gpc606_5 gpc129 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[35],stage1_11[35],stage1_10[35],stage1_9[61]}
   );
   gpc606_5 gpc130 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[36],stage1_11[36],stage1_10[36],stage1_9[62]}
   );
   gpc606_5 gpc131 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[37],stage1_11[37],stage1_10[37],stage1_9[63]}
   );
   gpc606_5 gpc132 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[38],stage1_11[38],stage1_10[38],stage1_9[64]}
   );
   gpc606_5 gpc133 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[39],stage1_11[39],stage1_10[39],stage1_9[65]}
   );
   gpc606_5 gpc134 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[40],stage1_11[40],stage1_10[40],stage1_9[66]}
   );
   gpc606_5 gpc135 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[41],stage1_11[41],stage1_10[41],stage1_9[67]}
   );
   gpc606_5 gpc136 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[42],stage1_11[42],stage1_10[42],stage1_9[68]}
   );
   gpc606_5 gpc137 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[43],stage1_11[43],stage1_10[43],stage1_9[69]}
   );
   gpc606_5 gpc138 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[44],stage1_11[44],stage1_10[44],stage1_9[70]}
   );
   gpc606_5 gpc139 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[45],stage1_11[45],stage1_10[45],stage1_9[71]}
   );
   gpc606_5 gpc140 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[46],stage1_11[46],stage1_10[46],stage1_9[72]}
   );
   gpc606_5 gpc141 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[47],stage1_11[47],stage1_10[47],stage1_9[73]}
   );
   gpc606_5 gpc142 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[48],stage1_11[48],stage1_10[48],stage1_9[74]}
   );
   gpc606_5 gpc143 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[49],stage1_11[49],stage1_10[49],stage1_9[75]}
   );
   gpc606_5 gpc144 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[50],stage1_11[50],stage1_10[50],stage1_9[76]}
   );
   gpc606_5 gpc145 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[51],stage1_11[51],stage1_10[51],stage1_9[77]}
   );
   gpc606_5 gpc146 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[52],stage1_11[52],stage1_10[52],stage1_9[78]}
   );
   gpc1_1 gpc147 (
      {stage0_0[159]},
      {stage1_0[28]}
   );
   gpc1_1 gpc148 (
      {stage0_0[160]},
      {stage1_0[29]}
   );
   gpc1_1 gpc149 (
      {stage0_0[161]},
      {stage1_0[30]}
   );
   gpc1_1 gpc150 (
      {stage0_1[161]},
      {stage1_1[52]}
   );
   gpc1_1 gpc151 (
      {stage0_2[148]},
      {stage1_2[52]}
   );
   gpc1_1 gpc152 (
      {stage0_2[149]},
      {stage1_2[53]}
   );
   gpc1_1 gpc153 (
      {stage0_2[150]},
      {stage1_2[54]}
   );
   gpc1_1 gpc154 (
      {stage0_2[151]},
      {stage1_2[55]}
   );
   gpc1_1 gpc155 (
      {stage0_2[152]},
      {stage1_2[56]}
   );
   gpc1_1 gpc156 (
      {stage0_2[153]},
      {stage1_2[57]}
   );
   gpc1_1 gpc157 (
      {stage0_2[154]},
      {stage1_2[58]}
   );
   gpc1_1 gpc158 (
      {stage0_2[155]},
      {stage1_2[59]}
   );
   gpc1_1 gpc159 (
      {stage0_2[156]},
      {stage1_2[60]}
   );
   gpc1_1 gpc160 (
      {stage0_2[157]},
      {stage1_2[61]}
   );
   gpc1_1 gpc161 (
      {stage0_2[158]},
      {stage1_2[62]}
   );
   gpc1_1 gpc162 (
      {stage0_2[159]},
      {stage1_2[63]}
   );
   gpc1_1 gpc163 (
      {stage0_2[160]},
      {stage1_2[64]}
   );
   gpc1_1 gpc164 (
      {stage0_2[161]},
      {stage1_2[65]}
   );
   gpc1_1 gpc165 (
      {stage0_3[157]},
      {stage1_3[53]}
   );
   gpc1_1 gpc166 (
      {stage0_3[158]},
      {stage1_3[54]}
   );
   gpc1_1 gpc167 (
      {stage0_3[159]},
      {stage1_3[55]}
   );
   gpc1_1 gpc168 (
      {stage0_3[160]},
      {stage1_3[56]}
   );
   gpc1_1 gpc169 (
      {stage0_3[161]},
      {stage1_3[57]}
   );
   gpc1_1 gpc170 (
      {stage0_4[91]},
      {stage1_4[68]}
   );
   gpc1_1 gpc171 (
      {stage0_4[92]},
      {stage1_4[69]}
   );
   gpc1_1 gpc172 (
      {stage0_4[93]},
      {stage1_4[70]}
   );
   gpc1_1 gpc173 (
      {stage0_4[94]},
      {stage1_4[71]}
   );
   gpc1_1 gpc174 (
      {stage0_4[95]},
      {stage1_4[72]}
   );
   gpc1_1 gpc175 (
      {stage0_4[96]},
      {stage1_4[73]}
   );
   gpc1_1 gpc176 (
      {stage0_4[97]},
      {stage1_4[74]}
   );
   gpc1_1 gpc177 (
      {stage0_4[98]},
      {stage1_4[75]}
   );
   gpc1_1 gpc178 (
      {stage0_4[99]},
      {stage1_4[76]}
   );
   gpc1_1 gpc179 (
      {stage0_4[100]},
      {stage1_4[77]}
   );
   gpc1_1 gpc180 (
      {stage0_4[101]},
      {stage1_4[78]}
   );
   gpc1_1 gpc181 (
      {stage0_4[102]},
      {stage1_4[79]}
   );
   gpc1_1 gpc182 (
      {stage0_4[103]},
      {stage1_4[80]}
   );
   gpc1_1 gpc183 (
      {stage0_4[104]},
      {stage1_4[81]}
   );
   gpc1_1 gpc184 (
      {stage0_4[105]},
      {stage1_4[82]}
   );
   gpc1_1 gpc185 (
      {stage0_4[106]},
      {stage1_4[83]}
   );
   gpc1_1 gpc186 (
      {stage0_4[107]},
      {stage1_4[84]}
   );
   gpc1_1 gpc187 (
      {stage0_4[108]},
      {stage1_4[85]}
   );
   gpc1_1 gpc188 (
      {stage0_4[109]},
      {stage1_4[86]}
   );
   gpc1_1 gpc189 (
      {stage0_4[110]},
      {stage1_4[87]}
   );
   gpc1_1 gpc190 (
      {stage0_4[111]},
      {stage1_4[88]}
   );
   gpc1_1 gpc191 (
      {stage0_4[112]},
      {stage1_4[89]}
   );
   gpc1_1 gpc192 (
      {stage0_4[113]},
      {stage1_4[90]}
   );
   gpc1_1 gpc193 (
      {stage0_4[114]},
      {stage1_4[91]}
   );
   gpc1_1 gpc194 (
      {stage0_4[115]},
      {stage1_4[92]}
   );
   gpc1_1 gpc195 (
      {stage0_4[116]},
      {stage1_4[93]}
   );
   gpc1_1 gpc196 (
      {stage0_4[117]},
      {stage1_4[94]}
   );
   gpc1_1 gpc197 (
      {stage0_4[118]},
      {stage1_4[95]}
   );
   gpc1_1 gpc198 (
      {stage0_4[119]},
      {stage1_4[96]}
   );
   gpc1_1 gpc199 (
      {stage0_4[120]},
      {stage1_4[97]}
   );
   gpc1_1 gpc200 (
      {stage0_4[121]},
      {stage1_4[98]}
   );
   gpc1_1 gpc201 (
      {stage0_4[122]},
      {stage1_4[99]}
   );
   gpc1_1 gpc202 (
      {stage0_4[123]},
      {stage1_4[100]}
   );
   gpc1_1 gpc203 (
      {stage0_4[124]},
      {stage1_4[101]}
   );
   gpc1_1 gpc204 (
      {stage0_4[125]},
      {stage1_4[102]}
   );
   gpc1_1 gpc205 (
      {stage0_4[126]},
      {stage1_4[103]}
   );
   gpc1_1 gpc206 (
      {stage0_4[127]},
      {stage1_4[104]}
   );
   gpc1_1 gpc207 (
      {stage0_4[128]},
      {stage1_4[105]}
   );
   gpc1_1 gpc208 (
      {stage0_4[129]},
      {stage1_4[106]}
   );
   gpc1_1 gpc209 (
      {stage0_4[130]},
      {stage1_4[107]}
   );
   gpc1_1 gpc210 (
      {stage0_4[131]},
      {stage1_4[108]}
   );
   gpc1_1 gpc211 (
      {stage0_4[132]},
      {stage1_4[109]}
   );
   gpc1_1 gpc212 (
      {stage0_4[133]},
      {stage1_4[110]}
   );
   gpc1_1 gpc213 (
      {stage0_4[134]},
      {stage1_4[111]}
   );
   gpc1_1 gpc214 (
      {stage0_4[135]},
      {stage1_4[112]}
   );
   gpc1_1 gpc215 (
      {stage0_4[136]},
      {stage1_4[113]}
   );
   gpc1_1 gpc216 (
      {stage0_4[137]},
      {stage1_4[114]}
   );
   gpc1_1 gpc217 (
      {stage0_4[138]},
      {stage1_4[115]}
   );
   gpc1_1 gpc218 (
      {stage0_4[139]},
      {stage1_4[116]}
   );
   gpc1_1 gpc219 (
      {stage0_4[140]},
      {stage1_4[117]}
   );
   gpc1_1 gpc220 (
      {stage0_4[141]},
      {stage1_4[118]}
   );
   gpc1_1 gpc221 (
      {stage0_4[142]},
      {stage1_4[119]}
   );
   gpc1_1 gpc222 (
      {stage0_4[143]},
      {stage1_4[120]}
   );
   gpc1_1 gpc223 (
      {stage0_4[144]},
      {stage1_4[121]}
   );
   gpc1_1 gpc224 (
      {stage0_4[145]},
      {stage1_4[122]}
   );
   gpc1_1 gpc225 (
      {stage0_4[146]},
      {stage1_4[123]}
   );
   gpc1_1 gpc226 (
      {stage0_4[147]},
      {stage1_4[124]}
   );
   gpc1_1 gpc227 (
      {stage0_4[148]},
      {stage1_4[125]}
   );
   gpc1_1 gpc228 (
      {stage0_4[149]},
      {stage1_4[126]}
   );
   gpc1_1 gpc229 (
      {stage0_4[150]},
      {stage1_4[127]}
   );
   gpc1_1 gpc230 (
      {stage0_4[151]},
      {stage1_4[128]}
   );
   gpc1_1 gpc231 (
      {stage0_4[152]},
      {stage1_4[129]}
   );
   gpc1_1 gpc232 (
      {stage0_4[153]},
      {stage1_4[130]}
   );
   gpc1_1 gpc233 (
      {stage0_4[154]},
      {stage1_4[131]}
   );
   gpc1_1 gpc234 (
      {stage0_4[155]},
      {stage1_4[132]}
   );
   gpc1_1 gpc235 (
      {stage0_4[156]},
      {stage1_4[133]}
   );
   gpc1_1 gpc236 (
      {stage0_4[157]},
      {stage1_4[134]}
   );
   gpc1_1 gpc237 (
      {stage0_4[158]},
      {stage1_4[135]}
   );
   gpc1_1 gpc238 (
      {stage0_4[159]},
      {stage1_4[136]}
   );
   gpc1_1 gpc239 (
      {stage0_4[160]},
      {stage1_4[137]}
   );
   gpc1_1 gpc240 (
      {stage0_4[161]},
      {stage1_4[138]}
   );
   gpc1_1 gpc241 (
      {stage0_5[160]},
      {stage1_5[66]}
   );
   gpc1_1 gpc242 (
      {stage0_5[161]},
      {stage1_5[67]}
   );
   gpc1_1 gpc243 (
      {stage0_6[92]},
      {stage1_6[42]}
   );
   gpc1_1 gpc244 (
      {stage0_6[93]},
      {stage1_6[43]}
   );
   gpc1_1 gpc245 (
      {stage0_6[94]},
      {stage1_6[44]}
   );
   gpc1_1 gpc246 (
      {stage0_6[95]},
      {stage1_6[45]}
   );
   gpc1_1 gpc247 (
      {stage0_6[96]},
      {stage1_6[46]}
   );
   gpc1_1 gpc248 (
      {stage0_6[97]},
      {stage1_6[47]}
   );
   gpc1_1 gpc249 (
      {stage0_6[98]},
      {stage1_6[48]}
   );
   gpc1_1 gpc250 (
      {stage0_6[99]},
      {stage1_6[49]}
   );
   gpc1_1 gpc251 (
      {stage0_6[100]},
      {stage1_6[50]}
   );
   gpc1_1 gpc252 (
      {stage0_6[101]},
      {stage1_6[51]}
   );
   gpc1_1 gpc253 (
      {stage0_6[102]},
      {stage1_6[52]}
   );
   gpc1_1 gpc254 (
      {stage0_6[103]},
      {stage1_6[53]}
   );
   gpc1_1 gpc255 (
      {stage0_6[104]},
      {stage1_6[54]}
   );
   gpc1_1 gpc256 (
      {stage0_6[105]},
      {stage1_6[55]}
   );
   gpc1_1 gpc257 (
      {stage0_6[106]},
      {stage1_6[56]}
   );
   gpc1_1 gpc258 (
      {stage0_6[107]},
      {stage1_6[57]}
   );
   gpc1_1 gpc259 (
      {stage0_6[108]},
      {stage1_6[58]}
   );
   gpc1_1 gpc260 (
      {stage0_6[109]},
      {stage1_6[59]}
   );
   gpc1_1 gpc261 (
      {stage0_6[110]},
      {stage1_6[60]}
   );
   gpc1_1 gpc262 (
      {stage0_6[111]},
      {stage1_6[61]}
   );
   gpc1_1 gpc263 (
      {stage0_6[112]},
      {stage1_6[62]}
   );
   gpc1_1 gpc264 (
      {stage0_6[113]},
      {stage1_6[63]}
   );
   gpc1_1 gpc265 (
      {stage0_6[114]},
      {stage1_6[64]}
   );
   gpc1_1 gpc266 (
      {stage0_6[115]},
      {stage1_6[65]}
   );
   gpc1_1 gpc267 (
      {stage0_6[116]},
      {stage1_6[66]}
   );
   gpc1_1 gpc268 (
      {stage0_6[117]},
      {stage1_6[67]}
   );
   gpc1_1 gpc269 (
      {stage0_6[118]},
      {stage1_6[68]}
   );
   gpc1_1 gpc270 (
      {stage0_6[119]},
      {stage1_6[69]}
   );
   gpc1_1 gpc271 (
      {stage0_6[120]},
      {stage1_6[70]}
   );
   gpc1_1 gpc272 (
      {stage0_6[121]},
      {stage1_6[71]}
   );
   gpc1_1 gpc273 (
      {stage0_6[122]},
      {stage1_6[72]}
   );
   gpc1_1 gpc274 (
      {stage0_6[123]},
      {stage1_6[73]}
   );
   gpc1_1 gpc275 (
      {stage0_6[124]},
      {stage1_6[74]}
   );
   gpc1_1 gpc276 (
      {stage0_6[125]},
      {stage1_6[75]}
   );
   gpc1_1 gpc277 (
      {stage0_6[126]},
      {stage1_6[76]}
   );
   gpc1_1 gpc278 (
      {stage0_6[127]},
      {stage1_6[77]}
   );
   gpc1_1 gpc279 (
      {stage0_6[128]},
      {stage1_6[78]}
   );
   gpc1_1 gpc280 (
      {stage0_6[129]},
      {stage1_6[79]}
   );
   gpc1_1 gpc281 (
      {stage0_6[130]},
      {stage1_6[80]}
   );
   gpc1_1 gpc282 (
      {stage0_6[131]},
      {stage1_6[81]}
   );
   gpc1_1 gpc283 (
      {stage0_6[132]},
      {stage1_6[82]}
   );
   gpc1_1 gpc284 (
      {stage0_6[133]},
      {stage1_6[83]}
   );
   gpc1_1 gpc285 (
      {stage0_6[134]},
      {stage1_6[84]}
   );
   gpc1_1 gpc286 (
      {stage0_6[135]},
      {stage1_6[85]}
   );
   gpc1_1 gpc287 (
      {stage0_6[136]},
      {stage1_6[86]}
   );
   gpc1_1 gpc288 (
      {stage0_6[137]},
      {stage1_6[87]}
   );
   gpc1_1 gpc289 (
      {stage0_6[138]},
      {stage1_6[88]}
   );
   gpc1_1 gpc290 (
      {stage0_6[139]},
      {stage1_6[89]}
   );
   gpc1_1 gpc291 (
      {stage0_6[140]},
      {stage1_6[90]}
   );
   gpc1_1 gpc292 (
      {stage0_6[141]},
      {stage1_6[91]}
   );
   gpc1_1 gpc293 (
      {stage0_6[142]},
      {stage1_6[92]}
   );
   gpc1_1 gpc294 (
      {stage0_6[143]},
      {stage1_6[93]}
   );
   gpc1_1 gpc295 (
      {stage0_6[144]},
      {stage1_6[94]}
   );
   gpc1_1 gpc296 (
      {stage0_6[145]},
      {stage1_6[95]}
   );
   gpc1_1 gpc297 (
      {stage0_6[146]},
      {stage1_6[96]}
   );
   gpc1_1 gpc298 (
      {stage0_6[147]},
      {stage1_6[97]}
   );
   gpc1_1 gpc299 (
      {stage0_6[148]},
      {stage1_6[98]}
   );
   gpc1_1 gpc300 (
      {stage0_6[149]},
      {stage1_6[99]}
   );
   gpc1_1 gpc301 (
      {stage0_6[150]},
      {stage1_6[100]}
   );
   gpc1_1 gpc302 (
      {stage0_6[151]},
      {stage1_6[101]}
   );
   gpc1_1 gpc303 (
      {stage0_6[152]},
      {stage1_6[102]}
   );
   gpc1_1 gpc304 (
      {stage0_6[153]},
      {stage1_6[103]}
   );
   gpc1_1 gpc305 (
      {stage0_6[154]},
      {stage1_6[104]}
   );
   gpc1_1 gpc306 (
      {stage0_6[155]},
      {stage1_6[105]}
   );
   gpc1_1 gpc307 (
      {stage0_6[156]},
      {stage1_6[106]}
   );
   gpc1_1 gpc308 (
      {stage0_6[157]},
      {stage1_6[107]}
   );
   gpc1_1 gpc309 (
      {stage0_6[158]},
      {stage1_6[108]}
   );
   gpc1_1 gpc310 (
      {stage0_6[159]},
      {stage1_6[109]}
   );
   gpc1_1 gpc311 (
      {stage0_6[160]},
      {stage1_6[110]}
   );
   gpc1_1 gpc312 (
      {stage0_6[161]},
      {stage1_6[111]}
   );
   gpc1_1 gpc313 (
      {stage0_7[156]},
      {stage1_7[42]}
   );
   gpc1_1 gpc314 (
      {stage0_7[157]},
      {stage1_7[43]}
   );
   gpc1_1 gpc315 (
      {stage0_7[158]},
      {stage1_7[44]}
   );
   gpc1_1 gpc316 (
      {stage0_7[159]},
      {stage1_7[45]}
   );
   gpc1_1 gpc317 (
      {stage0_7[160]},
      {stage1_7[46]}
   );
   gpc1_1 gpc318 (
      {stage0_7[161]},
      {stage1_7[47]}
   );
   gpc1_1 gpc319 (
      {stage0_8[156]},
      {stage1_8[67]}
   );
   gpc1_1 gpc320 (
      {stage0_8[157]},
      {stage1_8[68]}
   );
   gpc1_1 gpc321 (
      {stage0_8[158]},
      {stage1_8[69]}
   );
   gpc1_1 gpc322 (
      {stage0_8[159]},
      {stage1_8[70]}
   );
   gpc1_1 gpc323 (
      {stage0_8[160]},
      {stage1_8[71]}
   );
   gpc1_1 gpc324 (
      {stage0_8[161]},
      {stage1_8[72]}
   );
   gpc1_1 gpc325 (
      {stage0_10[156]},
      {stage1_10[53]}
   );
   gpc1_1 gpc326 (
      {stage0_10[157]},
      {stage1_10[54]}
   );
   gpc1_1 gpc327 (
      {stage0_10[158]},
      {stage1_10[55]}
   );
   gpc1_1 gpc328 (
      {stage0_10[159]},
      {stage1_10[56]}
   );
   gpc1_1 gpc329 (
      {stage0_10[160]},
      {stage1_10[57]}
   );
   gpc1_1 gpc330 (
      {stage0_10[161]},
      {stage1_10[58]}
   );
   gpc1163_5 gpc331 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc332 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc333 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc334 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc335 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc336 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc337 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc338 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc339 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc606_5 gpc340 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc341 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc606_5 gpc342 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc606_5 gpc343 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc344 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52]},
      {stage1_3[6]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc345 (
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[8],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc346 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[9],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc347 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[10],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc348 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[11],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc349 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[12],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc350 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[13],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc351 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[14],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc352 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[15],stage2_4[21],stage2_3[21]}
   );
   gpc606_5 gpc353 (
      {stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[8],stage2_6[16],stage2_5[16],stage2_4[22]}
   );
   gpc606_5 gpc354 (
      {stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[9],stage2_6[17],stage2_5[17],stage2_4[23]}
   );
   gpc606_5 gpc355 (
      {stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[10],stage2_6[18],stage2_5[18],stage2_4[24]}
   );
   gpc606_5 gpc356 (
      {stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[11],stage2_6[19],stage2_5[19],stage2_4[25]}
   );
   gpc606_5 gpc357 (
      {stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[12],stage2_6[20],stage2_5[20],stage2_4[26]}
   );
   gpc606_5 gpc358 (
      {stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[13],stage2_6[21],stage2_5[21],stage2_4[27]}
   );
   gpc606_5 gpc359 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[14],stage2_6[22],stage2_5[22],stage2_4[28]}
   );
   gpc606_5 gpc360 (
      {stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[15],stage2_6[23],stage2_5[23],stage2_4[29]}
   );
   gpc606_5 gpc361 (
      {stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[16],stage2_6[24],stage2_5[24],stage2_4[30]}
   );
   gpc606_5 gpc362 (
      {stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[17],stage2_6[25],stage2_5[25],stage2_4[31]}
   );
   gpc606_5 gpc363 (
      {stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[18],stage2_6[26],stage2_5[26],stage2_4[32]}
   );
   gpc606_5 gpc364 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[19],stage2_6[27],stage2_5[27],stage2_4[33]}
   );
   gpc606_5 gpc365 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[12],stage2_7[20],stage2_6[28],stage2_5[28]}
   );
   gpc606_5 gpc366 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[13],stage2_7[21],stage2_6[29],stage2_5[29]}
   );
   gpc615_5 gpc367 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[12]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[14],stage2_7[22],stage2_6[30]}
   );
   gpc615_5 gpc368 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[15],stage2_7[23],stage2_6[31]}
   );
   gpc615_5 gpc369 (
      {stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85], stage1_6[86]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[16],stage2_7[24],stage2_6[32]}
   );
   gpc615_5 gpc370 (
      {stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage1_7[15]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[5],stage2_8[17],stage2_7[25],stage2_6[33]}
   );
   gpc615_5 gpc371 (
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_7[16]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[6],stage2_8[18],stage2_7[26],stage2_6[34]}
   );
   gpc615_5 gpc372 (
      {stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[7],stage2_8[19],stage2_7[27]}
   );
   gpc615_5 gpc373 (
      {stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[8],stage2_8[20],stage2_7[28]}
   );
   gpc615_5 gpc374 (
      {stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[9],stage2_8[21],stage2_7[29]}
   );
   gpc615_5 gpc375 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[10],stage2_8[22],stage2_7[30]}
   );
   gpc615_5 gpc376 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[11],stage2_8[23],stage2_7[31]}
   );
   gpc615_5 gpc377 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[12],stage2_8[24],stage2_7[32]}
   );
   gpc606_5 gpc378 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[6],stage2_10[11],stage2_9[13],stage2_8[25]}
   );
   gpc606_5 gpc379 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[7],stage2_10[12],stage2_9[14],stage2_8[26]}
   );
   gpc606_5 gpc380 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[8],stage2_10[13],stage2_9[15],stage2_8[27]}
   );
   gpc606_5 gpc381 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[9],stage2_10[14],stage2_9[16],stage2_8[28]}
   );
   gpc606_5 gpc382 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[4],stage2_11[10],stage2_10[15],stage2_9[17]}
   );
   gpc606_5 gpc383 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[5],stage2_11[11],stage2_10[16],stage2_9[18]}
   );
   gpc606_5 gpc384 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[6],stage2_11[12],stage2_10[17],stage2_9[19]}
   );
   gpc606_5 gpc385 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[7],stage2_11[13],stage2_10[18],stage2_9[20]}
   );
   gpc606_5 gpc386 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[8],stage2_11[14],stage2_10[19],stage2_9[21]}
   );
   gpc606_5 gpc387 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[9],stage2_11[15],stage2_10[20],stage2_9[22]}
   );
   gpc606_5 gpc388 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[6],stage2_12[10],stage2_11[16],stage2_10[21]}
   );
   gpc606_5 gpc389 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[7],stage2_12[11],stage2_11[17],stage2_10[22]}
   );
   gpc615_5 gpc390 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40]},
      {stage1_11[36]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[8],stage2_12[12],stage2_11[18],stage2_10[23]}
   );
   gpc615_5 gpc391 (
      {stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45]},
      {stage1_11[37]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[9],stage2_12[13],stage2_11[19],stage2_10[24]}
   );
   gpc615_5 gpc392 (
      {stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[38]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[10],stage2_12[14],stage2_11[20],stage2_10[25]}
   );
   gpc615_5 gpc393 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage1_11[39]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[11],stage2_12[15],stage2_11[21],stage2_10[26]}
   );
   gpc1163_5 gpc394 (
      {stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[0]},
      {1'b0},
      {stage2_15[0],stage2_14[6],stage2_13[12],stage2_12[16],stage2_11[22]}
   );
   gpc615_5 gpc395 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_12[42]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[1],stage2_14[7],stage2_13[13],stage2_12[17],stage2_11[23]}
   );
   gpc615_5 gpc396 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[43]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12]},
      {stage2_15[2],stage2_14[8],stage2_13[14],stage2_12[18],stage2_11[24]}
   );
   gpc1_1 gpc397 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc398 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc399 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc400 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc401 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc402 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc403 (
      {stage1_0[24]},
      {stage2_0[12]}
   );
   gpc1_1 gpc404 (
      {stage1_0[25]},
      {stage2_0[13]}
   );
   gpc1_1 gpc405 (
      {stage1_0[26]},
      {stage2_0[14]}
   );
   gpc1_1 gpc406 (
      {stage1_0[27]},
      {stage2_0[15]}
   );
   gpc1_1 gpc407 (
      {stage1_0[28]},
      {stage2_0[16]}
   );
   gpc1_1 gpc408 (
      {stage1_0[29]},
      {stage2_0[17]}
   );
   gpc1_1 gpc409 (
      {stage1_0[30]},
      {stage2_0[18]}
   );
   gpc1_1 gpc410 (
      {stage1_1[36]},
      {stage2_1[6]}
   );
   gpc1_1 gpc411 (
      {stage1_1[37]},
      {stage2_1[7]}
   );
   gpc1_1 gpc412 (
      {stage1_1[38]},
      {stage2_1[8]}
   );
   gpc1_1 gpc413 (
      {stage1_1[39]},
      {stage2_1[9]}
   );
   gpc1_1 gpc414 (
      {stage1_1[40]},
      {stage2_1[10]}
   );
   gpc1_1 gpc415 (
      {stage1_1[41]},
      {stage2_1[11]}
   );
   gpc1_1 gpc416 (
      {stage1_1[42]},
      {stage2_1[12]}
   );
   gpc1_1 gpc417 (
      {stage1_1[43]},
      {stage2_1[13]}
   );
   gpc1_1 gpc418 (
      {stage1_1[44]},
      {stage2_1[14]}
   );
   gpc1_1 gpc419 (
      {stage1_1[45]},
      {stage2_1[15]}
   );
   gpc1_1 gpc420 (
      {stage1_1[46]},
      {stage2_1[16]}
   );
   gpc1_1 gpc421 (
      {stage1_1[47]},
      {stage2_1[17]}
   );
   gpc1_1 gpc422 (
      {stage1_1[48]},
      {stage2_1[18]}
   );
   gpc1_1 gpc423 (
      {stage1_1[49]},
      {stage2_1[19]}
   );
   gpc1_1 gpc424 (
      {stage1_1[50]},
      {stage2_1[20]}
   );
   gpc1_1 gpc425 (
      {stage1_1[51]},
      {stage2_1[21]}
   );
   gpc1_1 gpc426 (
      {stage1_1[52]},
      {stage2_1[22]}
   );
   gpc1_1 gpc427 (
      {stage1_2[53]},
      {stage2_2[14]}
   );
   gpc1_1 gpc428 (
      {stage1_2[54]},
      {stage2_2[15]}
   );
   gpc1_1 gpc429 (
      {stage1_2[55]},
      {stage2_2[16]}
   );
   gpc1_1 gpc430 (
      {stage1_2[56]},
      {stage2_2[17]}
   );
   gpc1_1 gpc431 (
      {stage1_2[57]},
      {stage2_2[18]}
   );
   gpc1_1 gpc432 (
      {stage1_2[58]},
      {stage2_2[19]}
   );
   gpc1_1 gpc433 (
      {stage1_2[59]},
      {stage2_2[20]}
   );
   gpc1_1 gpc434 (
      {stage1_2[60]},
      {stage2_2[21]}
   );
   gpc1_1 gpc435 (
      {stage1_2[61]},
      {stage2_2[22]}
   );
   gpc1_1 gpc436 (
      {stage1_2[62]},
      {stage2_2[23]}
   );
   gpc1_1 gpc437 (
      {stage1_2[63]},
      {stage2_2[24]}
   );
   gpc1_1 gpc438 (
      {stage1_2[64]},
      {stage2_2[25]}
   );
   gpc1_1 gpc439 (
      {stage1_2[65]},
      {stage2_2[26]}
   );
   gpc1_1 gpc440 (
      {stage1_3[47]},
      {stage2_3[22]}
   );
   gpc1_1 gpc441 (
      {stage1_3[48]},
      {stage2_3[23]}
   );
   gpc1_1 gpc442 (
      {stage1_3[49]},
      {stage2_3[24]}
   );
   gpc1_1 gpc443 (
      {stage1_3[50]},
      {stage2_3[25]}
   );
   gpc1_1 gpc444 (
      {stage1_3[51]},
      {stage2_3[26]}
   );
   gpc1_1 gpc445 (
      {stage1_3[52]},
      {stage2_3[27]}
   );
   gpc1_1 gpc446 (
      {stage1_3[53]},
      {stage2_3[28]}
   );
   gpc1_1 gpc447 (
      {stage1_3[54]},
      {stage2_3[29]}
   );
   gpc1_1 gpc448 (
      {stage1_3[55]},
      {stage2_3[30]}
   );
   gpc1_1 gpc449 (
      {stage1_3[56]},
      {stage2_3[31]}
   );
   gpc1_1 gpc450 (
      {stage1_3[57]},
      {stage2_3[32]}
   );
   gpc1_1 gpc451 (
      {stage1_4[128]},
      {stage2_4[34]}
   );
   gpc1_1 gpc452 (
      {stage1_4[129]},
      {stage2_4[35]}
   );
   gpc1_1 gpc453 (
      {stage1_4[130]},
      {stage2_4[36]}
   );
   gpc1_1 gpc454 (
      {stage1_4[131]},
      {stage2_4[37]}
   );
   gpc1_1 gpc455 (
      {stage1_4[132]},
      {stage2_4[38]}
   );
   gpc1_1 gpc456 (
      {stage1_4[133]},
      {stage2_4[39]}
   );
   gpc1_1 gpc457 (
      {stage1_4[134]},
      {stage2_4[40]}
   );
   gpc1_1 gpc458 (
      {stage1_4[135]},
      {stage2_4[41]}
   );
   gpc1_1 gpc459 (
      {stage1_4[136]},
      {stage2_4[42]}
   );
   gpc1_1 gpc460 (
      {stage1_4[137]},
      {stage2_4[43]}
   );
   gpc1_1 gpc461 (
      {stage1_4[138]},
      {stage2_4[44]}
   );
   gpc1_1 gpc462 (
      {stage1_5[60]},
      {stage2_5[30]}
   );
   gpc1_1 gpc463 (
      {stage1_5[61]},
      {stage2_5[31]}
   );
   gpc1_1 gpc464 (
      {stage1_5[62]},
      {stage2_5[32]}
   );
   gpc1_1 gpc465 (
      {stage1_5[63]},
      {stage2_5[33]}
   );
   gpc1_1 gpc466 (
      {stage1_5[64]},
      {stage2_5[34]}
   );
   gpc1_1 gpc467 (
      {stage1_5[65]},
      {stage2_5[35]}
   );
   gpc1_1 gpc468 (
      {stage1_5[66]},
      {stage2_5[36]}
   );
   gpc1_1 gpc469 (
      {stage1_5[67]},
      {stage2_5[37]}
   );
   gpc1_1 gpc470 (
      {stage1_6[97]},
      {stage2_6[35]}
   );
   gpc1_1 gpc471 (
      {stage1_6[98]},
      {stage2_6[36]}
   );
   gpc1_1 gpc472 (
      {stage1_6[99]},
      {stage2_6[37]}
   );
   gpc1_1 gpc473 (
      {stage1_6[100]},
      {stage2_6[38]}
   );
   gpc1_1 gpc474 (
      {stage1_6[101]},
      {stage2_6[39]}
   );
   gpc1_1 gpc475 (
      {stage1_6[102]},
      {stage2_6[40]}
   );
   gpc1_1 gpc476 (
      {stage1_6[103]},
      {stage2_6[41]}
   );
   gpc1_1 gpc477 (
      {stage1_6[104]},
      {stage2_6[42]}
   );
   gpc1_1 gpc478 (
      {stage1_6[105]},
      {stage2_6[43]}
   );
   gpc1_1 gpc479 (
      {stage1_6[106]},
      {stage2_6[44]}
   );
   gpc1_1 gpc480 (
      {stage1_6[107]},
      {stage2_6[45]}
   );
   gpc1_1 gpc481 (
      {stage1_6[108]},
      {stage2_6[46]}
   );
   gpc1_1 gpc482 (
      {stage1_6[109]},
      {stage2_6[47]}
   );
   gpc1_1 gpc483 (
      {stage1_6[110]},
      {stage2_6[48]}
   );
   gpc1_1 gpc484 (
      {stage1_6[111]},
      {stage2_6[49]}
   );
   gpc1_1 gpc485 (
      {stage1_7[47]},
      {stage2_7[33]}
   );
   gpc1_1 gpc486 (
      {stage1_8[60]},
      {stage2_8[29]}
   );
   gpc1_1 gpc487 (
      {stage1_8[61]},
      {stage2_8[30]}
   );
   gpc1_1 gpc488 (
      {stage1_8[62]},
      {stage2_8[31]}
   );
   gpc1_1 gpc489 (
      {stage1_8[63]},
      {stage2_8[32]}
   );
   gpc1_1 gpc490 (
      {stage1_8[64]},
      {stage2_8[33]}
   );
   gpc1_1 gpc491 (
      {stage1_8[65]},
      {stage2_8[34]}
   );
   gpc1_1 gpc492 (
      {stage1_8[66]},
      {stage2_8[35]}
   );
   gpc1_1 gpc493 (
      {stage1_8[67]},
      {stage2_8[36]}
   );
   gpc1_1 gpc494 (
      {stage1_8[68]},
      {stage2_8[37]}
   );
   gpc1_1 gpc495 (
      {stage1_8[69]},
      {stage2_8[38]}
   );
   gpc1_1 gpc496 (
      {stage1_8[70]},
      {stage2_8[39]}
   );
   gpc1_1 gpc497 (
      {stage1_8[71]},
      {stage2_8[40]}
   );
   gpc1_1 gpc498 (
      {stage1_8[72]},
      {stage2_8[41]}
   );
   gpc1_1 gpc499 (
      {stage1_9[72]},
      {stage2_9[23]}
   );
   gpc1_1 gpc500 (
      {stage1_9[73]},
      {stage2_9[24]}
   );
   gpc1_1 gpc501 (
      {stage1_9[74]},
      {stage2_9[25]}
   );
   gpc1_1 gpc502 (
      {stage1_9[75]},
      {stage2_9[26]}
   );
   gpc1_1 gpc503 (
      {stage1_9[76]},
      {stage2_9[27]}
   );
   gpc1_1 gpc504 (
      {stage1_9[77]},
      {stage2_9[28]}
   );
   gpc1_1 gpc505 (
      {stage1_9[78]},
      {stage2_9[29]}
   );
   gpc1_1 gpc506 (
      {stage1_10[56]},
      {stage2_10[27]}
   );
   gpc1_1 gpc507 (
      {stage1_10[57]},
      {stage2_10[28]}
   );
   gpc1_1 gpc508 (
      {stage1_10[58]},
      {stage2_10[29]}
   );
   gpc1_1 gpc509 (
      {stage1_12[44]},
      {stage2_12[19]}
   );
   gpc1_1 gpc510 (
      {stage1_12[45]},
      {stage2_12[20]}
   );
   gpc1_1 gpc511 (
      {stage1_12[46]},
      {stage2_12[21]}
   );
   gpc1_1 gpc512 (
      {stage1_12[47]},
      {stage2_12[22]}
   );
   gpc1_1 gpc513 (
      {stage1_12[48]},
      {stage2_12[23]}
   );
   gpc1_1 gpc514 (
      {stage1_12[49]},
      {stage2_12[24]}
   );
   gpc1_1 gpc515 (
      {stage1_12[50]},
      {stage2_12[25]}
   );
   gpc1_1 gpc516 (
      {stage1_12[51]},
      {stage2_12[26]}
   );
   gpc1_1 gpc517 (
      {stage1_12[52]},
      {stage2_12[27]}
   );
   gpc1_1 gpc518 (
      {stage1_13[13]},
      {stage2_13[15]}
   );
   gpc1_1 gpc519 (
      {stage1_13[14]},
      {stage2_13[16]}
   );
   gpc1_1 gpc520 (
      {stage1_13[15]},
      {stage2_13[17]}
   );
   gpc1_1 gpc521 (
      {stage1_13[16]},
      {stage2_13[18]}
   );
   gpc1_1 gpc522 (
      {stage1_13[17]},
      {stage2_13[19]}
   );
   gpc1_1 gpc523 (
      {stage1_13[18]},
      {stage2_13[20]}
   );
   gpc1_1 gpc524 (
      {stage1_13[19]},
      {stage2_13[21]}
   );
   gpc1_1 gpc525 (
      {stage1_13[20]},
      {stage2_13[22]}
   );
   gpc1_1 gpc526 (
      {stage1_13[21]},
      {stage2_13[23]}
   );
   gpc1_1 gpc527 (
      {stage1_13[22]},
      {stage2_13[24]}
   );
   gpc1_1 gpc528 (
      {stage1_13[23]},
      {stage2_13[25]}
   );
   gpc1_1 gpc529 (
      {stage1_13[24]},
      {stage2_13[26]}
   );
   gpc1_1 gpc530 (
      {stage1_13[25]},
      {stage2_13[27]}
   );
   gpc1_1 gpc531 (
      {stage1_13[26]},
      {stage2_13[28]}
   );
   gpc1163_5 gpc532 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc533 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1406_5 gpc534 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc615_5 gpc535 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[5]},
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc536 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc537 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc538 (
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20]},
      {stage2_4[9]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc615_5 gpc539 (
      {stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25]},
      {stage2_4[10]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[7],stage3_3[7]}
   );
   gpc606_5 gpc540 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc541 (
      {stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc542 (
      {stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[6],stage3_6[7],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc543 (
      {stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33]},
      {stage2_5[24]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[7],stage3_6[8],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc544 (
      {stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_5[25]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[8],stage3_6[9],stage3_5[10],stage3_4[12]}
   );
   gpc606_5 gpc545 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[5],stage3_7[9],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc546 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[6],stage3_7[10],stage3_6[11]}
   );
   gpc615_5 gpc547 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[6]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[7],stage3_7[11],stage3_6[12]}
   );
   gpc615_5 gpc548 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[7]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[8],stage3_7[12],stage3_6[13]}
   );
   gpc1343_5 gpc549 (
      {stage2_7[8], stage2_7[9], stage2_7[10]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[0]},
      {stage3_11[0],stage3_10[3],stage3_9[4],stage3_8[9],stage3_7[13]}
   );
   gpc1343_5 gpc550 (
      {stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[1]},
      {stage3_11[1],stage3_10[4],stage3_9[5],stage3_8[10],stage3_7[14]}
   );
   gpc615_5 gpc551 (
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_8[26]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[2],stage3_10[5],stage3_9[6],stage3_8[11],stage3_7[15]}
   );
   gpc615_5 gpc552 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[27]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[3],stage3_10[6],stage3_9[7],stage3_8[12],stage3_7[16]}
   );
   gpc615_5 gpc553 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[28]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[4],stage3_10[7],stage3_9[8],stage3_8[13],stage3_7[17]}
   );
   gpc615_5 gpc554 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[29]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[5],stage3_10[8],stage3_9[9],stage3_8[14],stage3_7[18]}
   );
   gpc606_5 gpc555 (
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6], stage2_10[7]},
      {stage3_12[0],stage3_11[6],stage3_10[9],stage3_9[10],stage3_8[15]}
   );
   gpc606_5 gpc556 (
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13]},
      {stage3_12[1],stage3_11[7],stage3_10[10],stage3_9[11],stage3_8[16]}
   );
   gpc606_5 gpc557 (
      {stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[8],stage3_10[11]}
   );
   gpc615_5 gpc558 (
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24]},
      {stage2_11[0]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[9],stage3_10[12]}
   );
   gpc615_5 gpc559 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[1]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[10],stage3_10[13]}
   );
   gpc615_5 gpc560 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[11]}
   );
   gpc615_5 gpc561 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[12]}
   );
   gpc615_5 gpc562 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[20]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[5],stage3_12[7],stage3_11[13]}
   );
   gpc615_5 gpc563 (
      {stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage2_12[21]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[6],stage3_12[8],stage3_11[14]}
   );
   gpc606_5 gpc564 (
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[7],stage3_13[7],stage3_12[9]}
   );
   gpc1_1 gpc565 (
      {stage2_0[9]},
      {stage3_0[2]}
   );
   gpc1_1 gpc566 (
      {stage2_0[10]},
      {stage3_0[3]}
   );
   gpc1_1 gpc567 (
      {stage2_0[11]},
      {stage3_0[4]}
   );
   gpc1_1 gpc568 (
      {stage2_0[12]},
      {stage3_0[5]}
   );
   gpc1_1 gpc569 (
      {stage2_0[13]},
      {stage3_0[6]}
   );
   gpc1_1 gpc570 (
      {stage2_0[14]},
      {stage3_0[7]}
   );
   gpc1_1 gpc571 (
      {stage2_0[15]},
      {stage3_0[8]}
   );
   gpc1_1 gpc572 (
      {stage2_0[16]},
      {stage3_0[9]}
   );
   gpc1_1 gpc573 (
      {stage2_0[17]},
      {stage3_0[10]}
   );
   gpc1_1 gpc574 (
      {stage2_0[18]},
      {stage3_0[11]}
   );
   gpc1_1 gpc575 (
      {stage2_1[12]},
      {stage3_1[3]}
   );
   gpc1_1 gpc576 (
      {stage2_1[13]},
      {stage3_1[4]}
   );
   gpc1_1 gpc577 (
      {stage2_1[14]},
      {stage3_1[5]}
   );
   gpc1_1 gpc578 (
      {stage2_1[15]},
      {stage3_1[6]}
   );
   gpc1_1 gpc579 (
      {stage2_1[16]},
      {stage3_1[7]}
   );
   gpc1_1 gpc580 (
      {stage2_1[17]},
      {stage3_1[8]}
   );
   gpc1_1 gpc581 (
      {stage2_1[18]},
      {stage3_1[9]}
   );
   gpc1_1 gpc582 (
      {stage2_1[19]},
      {stage3_1[10]}
   );
   gpc1_1 gpc583 (
      {stage2_1[20]},
      {stage3_1[11]}
   );
   gpc1_1 gpc584 (
      {stage2_1[21]},
      {stage3_1[12]}
   );
   gpc1_1 gpc585 (
      {stage2_1[22]},
      {stage3_1[13]}
   );
   gpc1_1 gpc586 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc587 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc588 (
      {stage2_2[14]},
      {stage3_2[6]}
   );
   gpc1_1 gpc589 (
      {stage2_2[15]},
      {stage3_2[7]}
   );
   gpc1_1 gpc590 (
      {stage2_2[16]},
      {stage3_2[8]}
   );
   gpc1_1 gpc591 (
      {stage2_2[17]},
      {stage3_2[9]}
   );
   gpc1_1 gpc592 (
      {stage2_2[18]},
      {stage3_2[10]}
   );
   gpc1_1 gpc593 (
      {stage2_2[19]},
      {stage3_2[11]}
   );
   gpc1_1 gpc594 (
      {stage2_2[20]},
      {stage3_2[12]}
   );
   gpc1_1 gpc595 (
      {stage2_2[21]},
      {stage3_2[13]}
   );
   gpc1_1 gpc596 (
      {stage2_2[22]},
      {stage3_2[14]}
   );
   gpc1_1 gpc597 (
      {stage2_2[23]},
      {stage3_2[15]}
   );
   gpc1_1 gpc598 (
      {stage2_2[24]},
      {stage3_2[16]}
   );
   gpc1_1 gpc599 (
      {stage2_2[25]},
      {stage3_2[17]}
   );
   gpc1_1 gpc600 (
      {stage2_2[26]},
      {stage3_2[18]}
   );
   gpc1_1 gpc601 (
      {stage2_3[26]},
      {stage3_3[8]}
   );
   gpc1_1 gpc602 (
      {stage2_3[27]},
      {stage3_3[9]}
   );
   gpc1_1 gpc603 (
      {stage2_3[28]},
      {stage3_3[10]}
   );
   gpc1_1 gpc604 (
      {stage2_3[29]},
      {stage3_3[11]}
   );
   gpc1_1 gpc605 (
      {stage2_3[30]},
      {stage3_3[12]}
   );
   gpc1_1 gpc606 (
      {stage2_3[31]},
      {stage3_3[13]}
   );
   gpc1_1 gpc607 (
      {stage2_3[32]},
      {stage3_3[14]}
   );
   gpc1_1 gpc608 (
      {stage2_4[39]},
      {stage3_4[13]}
   );
   gpc1_1 gpc609 (
      {stage2_4[40]},
      {stage3_4[14]}
   );
   gpc1_1 gpc610 (
      {stage2_4[41]},
      {stage3_4[15]}
   );
   gpc1_1 gpc611 (
      {stage2_4[42]},
      {stage3_4[16]}
   );
   gpc1_1 gpc612 (
      {stage2_4[43]},
      {stage3_4[17]}
   );
   gpc1_1 gpc613 (
      {stage2_4[44]},
      {stage3_4[18]}
   );
   gpc1_1 gpc614 (
      {stage2_5[32]},
      {stage3_5[12]}
   );
   gpc1_1 gpc615 (
      {stage2_5[33]},
      {stage3_5[13]}
   );
   gpc1_1 gpc616 (
      {stage2_5[34]},
      {stage3_5[14]}
   );
   gpc1_1 gpc617 (
      {stage2_5[35]},
      {stage3_5[15]}
   );
   gpc1_1 gpc618 (
      {stage2_5[36]},
      {stage3_5[16]}
   );
   gpc1_1 gpc619 (
      {stage2_5[37]},
      {stage3_5[17]}
   );
   gpc1_1 gpc620 (
      {stage2_6[46]},
      {stage3_6[14]}
   );
   gpc1_1 gpc621 (
      {stage2_6[47]},
      {stage3_6[15]}
   );
   gpc1_1 gpc622 (
      {stage2_6[48]},
      {stage3_6[16]}
   );
   gpc1_1 gpc623 (
      {stage2_6[49]},
      {stage3_6[17]}
   );
   gpc1_1 gpc624 (
      {stage2_11[22]},
      {stage3_11[15]}
   );
   gpc1_1 gpc625 (
      {stage2_11[23]},
      {stage3_11[16]}
   );
   gpc1_1 gpc626 (
      {stage2_11[24]},
      {stage3_11[17]}
   );
   gpc1_1 gpc627 (
      {stage2_13[24]},
      {stage3_13[8]}
   );
   gpc1_1 gpc628 (
      {stage2_13[25]},
      {stage3_13[9]}
   );
   gpc1_1 gpc629 (
      {stage2_13[26]},
      {stage3_13[10]}
   );
   gpc1_1 gpc630 (
      {stage2_13[27]},
      {stage3_13[11]}
   );
   gpc1_1 gpc631 (
      {stage2_13[28]},
      {stage3_13[12]}
   );
   gpc1_1 gpc632 (
      {stage2_14[6]},
      {stage3_14[8]}
   );
   gpc1_1 gpc633 (
      {stage2_14[7]},
      {stage3_14[9]}
   );
   gpc1_1 gpc634 (
      {stage2_14[8]},
      {stage3_14[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[0]},
      {stage3_15[5]}
   );
   gpc1_1 gpc636 (
      {stage2_15[1]},
      {stage3_15[6]}
   );
   gpc1_1 gpc637 (
      {stage2_15[2]},
      {stage3_15[7]}
   );
   gpc606_5 gpc638 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc639 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc640 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc641 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc642 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[3],stage4_4[4]}
   );
   gpc606_5 gpc643 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[4],stage4_4[5]}
   );
   gpc606_5 gpc644 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[3],stage4_6[3],stage4_5[5]}
   );
   gpc606_5 gpc645 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[4],stage4_6[4],stage4_5[6]}
   );
   gpc606_5 gpc646 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[5],stage4_6[5],stage4_5[7]}
   );
   gpc2135_5 gpc647 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[3],stage4_8[6]}
   );
   gpc2135_5 gpc648 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage3_11[2], stage3_11[3]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[4],stage4_8[7]}
   );
   gpc606_5 gpc649 (
      {stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[5],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[4], stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage4_13[0],stage4_12[3],stage4_11[3],stage4_10[3],stage4_9[6]}
   );
   gpc1325_5 gpc651 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[10], stage3_11[11]},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc606_5 gpc652 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6]},
      {stage4_15[0],stage4_14[1],stage4_13[2],stage4_12[5],stage4_11[5]}
   );
   gpc615_5 gpc653 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[7]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[3],stage4_12[6]}
   );
   gpc606_5 gpc654 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], 1'b0},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[4]}
   );
   gpc1_1 gpc655 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc656 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc657 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc658 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc659 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc660 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc661 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc662 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc663 (
      {stage3_2[6]},
      {stage4_2[3]}
   );
   gpc1_1 gpc664 (
      {stage3_2[7]},
      {stage4_2[4]}
   );
   gpc1_1 gpc665 (
      {stage3_2[8]},
      {stage4_2[5]}
   );
   gpc1_1 gpc666 (
      {stage3_2[9]},
      {stage4_2[6]}
   );
   gpc1_1 gpc667 (
      {stage3_2[10]},
      {stage4_2[7]}
   );
   gpc1_1 gpc668 (
      {stage3_2[11]},
      {stage4_2[8]}
   );
   gpc1_1 gpc669 (
      {stage3_2[12]},
      {stage4_2[9]}
   );
   gpc1_1 gpc670 (
      {stage3_2[13]},
      {stage4_2[10]}
   );
   gpc1_1 gpc671 (
      {stage3_2[14]},
      {stage4_2[11]}
   );
   gpc1_1 gpc672 (
      {stage3_2[15]},
      {stage4_2[12]}
   );
   gpc1_1 gpc673 (
      {stage3_2[16]},
      {stage4_2[13]}
   );
   gpc1_1 gpc674 (
      {stage3_2[17]},
      {stage4_2[14]}
   );
   gpc1_1 gpc675 (
      {stage3_2[18]},
      {stage4_2[15]}
   );
   gpc1_1 gpc676 (
      {stage3_3[12]},
      {stage4_3[3]}
   );
   gpc1_1 gpc677 (
      {stage3_3[13]},
      {stage4_3[4]}
   );
   gpc1_1 gpc678 (
      {stage3_3[14]},
      {stage4_3[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_7[18]},
      {stage4_7[6]}
   );
   gpc1_1 gpc681 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc682 (
      {stage3_10[13]},
      {stage4_10[5]}
   );
   gpc1_1 gpc683 (
      {stage3_12[8]},
      {stage4_12[7]}
   );
   gpc1_1 gpc684 (
      {stage3_12[9]},
      {stage4_12[8]}
   );
   gpc1_1 gpc685 (
      {stage3_14[6]},
      {stage4_14[4]}
   );
   gpc1_1 gpc686 (
      {stage3_14[7]},
      {stage4_14[5]}
   );
   gpc1_1 gpc687 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc688 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc689 (
      {stage3_14[10]},
      {stage4_14[8]}
   );
   gpc1_1 gpc690 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc691 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc1_1 gpc692 (
      {stage3_16[0]},
      {stage4_16[2]}
   );
   gpc606_5 gpc693 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1325_5 gpc694 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6], stage4_2[7]},
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc695 (
      {stage4_2[8], stage4_2[9], stage4_2[10], stage4_2[11], stage4_2[12], stage4_2[13]},
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc615_5 gpc696 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2]}
   );
   gpc615_5 gpc697 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[2]}
   );
   gpc606_5 gpc698 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[2]}
   );
   gpc1406_5 gpc699 (
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2]}
   );
   gpc2135_5 gpc700 (
      {stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1]},
      {stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2]}
   );
   gpc1406_5 gpc701 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5], stage4_14[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], 1'b0},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[2]}
   );
   gpc1_1 gpc702 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc703 (
      {stage4_2[14]},
      {stage5_2[3]}
   );
   gpc1_1 gpc704 (
      {stage4_2[15]},
      {stage5_2[4]}
   );
   gpc1_1 gpc705 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc706 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc707 (
      {stage4_3[5]},
      {stage5_3[5]}
   );
   gpc1_1 gpc708 (
      {stage4_5[5]},
      {stage5_5[3]}
   );
   gpc1_1 gpc709 (
      {stage4_5[6]},
      {stage5_5[4]}
   );
   gpc1_1 gpc710 (
      {stage4_5[7]},
      {stage5_5[5]}
   );
   gpc1_1 gpc711 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc712 (
      {stage4_8[7]},
      {stage5_8[3]}
   );
   gpc1_1 gpc713 (
      {stage4_8[8]},
      {stage5_8[4]}
   );
   gpc1_1 gpc714 (
      {stage4_8[9]},
      {stage5_8[5]}
   );
   gpc1_1 gpc715 (
      {stage4_9[6]},
      {stage5_9[3]}
   );
   gpc1_1 gpc716 (
      {stage4_13[4]},
      {stage5_13[3]}
   );
   gpc1_1 gpc717 (
      {stage4_14[7]},
      {stage5_14[3]}
   );
   gpc1_1 gpc718 (
      {stage4_14[8]},
      {stage5_14[4]}
   );
   gpc1_1 gpc719 (
      {stage4_15[2]},
      {stage5_15[2]}
   );
   gpc1_1 gpc720 (
      {stage4_15[3]},
      {stage5_15[3]}
   );
   gpc1_1 gpc721 (
      {stage4_15[4]},
      {stage5_15[4]}
   );
   gpc215_4 gpc722 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc615_5 gpc723 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc623_5 gpc724 (
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc2135_5 gpc725 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1]},
      {stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1]}
   );
   gpc615_5 gpc726 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], 1'b0},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], 1'b0},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1]}
   );
   gpc1325_5 gpc727 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], 1'b0},
      {1'b0, 1'b0},
      {stage5_16[0], stage5_16[1], 1'b0},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc1_1 gpc728 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc729 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc730 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc731 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc732 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc733 (
      {stage5_12[2]},
      {stage6_12[1]}
   );
   gpc1_1 gpc734 (
      {stage5_18[0]},
      {stage6_18[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA162_12 compressor_CLA162_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9477c4664fd25c48b83b5f13e4d952919e38d2d194ff1169bd733e93a3449bfe663274a87b5d49110e453f0ea1491d9c9e69e2e5fba68e93184c19e36f28e1efbcdd50f5f5d885810f42f06b5fe2fe3b668721d8cd23b101809ee66b402bff11cc7d09f18468b88e27adc4e19de275a88eb2598556b1c1429ca16a0eb04472ccfc8db7a1f6edd5d61a33f87aa4a205162269ce8b9b760fb827f4c5f7facc224356ac0fe82b86a84457a32a48c0831e686a2dcc61d3d3aa5e22870a7d372c8054d6e425cb105f51f11258541c18c22bfb3dc3952e6c94336259fe6ffb3f5c6432bdb2f83a24119b00c1edd0c2216a0eb3f76712;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfb89cd6795fda8dc51a9e5f774ee1f3330b7a4ca36e95a936a7f03bdb5327f52e77b520b57b2712a19c5d184fb4d84faa884bd1b94417734fa891559152e8be3c73a62459cfe52aaf1fee651b9f41efb14c6e8b2dc01cccf43a6d101b741e3cc6ba5f6dd6c46bcf2ed95131b2aaa0bfe28334460c6f513edb70c4e4e688bf6f5ce212bbd743cff0a2a63b805a0cde509e5e47eba1c87bd04c88c55570bf975fd6bc85f29742f2b66ae9217e7fbcba3303fbaa8b071f0796efe6a972b3f8866667597d37e7ee94162b98d5f755f870bf3a54d53882e8049a74060f75ebe86492b3d2593e79e31b568818337cce397da5e51de88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h92a9d6620d4d2501e1f41f1335d814df6317e799caf0f3682ef6041de1c76530416407b3e852dee4fb15dbf4d5aca78e1193ff1885f967c0669203ea5e713d7395633e0b2737acab400a04d572a22ddaf5f32ddbbc93d58ad1cd9a3758f3d989e7362f66519bf51bb6ea4d61a80df58969df10254bec5e3f15dd194903d8eeca05ad17a283b83609e0c372a8195f07b8042a34ed18822450fc2a740ae801e144a5b943372ea871c0cd69e1dd2c583dc3c3db038856f4d6fb2db7fe81612fcb4295524e5e1d5b450d1f2051280362fd5da6bf81277781d5cf67070731d13e9a340c7f0bdee7233e5cb0db07c479d49612f5cf4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9d8631c306f163c57c06d8567765daf52d806c84bebbf44f93161fdd9ff928021f1293af1cafcf5f5e4639f86450ee84c79c307ea734fb14f35e9fe92e9236f25cf3423e7942955046ef0c0184c3888d4fd8de237cc7bbc044897981e3470757af08f20a7ec3d217add66be499cf01427c3c5d6b46e154c3382b2c43b42350acbe65b4726eda4b5f6095a31f027c0f688f1d285c5dc536de69874252753798c13306122f1a7b6160e6f45b509d4f112f1814a4275ca8da28aa24471b11f81fe55af185bf2b4208e3befdc224f81324991db5d030b8e1e01af8f3900e90c071f179a90f894a3721061c0a23a15805ab33a623ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd074e11545aea58cd8539a73a41135cd0b9c2d7eea96508cb0dc41cfd366893341f88553dad99426c644407acd8f88f29d306bf1dd7eabe5baad221eefc3fa62baed9fffb0834df3cda468b533819d8d224984ee9a6110cb0d20e953c38249efa1eaa4dcbdef6567d9c0cfd36b0388680d7ddbc08d401e33d8aac75e8a8532a9bf99e1125dfdda3c1dff24123ba9366f59e3fc954516445f779a795c8cc5d86e2f10cbc68b72fd966c9cdf5e598a0c4475c23b578d86329f57244cbb11873b7355ba7a0bb8418ad5fdb807092671bf5330a2e6c34d16128ffc8ced90d49c4cd6603dc6c4577f51d479714949e8ae815cea461a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc3c76d4643c0bf06b11201d9da5a2308440d35304895f3cb591f25ff5399fbcc95427e66ce5a90c0cbadb18835ef747cc39fbc817a5a8a7230452452d58de009e4a5b216b30956a6069c03ebe820a7dcb093c0dba345b3f5f3b312ca5da5c8fd66a9850cd6db5779ba8dcb5d96828616cc6cd5ca9b1895b4ca55820ac2b5d9e95206dd7a4b03b184b001c774815fa626d91a39f8f8d5e85ab45fb5364e0a77e3474f10b7abeeeac309c135c23a43cf070b082203fa5f10f0e77f1f6b5da7f97c89c34e07724bf7b40675233b0a994fedd32f2e689098fd42dadf5e4293a1ba5995182a2b0788554a0462bbca167c9875d5430b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he4ba8fe619e3536d4fac55e6dcaa4bd43f8a76af723ac865d5e7d0646ca23d1f42ffedfa06950323dfa4d0fb7f0dcd4ac6898ca8b2a2adef53f675b65606d369eeb92a805aad688232e2ed2b7a10b78b7ca3caa32891106f8c4ae13930488601f3f64666e4a325596cbdf62ab64efa4b0fc3a0a4ee27be23b099e3063fc2e7773c778986fc5941281f66b840ebab37513b63d4db2fe41aecf260d04ce8102aecdf77cfdbeb481a5db91f0d3963e617a9afba7c79ccb546c54c3d9ae845a7efa03cf698644ae3ae3524a36167c8bd9c7dfdb2e302e5ea41188d14ea39ebe71202e57c0a77c3e5c559081b5bd81ea7366efea3e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h515cb625cce20928cb842109a44e522092114459c1909b17b45a07ea3b52608334537e143c4424d098bec94bbb8444a7a660d4ffabcb98b1775ded0eb3db61e9fdd09ad22aa7ff34fe300d1d9a111912487b2419493bb5c727c35dbef1f18f56b57603017fe25a48449106ed62d263ab7bc812836b11cc8b28f515f5e1ce9197186afbf590a2848b71f20b4e031ec39f806f45f26b477c268b50cfcc9e55eaf777d9e3d5056dbe9b298366670b21b7b43108982b64f3eab668fe9560cf4fbd4a6c8a794b2d797fe532d12e8fe83eafc9948d9b4b603c09e78a99c09b0aaa398581d19c00d3043cbc0b230099639bd1f95b2d36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7b3c1a3641cc707abdbf8124d5c40bb8d5ea78c6d1e0ec0fcc41e30769f0e2a95238fcd7f475c5c228364d904f3f0d61b5d0a45d3886e6398090103971a88a30678a552b705517ad272b94d22f511e9d50c641546d2f2dcc0451156ab70c5ee6bd0354d58ba68ebdee82a480153ebebc481688854fa2f033b2239719ede38c2de2a14a97e8c22fcaf6a14e1cafdb69094d2a593f7bb5fcea36753dc7dd3a56e50b939835175c6903e10445c8ec35261dbf066959972f13463ffe6d580b65c35418eece4123f34deace5684ccc02a5befdbb625d3e5b9531fe2bea78310d00ae0437e8798a98f2d7c22d2e6805b1707ff891881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he93e872f2c723c0832491fc2e4595390f98a6758b858f0f13fe3d5d196aff8ca26936ae47ba9d8cada191abca3e931689913aa83827ab8fbb27de179a50dc5fed04a1b9f4d75ab80533616b81a334b9dd78c0b0b2048fdbde131e582552423cf15599b18f104ad0626df66bc789ac5a0a3f02eee51ad890ae4354afb6c5a4353329162324f0618638c5694290071940e168f0da43e7c110909c7ef92cd19c53b298c0462b54178ff7d25b45f7a8577b8b334b1f335a37b7dda8337281bd739cdcad9b42a4876fb27d2a232aced5ee503ce6b0322609260ac248074acf96f929669c9bf60e5a5937780f16bbfbd68180b409254;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb8e1334849d682fd0571605f75097355877cfed4e081dcd45a89b1aedf5a0fb1644772c1a62b04bcd6961de018c50c1fd2c23d0db0eb535666e372d10861100d94d3f63a4e73dcf50744a0e82cf62bf64fa802032cc11e315267d0b2129a01f0de31c55ae57e8ab5e618fc212a0e64b050362c1ea0c2c3aed5c519405cfb3da9b31112a7f7bf74bc202cb5e05b3715abe237df4c80688989848965e8f40bbcb2a66c33992d0fb930402ac9c8918e542aada2329e3189fd65f5d86305c09bd2050a351dd13e436526a06137260c13930c4a68032e43af7ee15e5c481f1a9e91055786feb4adc5f5e459394d6bac34ed0ea26f3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9b0aacbc2b36a0bb09f3b1d65cb1d5d011bc08adac9d446475a829f2bc7d221ee5af0199780e0582ccb2fd1970e4116ff74d036bc4c84f75d0d888eb225e1e7773adc40dc3989fdbfd6cfc32395999b28c7651c5c9979e1c0e1c573da5cdbda63a6731eef52f9b92edce8fb65638d0d1ce53ea6948b6e52c80cdd1818d9f9efc24af9b1fe54f0c5180d10f5abb22d347fed42eed9161c22724497a68534f6da9117bdee8659afad45daa8927b761e580f1a4e41bfdea64d8dda2647f599a9a469f64f64318e8dbab0a311fe16905c3af76fe7ea3264d7dd64d667b0165120a4f48e1cefb3e82308d600035766fa3adfd071a8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4c3cb37d0a01da39682c9c50f9a4ee51715cea79f43fa1444ad4679ee611978502ef1c2c0c89310a22e287a71e4afe756ea75e59691b486491cf56d33a88c32341d00ae84737270f6421fc2ad89236239d6a84618c8cf652b9ce772c26f97ef1eea1aa075dd605d9c083413f3fa9353d8348e95340c877f84a39b6a61c0cbf82fd3eed58de6cc386c5230ec6fc2202f568a7155f4d1734b0a9226187cd2bf8666618e61c7276f1c1f6ec166fc57d6a12dfd85fa577832d9deb57e10ed21fd22a7a2f81f0efe03a7964fef836600ed63afe2236f6bc47f23e4fc5475f07b75afa5b0d6087522c93420ebbae0d9c669db1401ee7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha3c25b5e0a17638a1da7bac08b8f68fbc011907010e7179318ac64168f3a79eb88799eacdde7d88a31803fae88902185a50bc53118f80e5058d6efcb5459eb9e764d0b7683f4c89dbb42bde2454fe735bc98b2b69eabb51c6940173df250fb95ff7dbaa2131a5a6a02035f698822774f995bdd685bf1966e25fea90725f33f25ce2059d9353b88f1917a163bc4eae040a9868c9663df9ad6acac27c3305da2805ef0e1a07f02b73c242069775184241aee5c36ff4dd8426240cd49af7a4eafefe335386cf87de2f74c2e9ad2aa7a4ecec6a071389beb9ca8cfcb4fa0f8df33ca2e6e1f8c750626803e502e81f082ddc29f61e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd7b0f1b8e2167bab8096dc9bb44f9379a08a8a61a1b26cd685cdcaefbd8164c0b122bcf3a7505e30c44949fac121fd0056224b286192aceda0d511f4534344fce012b5f2b18c70f9368e20048605dedca71e77f6fd7cc25e3b550b623e5c73de96572758aaa8f72158311d310f9fbdfb7aa72211c8af24bfa266ad88d4f65dd443a55233c9d426fac889baa0f4f064e79d2d1dedbb170745507e2222c7414ad084818c8ff3769f3339eb098ebc061dca5c63f417084c323c9354cbd26fdecee8aadc266b370cd0d62eec48a7531e97affa8701f249b9762271852741d1af63d76d804db37759066ea618c1c8a41cb0a0da61d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd3294e61cfc40c0ae76cc9aee967b1d58fb31a8341680566b8bf8b985f996bff6d9b7eec9e34cda62e0bebcf9bf91723aeed3c0320d6ed2949d25e75910b3702cfa71a896089f83f98194b2ac27193da4e0c5c1441308b85bf92964581ff86f6456d44ca1dda6d55fc1aab32638b850972953cdfd67de5a7b249f9a231b7320091c94103b6c152d6695fad520ae0fb0ffca7b43d116bb392856ddc95b7fed11c43fca266d2698fa14e91db128a17660a375984c294db529cf8328569949607a2a02bdcc4e680e38802b6d2c284ddcc6b872d967462e25bee0631c2c6b3c9f5522958b0952f0ce85b0a2ec943ccf79cb406959c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he270d3d098fa70fb032fa1f8e4acd11a3678110568180d4e0c19f8c4414b8b18870a0933190242772aa956ea73a52c866310d5c9193fe2bf52ed783547e969cf75d048babef14aac03cf8c54d7876b6df41a9189dcf02aed020489a868290e49d631c81081aa9625ab917de1f00fc65618d15ddbe6ffed812d8d47c91c584960134022161d84e28b47e7d3af459e84a2a2bc4d5761b64f0b1d85aa0a95bd6e8d0e25c9dec3e96245641c1c413209e092fad7566f15edd6f5ff9ed29c783afb7f7c5948193d227fc01ea99ad2471aa58229cef687ae27fef6e29a9ca6839b11301c4dcdaa6866d4f8b2c2d0805bd5d448c3d244;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hecb88a48e74a67bdc439d030ea5c25963ac121ba373d6ef64cfabe0b16e2d6cf25184fe28caa748f1491123003edbab92371078055831cd5cfd6a1b17900c01880ecc1b876e1157b77b7486c8d5696cce47245b0872c4ddfbd78930c01cbc8c6acd5923566baf63e5feb7f17c8bb888c2a369961a659c95f4738971554befaf3b42118b9f52411b1a01fd5fa0128165a808a9f324d7fe2024935e3bde029ace6cf8a00aef73451849ae85d52abcd6d8bc161a6cb455b4de09bbfbc245c152dff785c97df23bdbdfe984ebc10ced2ba74dbe4bb7e774f73cd18358373180c8c90fe9e813ce2dd183f0b7406a426f309d9816393;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h6a0d2bd24d66e6da6c5998f07e3aaee1649e2306b498c41b8a32f6451b265035cd4e90fe38b91cf4fe8f8b08685a2bc1fe55af5a01f0e17f80525d8e471824347b4abebc84c36a8549d19d7cd4eebaf04473af5332ddb301eccdbe72811a6105806fc9012cd5074572c991ccd328697f49cd19e002a0f8fa293db5cd5e91c34f98e190fbbc748bde7434170bc1d9c45d71916696562af68f7b7fe79ecc0fba4d4d1e7e6b46a190663f0e0ba1d2ed558456571441daaff281de4aa09cade0281cbf057f827986ed44a7c13cf1e76a365ddac000df6ff323b4ae2c3c3538f53309634904f9395e41c3f13a20b32a354987a9e85e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h60276e7237dce438b738cf1350e1a1420c01f24b850f182be935ac0a8423904f7b82fbff5ff64f9a344f4f0f74036e4c4d8b5a872ecfd70386bc8d9c9ead00b38ab1d38a66ff5ac27495d6a4d47c3820a6f60238a32a8ec5be8812d5421af810029fb640dd8d8dd38fdf050468defeedee4422e75acd698f934337db31e9de7befe3a792fe31d35900b43a6bd2e55fe1ff10dc4f4e68261c32e6fcddf5ad7bd50a5aecb47fe15b33c1abfdb438c40c9c17880d41d8e94891259049d7044e3c1dfbd57c98cc0e6d41a483f6d9e5675a342f2da3effb6e24436182bacfc047603c03efc9404b425283cad4b0f6deaea34cd274fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3a7282fb6aa72167cee9c3264eb7f69c65197730199b45e44d020030359e679e6bf6d7f308e30e6c2c5117942ca9a1cafab12c97bf75bb5332be35df174fe416a8ad1b6157e4909320bb982866791c66960e44ea705a954530465d3b81697abec4dc6401da64bc54f96953bbb4c0877b00c60327110b2ba11b6c1c8d270541de3e62c89c2d05ad61f129ed2d6cb722506fe0d2b046add9f9e979ae8b9075584146a207a28811c42e80d722d14075e8b5ed47fa8ce94464e40c4c770320601f44f4a30bac0cba4675d628a671003e963c5a47f20d41e96e4c53f25dcbb831c51602e03d6ece1cf435077dc8199931a2b9cb6223;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h83ae09003a97b12faaf547f2cd16e062ab531dbbd0af002c77595b20bdadbf2f8392164baef34187c86fa375f7419b922e8eb9625b6e3d75ac996297a314587e18df2ec69938e7817e3e355e1b8ea26c2a2f514da724c13d0e5f290f138b8c5215b17c3bcfae90b9de3a3608ae510487407b8d3a27f9c6555ecf11537ed08dc60a76aba44bd2026453cd166b07bd4b3e065cfe1e9b73c6471771bf935fb0b9d309c37981c98223e47656c3c365ed6f8b55a4ebae887491fdfa5d9736407ef0d11c50e0d83efcef6d4edf2e92d784dca0b5f4dfee00df63499a153bc15c53c9ae36e72bd6c1500ae5eb281e5969604a0cb6c8c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4b5fb840c9755749ddf5b32c000df2b2574ec0acc23da9f74c10872120788da842662403447778bb2c099aef4ffcf7a53a457197ba5d2cb671659c444099bab60b086c6925f25df59d15019576b8fabdcf74dae53e82e3b526dcae44636e7b15c3bba62302f084e56328b924366d0e906fcb9f9b2390a2376f72777b0a44b2412a86ebafb15aa3235d7280b0a77a05525ad3c59c0ad45871d83235b1299f6d19db76c13a1ae5d5799d08d7b26fecc9fcec8997fc448c8edac6a7dfbdc58d3ea49f08f594b5950765cabdfdad960c71802585c9a7e555e9addc2ec5f704b439e9bf8e45187cdbf5436cc558dafc09727a59c2da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha56074acb2cfd297d83616644109869a55c9200a83fe9b0d309acd65bd54c1be376ecb076e860dd569feff97c06168c68904f2324502405a068083e0ebb0673ce7bfaee8780734579f112366bcdda6bd0ba790f20bfc9085a600567a50134efd264480b70491adbf7e187e56671eba0fb9c453424e8b9fe98936fd3f03fcd899f71c1fb00d63f4d56ad055c533c3d554c901a3ebaaa5c70906b9b4ed424f2a1e21a3898587f07326c3f3c55476a062252f7905ff3e7a2f06199b67f543752d3078bba7c66868659fd4fd054d0fcd263c56da9f137ca49257761e6f253bcfa2508a0d452c39a211e20878db1c2adeb70d4ba0a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf2a76ddd2c3a03734a5d2693584d492fbf6cd8fdd7b3b15f6e5f1a1e44bf931153b8eb9d006cf2ccbca5bd856942ff9510aac86056b8d9a305d0e5c6972284d4ce99034b6f220f595b5de8fa191be0577666463962ea8d7e7857a0f147d5a6e28df2740776688b214345e19dd0ec8ef2f07df9c179a8a6c330af708a384b2215a027facfae673d41f0c63b9b503e1049e48b4368d62065c9aac27d1b7c096cfe49b922490af5d225e07fb38de33a70d5527b96c123fa7ae0b13a8b8d7d92bbdd9017259fd949edbb23c8f75b103c7af8c55f15b249227f144a56b6d112c83efb5b33e3455fdb9a14beaf67eafca42575f49b48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h95261a99f3eec84bd697c342eec618f52566d51fa62703750874d6b7b93cbf134a716734e52ee8fcad6b4042c98c6a3451304dafe8e01ea0fe2852efbad56c0498c25aa3cc83591b1d72b824b76182b4a3fe0545dfa727a4e634aff4e62d3999630dd833361b60b9cda93ead2a3d780a350152106efd4e8c5f50690af89a8ad5c63130cc76ce416135dd1887470167b3003dda1963d92b8468e686bbeddd8e3e09d4f685ff92a7608bd9e8aa0dde7a2b4ead88cd2007b51ddcb3cfa192ac1aa316e3f2db3e738e5aa2461e395581a539717e5a68b3e1f2a86fe48138054032c14f83388463c7de7c79a4ae1e3375534685809d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7862ec6fad7b523fcfc681590b2c70473fbc84047bfa2dcd2706e66114fcb7c57330b4946c1d8dc272c4ae3dae55da78d8f10f83f05b5517cf6158c601c831cde91b7104e174e3f9983f20f0473cfcd1decead8758261bad7b28d5a7dbb234d0dfd104b83b3991e3adf2ccf790fda9b44f303489b02552f3cec7fcedf17b611b3900e3a68c47629547cc03222269456894ab19504da0e06709e508842f85731c40da8aff05dbe5a5fd31fcf3909b8eae6666658e0f4d488b1c6406cfc074dda8fae9358850786d0f9d28bb818ba36ffda7624ab0b4f7ff48248119bb4cd020646b378ff794808354a6d5babbb6cd3fbda27bd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf0945463c3678ccf81a37f48bb9e922d68967855d7361f854be6e9ba0e519a548881adb82a7dc241a679d71fb3f132a579084a8eeb43a5db07b569baf2f2fdd209a9381b258d750c9c191e92d23529a72e4a333c38536efb6319a7f6a279241fd018abc04f8bce3d67e8869d51a477b0011d6d8e3cfcb06ee23b88ca4850e8d7c8eb6492781735d911361364135a2e706435682fc6b2a499991a3768cebf1c699d3b710ef10c00912c346a4841b6e80b15e7114cfb7c634995b3cf6b926c73facb66d6794bbbd383183985371e1e3b47808e796b53ab4c51249bc28cc238237f40e568f260ef2f729f181e437e436b9d34ce16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd50f7d567cd175d23030c54f947eb47482fa899bdcdbce12a0d6359d7f5e2bf12cdae2ce7d05c928e57a8fcbb3714d63ef3fecf47c4a6bee5c96a746a763cee101375ee1f7da9e316c89441c927030e09ffb96298adef4f9c2a021f79b049fe6b77801c41c21ba239c31b484ce947b07712c83b872ddd472dbd88d2843e78c43734d2f9f924778672aef5e054f8bee78ad50a6f39d45e7cd84a34040c00ef98f88a263b31807a349c3edde41b7a0c537348c1d1a3a815a4ab7e9f0f19e31517b9ab196f8c5a0c66da297c493604c46767287b02ca7c8ee926e2221d7dd3d3c5d27151f5063f9075e5008de784fd995eb450080;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbb0c72dae0b5ddaafc39d09ec3ecbe5fb0cb176908db11091370fb9297d61fdee347d5d096747bce1ee0e74618ea23bdf60b0e56ec531943e9694078c1014ec1572a32425d10b1b5a5d9f6542d4de3079cbda21ed5898608968f88fca6c48221d9aed7c8998639cf3579a6273d39b3811cfb28069949d0f087bb635f10ba9343718d12a2e07f275174afa3122c1e57fba7aba93a1efc3e34860e26ff19bb68d1179f947ac899a995cf5ac899c2d638bc6876c5fc16d8af4ab03c020e9f423c9ad7b7a224328ccc618c2b58e494a178f4a757f664738a0b65489981f2419cdb0641767733ae9828f0906280a1ef1d23c90bb3ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7faf328546fc9557ebea9ade8e98fad9a7c1acb57b46260d1aa08588ab4ae64a442c75b4570f601695906870e9a7f1bfad50b92a45eb5d2ef276ef1374c0806af39747b489a0ad5f8b4574bfa3b88dad5d80b6b773d94234968fcd38a2fff52a124d3d66fa1f51d1ffc577e6e97359202c535ac7e53351f4f5d3e2c01a0c85bfe26cebb700caebdf441d9922c9c5d450f6345533b0fea75fc72c794ec02888dee3e13872489bc3f375b9bb3bfc185d6c95f9bd0770432e89cc3d0090b3d865d23922f645418ca8313411191403c90b8fe4bdde9e2a655ca298e76a160a760a74f319888df22b35bfff847d28143999ab6635a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5ad81ab76093bac3c7e09d050fc764811474ae3dbaf808cc6d9ff7594eaac07c19e6817d08d17c8e90c2a336cc39b37ae260893608926b17a0349aa6e7c665bd96dcc781e33f6c8abbe0d1d98f176c5947f6f1aa98b4fea35e545fb1d712c74b5fa65dadd25dd7e84dfeb712bab23da2737ed598e4476643feb061a6b2777b097c1a1f47ad7dd09b79794750c9e8f638add16a16b7697a50fef4bd24e8e85da83059c89abf968a44d52ef3596afd44f1cdceec2ca9b4d4c87dd6c6f1e83ea61f79cdfdea2839de6ca35ae8ae6d43e9f44ebcd5a3e53909050f2d5c73ec9631d62c8fb2349ed16acac43a766268a5da0ecb17fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7d0dc37105b73385f670b6ea45b8fde4f96b3ee6831bb44a098ad818baa69d6c1cc1776da378ecbd340c421e1afb841445cfa99cd25269f5b98eb8db0f1fd3493d791d55444aad70bb44a461f198033165516931fa5b9241db1aa8d77d83829f5e5ceb7d82ef61f4e4d17056645f50d45a75cfad31d89f74e5f7c0fef9cc5a6d16adf46045a6ca7060db41ec1e68d44b1a4196350bb3442a908bb57e875b184cb6fb996f2451f86b0a7f946e6d7899c7dfa96e8da31cb00765d3516d91d2a5ac2cb884dc1d823fc4fed5a310782226358afc07ddb1b74ad1bf7f0759f307f3e831fce1928d3383531698be18a21b958ab3ced6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf6faf38d25e02aa03147fcacba8baf23f46a00a97008543ef0d6bb65c1e9b78bd7404aaf81d46f8168da4a7ac43b5dd58407f6226fa7b0f6149c1321e68186fcb2293d06d6361515f6ffc47471ed674e543b3babc8303ece784274e5ecdf1f21957e6077c10096d706c7fdfb5e5737b102d603f45fa0af793e19bc5854e1d6c3965926c2585e91bd79f3fde5abd87f91b71a05fb26da0d37986f96ab363717734d7597327c3bcaf791dbfcd051421d91dfd872c6c03bb189ae53b1dc4938c3b9bd69b10d72e36cd16d2954f1c3b9bb8c74ceb426e2cd2a07edc4f07fe94ac64d6668de46f3df2c5d4a192115b1b3872ad2e58a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf7c90aab9c4fe5d535e794e86dfe57e5b774480796999d7402ff221458e28f6268b504559269d9c6fc33f37ebfe8b3b84df1eab59a6f636671682889aec60d47f0c1283db0ffff559a1ec07791fdb68c7eca96ada9442241ca1f5ed2187ed9301af50fb2f83b360dbe4314906ffc0599b39444129e26e99755635cd814ee14ce14716f73aefdd6712aad0a0eaca0d8beb9a2d1e9fbc18a4f7c003ab91b7d2c8a257035b26877365bdc395f767ff46fd0a3d842cd6f00d9c2e3632f6d3c9e26f74e5c364af5c78f11378ae5f565c42b6baa15b45e63665d26634d457da424e8cb9e75f9c8b49940cf5ec2295fa84e3c986872ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd87dd684a0b85a0db74d691c14742eb6f315815c4ba1388a4945f5860c401208bc3be65e58cfb719befb5abd12dd7d2579c34bbee2a62dd18c6da567e592292ad7f9681801777123447e1227f929787da511773ccf1312edb577f3a0967f8fda165f127a33f554aa51eb5093a6b32c1b6a3a9e740a4f26c871a80c9f13a3621f3afd361c189c16188eff4022b86eba88c04370c4c64ea3897076dfa3ad9981f40cbcb8f8978b7f15e74255830def231d98b7765167b484476a7e915887e607082b2de288a3aa69fbe97877fbdbac5a85ee28aa029a646559b6ecb8098294e3a29d88f6c19bcea04323d0c203e2a275e560eec8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1bd114059de9e1c90d6c2c8b7816f57bb4f95cf4f865b951fe2e01e5c89986df47ff55155231115cd821fd67f781dcb548572664fc8e86bd5a763a9ba0ba4f714101cf06eb83a101f4e08ad7358a08223efc394ccfe3bb9c0d2297102d12908505bd0ada48b56ad9a82154665da16b65e36606624672baba614df252fdb634cc5f33f482eb90139aec6fd6cdb3a3ede993552bd4b109af04e30eb7a554024c66b4efaf867947fee122f79e9bc90ab45a4a3e1a7f0bd12e674a2ed709278497c2a94c2220598a359e0299b9a9627b50dba432d654e376184070159268e48d21750cf87c22130ee76b0526a87b3619c30333e7ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9830a3c5c31f9e1a7e28a5cd754f8228720544f53cce70a35652117baca77d7cecf22bc0bf137a892898bf99b8fe7df3af0ee7d72d47b6989f83f7b45567fae21da8312f45a4cea5454e4bb211d3e808e4b2983f1dd16ba8a4dc803d873a7b4481e69ac16424a8b2358ec1460b09151731991f01853d781dc215a1eb5769186f08601b327b66679f038519ad605ebd536b9d0ddad702a5d7716e911495772f252b1829ff88d4305a4dcf9cf2118143ddceb6b7948ef7d7eb9aab77f5ef9d74a4350773fd4199d85e8c21dfc912c658ee4321cd310cf9099533573a5be11ee2370218db50eb900af4cb2d66798ff28766b6ca58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he19e71c04ecc67d97695c3a90c6adf625c91b233e5210ffd4b23c05eef98d49b086fc8d6ea57ef26a2d2b1f47b83b954595243c45624fd65f2409e267b414c148604814d0e2f634b1506ea1f35b714d95a6edb2af0296738b72c247635e660c51d2bc87a5f1bb524dcd1f459f0e3bfcbc692bb0281df1ead27e07ea8215b2712bc90f7e17d114e5dd276f0ac027e607af7e1875a240aac8adf199c5c862fd6b09f632bd352f65772981379c8db1d31c37e8fd7c44b3318f57e880d6dd858b2f4c0ad5a0f324f1773d567a452310de176e3744e5ab4bdaf563df1061ec534d4c6dd737825b89422cdf32c147e71bbbc6c6e2bd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd2e3f0de922e0f408742199e6c0a621ab8c2206f06053ee2a5b95e955e2bc00e84648a1ae7054a38553e473a2a6f14b4630d99812fd88a405faaa0f053d3d3e80630385eb37cc994655e8def8cbcf5dddade07e6a450cfcb5de422e4ed6d90eb5295b14b6423abc19af16693bce947331cc7a2189c46b64fc5de427dbd558be59dabde932100e21d0998d856cbeb23c4b9803a5293fd857bfa5db71d0960a5ef2f467046164d7029a0361504eb50fd36e4eb7ea2244a2e05d63eb674008584e0e72ab03f4466b06d25f4168c2a8534a1693ec149a587b4872e0092d53bd3e36c6f9d513a53abbab8d8d1009d9d55b3163906bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h75a546665cb99eb84b1c4ed7905e18d2f03d2ea6f6567a90ccd65cbc989f2a95db3c294afdb1964f955933e3eb07743b25ec209a3fa198e8a172638ff92b6c0cf602a68ad8d8775b4389e9793e55ff21307ba48eb45414407fde453c241c228ed6f87bbdb4d6f8207e14bb135f25c7fb47aca8ad1628d95c9cf8a643c1b48eb86e137d9165c7ad21e7ca381feaaae70864b1f7c5b4647ccf47375462083c1b42a05c8f6ac9229dbb71fb419e857605d7c31eb98d9b5506beda390b6a61104808331640df9e8ab1d6c295b63ffa10a5ce9b669857c656f98bbaf0bebc9cbd35889398279c6fc25c808d9956fe783bcd88fca099;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he5fac0825c8689bd6d53b9a88f36cc18333ee69c52d3bc44b4a88dc5df1ec97c267e2a3c5a765dde64e130d29f395266fed395b47bc404508a2cacff2d50093a03331ba23e908c0cebb4ada7f981d96f338e78730764417fccc47e2fff6a1f051e6a86e8fd787eac2fbe303cd83b3ce59bec12b41d140370e2f5a65b6e70bc9b6f082e1607f9244c867228dc68099df72fd95f2bd1d66c977eb1f5e60a6d30c7046001c6b1154de5ce0f502301b02fd47712dcb0bda42885697f770acd201934e7ccf96ca93e374deee312f8f4b96b7169936408591197b75c3d82daf221bbf1683d124ac5f5ed865f6afd225d490539ae27a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2af6e737f1f65a0438e3949409373a26adaf6d6ac01de95e4a94040f1901c9a9e46311d41b5593c55bff0ee9696f49a069ea2357fe32858c2234a08e146df7947af61dc35fedfc5342e50f257137f8c0caa3efc51e658e091ad3865761fcbb70f08918079c505a950e6593809fa3b8007631bcee612e3c1cda5cf6a335ff59fc64f98e11989c853869d4a7909f5ce0fc2cdf0ba69adea05d21a8b9f36e7909d4bc2b1429082e6edd652f37e99b02a4f4511a0ab8fa89ee1edad79a746d4e9072512d1d691154db2e6d530200873c3d912551c6d7c3b08d70d08333ad6dc238a19aea68d85d6ca6dfffa364e98ac396c1c402fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h42c50c6f896c0b30c579c8ab2c4bedbd5cda407f1ddf7f30fc120c94a119823ca09bf219b9ed9ddd2c21a3952398142402a345a2fcf765acfb69e62f0c02e2b2b8b60f675a1051cb211b2634857c680b53395eaa34133ad0781e3be9e62093fd2674cbacd07d1e961e363d348b57ecfcffc5bda2a58add3bc1626bad1e973ca1c49ab326f5a48c57b1de27fa0eafc963c87075b1cc6a13a01a85e73a0b1628af3d06f19482509dc9df43f5f43b8457323f821b85e5531abff4fa9d1206a992934a9ebe1c1dc3fdb635cfe5763ea0402834038362aa753f30e90638a7478ff403a932e8b7bb4e01a5d86124e148502f220ed92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h8f439a3db58561e9d6ab25b0a41ca66d0d8636a1ff22b7ea99b2b72f2e0355a7e0df3000944bcaa136d61807266775c5a474d603fd793035c9e4a9667731d69161b854494b8dd8621ad99eb9e197f72f0130fcec52c4f82d8be9bc829d06a25dc615bb200503f2eca3f9317d9da4a9f829be3b75e4cb250ac3192330d3914486a96e0cd7f01de3657bd78507f4f771f412310d5e6810eb44ef8f2da59e889d0caf6ae598fb03c19f041ebd50ac5a909b4646c561ddf6833dfc542ca889eaa12d2423222739e2348b951d29225ed7570c08ae1acbc71a7782b290e0a97bf0a277235ef00bd0bcd931874f483d4223f8f07e3de3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdb1b965163c76b60008432b3f1e33b34c1599a3516adfd3b8519b7d9cd9b203f213e908532254ca0e55085b7d947e3485dc04f83acedd20c3c8feab33ab7dcf8e4370e4acabebdf5c85e2dc73d461195957b0f884cebc9c50d21fe1c597f2716cdd50198e289589504f8f7c849af392b8823e287ed1fd785101b7e2a6d5015d7eb823489a01026e48f7751f58d0cd4c4c913a021ade720afe84ac71b86ff6afd26c28110ebbb861bc990d1f32b1bf545de5707cca72d213800b42de43629b064a15db5d5e75a909c9142ef96c07129c6ca728b264a7dd3c477c153cb15929b349a490127a1cd97e7267e9719dbd76f405adaa0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h46be68b833a79dfa7b7c6deb2b3d3926233617b62965483c60927041d685e44e747576833c7a9f72cb93bba57c9258c8c09a5dc71bf6518bd0c50ab18d708afe6bae49912a9b8b5b396fbd954f0af96324bf3274404348b401db09694dc0f70b64fe9efac9d09dad3f35dff9d21c0b91457609c05f85eb5b5e45a96ac8510b4f69c35abefd56ea935d99cecc4b7234eb2a6271983d37c5d4654abcb58a84be4fb09332a4e026a831ceaf26cc8f2e3a74964b056d23982d1216ba7073e3a71f99da18bda17de43fe5b342cb50489837df1765bce7b367b1402823ab3360bdd89ad20a5648d7e2d75d4e84f1367b3a1122292ba4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hccf58b0599a9f399c372ad4ae30b441873119db704ba4e3d8509b127bf9491e8fd432274d0a4dcb23285fa3dd379f1576934631a1503dbd7acf6ba0adf567797530cb0d3bc8d678a396606204eed2d1024118463f2f3d1ee39ff0a5fed929264874e031af2d986b5bcbb656d85fb862d3999281bb7dcce23a9d0c1012733d8cc363c4286b897986485073602e15494ac08e5024965e04482556578d34094a58b2e51a4a4fe6629b2c77c5c808b753d65a5a3d39073808e2fca91157664d97b83ff4fc1db3bd21702b805b72eed50495e1122367c7996b3ec1626817bcc09920db5e0fe1bbce14e77eb5ce109953a68b9fb6848;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h6cf40f5296deb212a1e212d2956e59b74ced8eff3991411978e53815fb9872b24cef2e3776c8d780d730e7b1fccf7723dd18032396d0e7c0b2b14ebe32f04a5b751bd434ce78a684c1aece760fcfa23cdcdef7bf86a8685e9477dd60399dae59af468eeaeff948e98b0c41025a4ac858f56d64a771a9df4c2e4cfb9ff806b7bf27dd950dcd5b797a6491ed7f272a5499654d88897bf0de66ac6a826041ca5293eea64289200a6243999b0eb2ba3c24806053b289e249ca6bdcb3d4cffe18bb912deffd7f09101995dabb2c900382633b900907abbe3b4fc2124793035e9991381ba6c1382fb170cfb0c5ecb0b6ba5cd8c84e03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf862acdd6f33db75dff00903911923694aca4056ef034dbfc9051026496721ca51b0771b4d4752b2e0aa2df069427c09b59cf65e116923127910559d593ea301b498da347a825b32ddbb11058c39a5a0aa75ce6b68a907e25a2c3fe321f81bebcc09725aa91a293378b0f5e3626e31e3c83cefd523d33abaa852bd27edfd9a0c577d8be6762dcfe1f6f49f82126654d01a385ce69194467cd8a07eea564b7d912190816c7b6a14c5b959304a1251b32a3a5846906a780731b17fcacaa58dc90ab4f1960ba46dc6facf7c4d1d50dcb2706dbaf91b20994e8cb42c8bf37624d50371b9ada1f14d082e836f81bbdd00ce1b8edf53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4ab3403ac504c22c3d5a0c6e7ce3f802b633aaf94e4517be3d3e620b61ab9c161939f4b6696e01a9856f8d43977bc0a65372cf8487a9678f990e91173c7264b877d19ebd4576da53759d6c3ae85bc6ef718f3e86d2e848f71dd3c50120da51e66eda0ee5211a780d70666a18870a8cf868adcddfc79a54812592429eb6e44aab31260cc978e429dec7a68f2a593f1ee3785c606466c539b5907353a16fa5a76c40a1ea6caba83c05627f071a50bdf0662db56be1a375ca0938b84e37ff2e623570374b5cfcd995508526b5610bf76810f9ee96ed1cfe11525231d412cf52174018dfeb4e7bf47d93b57efe04239e062f3c583c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5dc539c2e396474aa0a589408e8081e6b40fa59a10d64389aed217e5e444b9e8fea1b24eac8ba803bf9cc2aed57c1c8d141d3a7cf40a379547f203a890d04d062835cb0a51b10550c03d6f316420ee610028f6dd8c11fde04cb123f76abe189440d9e02f1b3fc2f166380d5a9be46a04da8ed8bbccfde7b6ceee751e37fa6ec28ec0c19516d8b9451e0bb5e4bcd4ea75cfcfa499c54cfd885dbda11b9f70327093c59d2f69d03e6a4ceef07c749add3c1fbc82f77a15fa9c394b4ce875dcc517c73ad480a831c5c642e75692c385d4fa64227b4345b79694020b2d06b9b03d92ab322993ac3c1d4904abac8fba9cee40531943;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf094c34671fa725fe20942f164b974e40849a77b24850b6b87dd5ab4bc6747962d06849734953499510994d262c82c48d7d31158c3462ad95f89671f6e2a771dda13fa826ab83840c15985b5cbe8c4d18f905a88a2a113246f6d0e2206a6c84bf8d2a2e1f526c2386b233e15044f6b9151514f05ed821809f0f4c6675849b8f290199331ebc5047dd85668e22db35af5ed55e35258245a05ba895668e9b0c91a68e573ebc7fb714c222ed5052c896ebdc83c29d879d1366aa0fa74a10f6557710a583c5ff914ac348b1588037a20928f6284a698be9e7b7dc383388e28c341e95e24d1c6306ac9d83251246238ac8130ba4515;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h15cc6c1403cfb4fddaa9cd7274d98df273b418654045b7280428a2083e6aa0fe2b9847f8b59b90f941f7c8ea5ab0aa3798fffadb1be03de6ffed694c23634ec750cdf2453cde17e07d99a858e7a6c073a3de967a1355add2e1802b32a3d1e71d9a8f69f3f38dfca6b8671f25b38ee1e9099d154c296bb8aceca35a81fac00ab105cbd312bd113df25c0fafe119e808c1909d5710b77596de2035e87ecf3fa2f9a3dbd371b7a34d6571cb2003714b36372496d793aeaa012b475886d3b1d99f09e1d306536811a80719108400f07c64840b53fa171e33febb81f2d4f54d6912b092ef1f11ea60680aedcded20e10b2024d2aeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hadbf31aa790513270e0e5c63a7b87e2c7ee0db4886b5bc7c9db9d57a74e36c8d226f27cff8ca21ed80858ecc679da7b2b6b530f17dd9e114aca06ce8e9139bf7ba8c1363d39b80fb2207fcf6fea4da7eff72fa0de5940a7d830d57c98982477f9ca4468fe2141817336f6a4ccbd3794cf16dcc45969bcc8bd33e8e35d3581749871befbb3a76eebe5771f1029379caf9721c949550a7352b6f422a3cf75e23a649f57da0b548fda52ce61d1b8847ae07e039c9b6ebc87819eb1f4feba272475f5f9ac701b30da50f30388e844266af2af080b9b907fe4b94976b6d2e94f619785d0974b24a762f876d266ad94c55b8baf326ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4b958804706ab0788c76ff6db60e07faece4f182ebc6c70005f4aae3201a1ba661dbffe1b1a7396100ba26fe485608b1e9f299ff9ac0239e671c61cf931cc1cd9a8d55b44cbc3d3c80349aa9b24ff93d18fb76279f9bc5b0939a4b334e6bcc1c988ad8fe7fa497e6ec0ce5623cc7d1f02f3b49356094d2b91fc224d088c13ada78095150b790e8234608673e574c88dabebfa28a803b73e1ff31f0eca9a7b5bf6ee8aaf401ef2e292eaec37df51c49e6be23047928321f645daa5fda7dd1315035d5d187a35f9cd5154d807159be598cca5284a4f18f6a3ea3163e19525fac3b6ec4c5d6b4883b0326766688c83e896ec021c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2a65e64d90cf4ec0363984fd2f3c75e8b9364401f77d552c30983a4657f05a461cf9fa6389e8c1f731f86c140ddfc8b9a58459e9dffbe4d778fd90b9f60f1cb712e51073d2569ea07f2686f75330a0cd68234d87fd779bbc4ce08ae67d7bebcee96c4b9e2d178e7563cf738ef2ed82729c582936c3226f39dc620c7e19bd9f77d504b4853eeb266a018ecb2f14fb83a875d3f0e05db122c2464c998cefa185558d6f6446a7038722b2b5714b3e47004219ba09e1c4883120d6dc7ec1a140e2215dbbb124d9b27a007dccf8e5f3ef188bea5fcf9b97bbba38b378388170dc0bfdb5f65e2e96449fd4fa7480d3863187c80674a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1c071ce3be200d8f8b294cd47704415621caa142ddd05baf0c81bec09b82a73f341ade779ed55715e371262fd61cd0483e19769f9b039b40be0f83f120d4893ec5353722f89dfed29f45a1e2050301e25cbfd41ef9dc72f7f67490296041e7da8159891d77239b3111854ba14ffb5dda478d2c96f42b6acced9fa916c7e8ba53ed9ffd5239e220b630960e23dd201b39378a9a58421bd6d87a7d88e8c68d40fa5a210c69193a6d83805cdc8c0a4688da74acccff767406b299373056002739f2480b25953037ecf95d6c9f75a5ac6cd2271f185efb0bd4c3bd79157580b7cf8dbf2eb8878f668f9805356f915a75d5a78d7e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h11321bf5f4296fe9562e279022cc42ef0fb6cb0a230526bc91864fff146f06a38cd08388e2d41a118c685fe3a4dc03ab55f8c9d412f68ee5b61f2e796af5386b460fe534097ba224f9e29e7c25c4b59b14bf1702d84ecc16d6e91f81cde7a5c2140007252ee4a5a15f913499bf196b15fbcd85d6cab798c5ae826e6aea6325bc3598d23dd6433addaaebab0f7aad458d3f57d0cfe26b2c5e5b9b50a715dc0b67301380c95d2f87ee21ed66d02c8db07ac7adef0ccbf1cf6ecfdf7deff4deba5016da61dfece69dc10649f07c3e6dd074efed9f85be819f7864650f44a563ddbc838ab69a06baab6aec76fd50ca1189dd9c9f61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h926a79bb3d6698002ccb527eca7ae0a3618d0c197a82f39b7aa3e7e39782a90508ed0fb26dda4d03f83d02fd2e5cb0cb3babb96db8db7cc06b95d5b3c79f1f57e49984ef758703b4cabf29b0177ba46b638214483598d739ace2f6d95d51f54c8ee41946c59222740cd08dc7d10abf623727f0583daa94e6370eb7dfb42576e0a796a3863dc5ecd472651afc480bd9d555c849dcf42896211c116093467673cdb8f746a85b3cb565619d08d91d4cff77bbd4fae9430edd78bdad3adbb32b5ebb505d6fe1c6bac9103e5d84a259df9844ec992ea39e2cf70525debcd7bcff16ab3dc680f742d232cfea1ea2cfa0967bc89476d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hed81f44f16c8b53d76295401f0cfb334fd5e0ca1bd80515fe73bc2c88cd9b12dce47a76005206b36e2bcfb9af6dab1cbbfd260050a6cf49f54cb3897ad9f1b8336f2a43744f4f70354d4db470afecdf38f77c281abaa7a62f8c1a26d6d1865da35ac2108bff380d604a3e5e9034fa680be89e5956bf6ce04af4e6067c9391c2135e4f1b9983901b88d9eafa5621255a895d6fdb2a5004c4411ac60239175122c8af3b1b0ce0820398742e4a7e61166dd2180c5997294c19903fe45b9621029ace7bf508695d1d02a6598a97246e88ae275aec53e689d68f41b00c9a87162fab9e76af96d02a1cc0996299e487b08bc5aa12b95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdda3960dfda12a1f2b658230a87a391eb11d8342fc72acd23ea1d538ddb840bd6b15d89a8ade63c8646bfd35913a71869e522ef80a53a912102db5b8b4bcc4886ca01082460cf335c637ab8a099b4559c76740af0c224d1d642ac38a088e4d2bd2ee055c1e9101e1a7ffd0689c47c3ea9f9e07b22288969d9d88ce350263c0be6de29be8c01f90c434130354cccc90a966acd6bf9f038831fb4d302e2b75fbeb3f4debc2249d2a0d7b9b4181e4db5957ce9bcb01835b57cd953b7fe896cec9f8573f7cd9b7eb21cd6f28d85046a8186a61766be11c4122b0203acd5f841c0fffc75f248912410eded8608bdf95a73d2b9861f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd8d453213f9cdc10f533929e4a45872a9e36d80fcb61d08ca2e6f9f1a55dbe93283676865ccd17a9876d684b84d7c99f5eb2f58e2a61bcc1af94225c1bbaa439f8ffa76aac63b4fe4f6d74a7911b16d99c59426266b262e404fdc2a51ddd3eb2f00610fbeda8a4fa2ced70e7ac61154527912c30ee8282e7cef953ecd8dcd4fdbf8014182b594ba20b3c0fcdc45d5d40bcb80ce67ecacb0625eac3731ed543046581c25dcf4bbeae002e8f930234179b408ccb8d50ad1f68e93c7a29873e6372f1eee91b63235f6db7475e216689240281c0afa9a114bbcf88f4f4d2befd23c1951f48cda385c54a1b7f224d88542d16f4a072;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hefab37c1abc5b32156a47980630d6912d34c5ac4832cc4a86c73de3d15259eced4d2ad7dec8179d6b996c4d291e659a876b5f2e474408bf116dc8b1a96aba55a54068dbb51b11fbb54fbf426772a6e619ff87880bc55932a9103470b79026624356d15c00e7f203a06b5305cd0b2b1a0a7e5f96a37832be03dbd171211269de88e0695f19a441f0f2119d4a99adeb82f1f46f6eba7c3b52b29b7d75b339d4d0e09bc63263078c62311cd431a7a88467f6d956ce92fee4b6ee93ce1b423961017ecab6836fe0a0975a36aa2924d9c892d54e973e138e8c978594f9c6fbefb8b94c307b0c636dba1f67c62ed86794efb3802c96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha45203921d688b4c6d5f01b612ff51f3d19ec0d268bc2dcf8df810d19fa218b0313c9e75121d8d64f75fcaa83378a821553ee8709752502f5d242cdc833e2e7119d26a6fc22d6772efdf4192049f39e10b674841df43d8c8962ea9a306806be4267e0bd4c64c148ec1a382617a01e675750a3e598ae07a8566ebb97ea7ab317ef456706e6667fd8cb1050ca80262f0390114011c6187bb0342296543a008a2dd7b8624f3b7f65f101e7f6fbcc93b03737e2496c7ae387cc963bb10319850266ab0a5c9d1a2f53545a88a7e1c8e7b9c91cb5f2505206295777e1975420d92c575bc15ddb3ce4d8350d44a2815edaf70ee0f1b50;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h89340229951f2a1e832e82a44fb95f57c8b9250b47105133edd320582665175934199476765b1f6acaabeae933ba261592c469fc7174935cc9cfff3753b4d58ab9f085f5b5d8b59a89bfbc797cde3572a36105bce1ef8d4a18af48cf374d927abd386d25f57e929a1fcbd61a6b2b87e7deaa07895db414ef8ae888b15afcdc1d84e48c14049d5bf48ba664a604db3257ee4a558aeef4d220accd9ee8d24af4315efe2664ea5465a5ba13443cd91b2ad158b690d654f75c2d7293ec753e17d8179681a8a624b5233dba8036a197a1769bf5f420ace344b1d55e7f2b1fb94bdb58848040f95398e54929c09f7e1afbf5540e95a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h8255880dc40250719d2db8ba1b7eed4d44a0b8b9429ffa33236bc006d871498e99c7a1257b878258491fb9c0d225866cd1686fc37a79b4505980743e50671ceac2d8862791c9ee532d42df6cfa989cdfa36a761e80031fd3978d407821c066fd8b7862cc7b46a7cfed2eeb018f670ee70564a6a5551c62a4824d2540bd5f3df0e17942a81abbc33e380d3f2f29d0b3590827e14930684e0127b2479b7c272f43b231177a80f2aa745b8f74dbfef6e36c93691530ccbb57f142567d590b67dc7a4a9d1d85c6596852a38286886e1c37eadb724e07061d7dee4c948a59f7fd1c55d2d92655af1066f75e70df49217bddfbb45da8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'had6506045ed9e908e44001590f36f7ff19f6dcdd27cb70a7a148951d6d565be66f166bf113ca046e46236cd0abb964591a24660cdacb3519204c1d127b91fbbd332e3fb9a00f25f84d59234e35258d86806518e1b2bc7621c8f40885073847a96e8a52a782e0690a24253787709dfb4fc000e3edf67c42d754f542c54a30a09c306c2f897376157464bf5aad6025e93367a696cab64d407fb90267f12326cc775e0209480318ad42f716112f5143a8bc87da0d415b42dcaecb1c4edaf519e8c5222b4e2c4220afd15eea1f4cb4b79b840121e2d95ba4a8d1d07bf7b1017786c5a9707e0799d551594e1a43fa0aeb50e54e459a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7e8b53418cdd839edea9beebb690aeaf1faf3a58c443f7da0efffc4cad185675f4839de8251360c74ea4c900943222e57e1669be00c0baecf486f7dc9669363a4f2a6fd3c88a07df2533d2e6a23beec3fc2abd38ccde800917ae7dfcf0a7c74d6d2c8927d13eaa732a3dea3713d48d7a625e315e81f727f4d5ee2496363a9adb488aff42c7e8b68e121ac40cc30a9ab5d13aaf97e8c352a24f97ef11a0bcb0b90678fa127a1ef72ced015390031fc6991b9dcbd77d7d0df0856db9b247df9b726840f16db328aebac0df05175cba6debcca2f12b1132e0bd08d4294e96e5f44dff4bfabc6b9437c6c0fbc0431de18b724ba4d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h44f4acc73c05fd7fbc7f1a81cdfd4631a32b8d70ded7ea3e91d77a85b9b2612b4ac21aed2faae6a30fc533fdfe6ceda8bd66a493cedb2e2af95b5ccc1c865223eea16b4d181be0c7346d262e36291a68d6c7d364f55f7c40f8c10ba77e94b1353a40b6b878c008beba32d8e1b61c04fff12a78fa4f6496a5153edf645fb66fdbc170f64973dd3ecad159b1acea253ab7f475695cebe8a756b80a1b6281e640eb4e697f8f33b15dd13518e78a8699bd417324bf19203b3143318b87a01e181c75b2914d4c2541de06c36ec2ae7ff165f8e071b6a8c42ebbbd295034b4d8ce527f12f8f834fab6d63b67d7a9b4ad69454a7394f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7b1cae9deccfafdee224019502c9c3ee858c34a53df6a4133669a78cef8a8860b2d20ae032abe780a93d844caaa7529b24effcab5a3daf99287d16763810a5d9fc447727888458ffd4485b0ef07aa10ecabb05acc2bcba1c5855c944125b990685262bce2fda9a28e1976d98f6e1f67e155241270eadcfc2803395c29cc72e72176a090864b4595baf643e6168025e456efba6ca37f7c292388914e2f07957bfa6b66b0a803e25850c0649c18010ca2434ffb207397aafc4189ac2c6d9ec9aa920b682033ac84395f7bc15eabe656beca05f9b2c3c2f949f0df14a32a248793718a7228c78dd18cd13f6a59d53175adf085ccc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd2b7210bea7e63bd8d45aa81d2548a6b9866a9f9b958e94352a0ede588ade93685668d47eb75ba41f9e5093ef7a8ecd20ebdb2998812ecc3c2eaae5292f3d9f6f7a1e8522d8c04e9a3381a10074f80ed41ffc7f89b14dbdb6c6cfa287582d200e47bfe653809014fa5febcb73a8c03625be8c8b6ef65c8841b6e9c38a31fdb59cc74ddef5b5b59b0ef2c9be747b0745fc4f86304661e68bb417e8795a4b969b742b3e0c5b59a108cbe95809fa54836936f363d27cc7af3cf7f4d19575197e501dfa2805fc57fd9d76ff3e17ec078da06414c3bb5efdcaf7e4b5b22467e72250baa7aef059d510a736557ad6e44ef8e4b717d4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2dbcf2434202ad7ecd810f709bb9d2094a5afe48def2682fe19e99e7ff1fa2156bee7e1f5f504256758f0389ed59b3270284a5642e078415ea39f339908f28c7b083cf7be53d3a48eab62b00afe4d09ebf37cd0e03ddfa14f0078d79e8cb169b93f07f4e90358049ce9625391f46d9e8e958dcbae4aba8bcf59079db8d0679f5f44a4263c7bcf8a5dc3383b8083a36a7ee3ef223415bc59d9681c597aadd1e11d51368b7931b7cd7a0958dd51c62eec63a1cc7304b41412c8d05097c6ffa3c33f890f003e51ea582c75bdee3fd0f96d95df8aef01fe6af6e362d463abe53c381426731db1b886346cee123839161b7d2acd96c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbfb7a91bfcb0805200116323fd42a6db1be8f294bc48f77d5f749b5e493d5a6af0659507add4161e0861f404e962769d707b5b8a0ec4b667e5758d538fa8edf1bd202b361d0ac5642e0fd9b085e4f790c55845b18cc9c5e7bd66740a41b8cdb374e302120ded115b2d1ae75b8ec409d7cf729fdd722359e67ae1730d5b90c75bd5b428500691d1df61c31b2042c9de2ab17d0530ab286e20fcc4d63ae01818ce61fb0c2c0275b22d48813c7de15f2f2d2bcb188805ab67a758c803961a5237823e7ef1fcbbd93615a29db2794a76e1d222c8692ef936709c2c20cd2a706702fab29c1dd97b434e7539b70df497c9e47da061a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h63717f5db0398de4f01c2a399ba78a63e7ec363c31bca5346ec4f4fec4fddd31e0ffdb00fa585494231de828244d1442dfd5d2f53c6632c767dd2cce7fc2715b9790d23a2b2827f72d51270da13b35f1cff8bfb94295af89b39153e98ed22053fee638cf43258b4c2856797e0fb4dc118f618522c55c42d6c8af126462682802bffef9c2c7da1f6b2d307d4fb96d50c7b2694e16311f7e1f50392ed7e3da1e657262ebafdb865bdf3928fe7938e5532e762629df7d4b875cf20ae4868f34f222903e733930678305851765d4f54a28b102e74af0ed7051f1a1760250df4a69dfd56d3806d5fa5cdc4fdacfe62c74645d641aeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9808ce558690dd2486d8f890fb60675f9b78e6e2fd2ddb73412a5e9dcfe2e70df3ff99b3f678a151cd20da1e5c9c1bebe4ef98203beec5b418a0e0a7c3cfb2a99696aed94d5838954b5f4b9144b5ebd0a7f2a5a6ca226d46e2336d4742cd3a94548d06fda36417ece574f95c00b055370d74a82adbe2f067f72217a64c468ef6373e0f5ec2143c229e25664e13aaf83c5040c5d4d4d83db7c901d84ff2009e9dccf27167bab2e5cb0f22bddf52d626fd05f3f42a35d46af6f86d3151f8071ff6877e574c36eab94a0df59725cb82f1079b3a64a6d71c6735b4c10d4dd442384826b629561285c2dfd210c2dce0344430a1df53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4420c3cbcc2e5e761a59b205e022d4d8eb8f67ab234364919aa551bb23183ef2ca0981936b90de86d94fb7e9ef6e6baeaa8cdc0851a6d04a9319f508c49c737c7e4071af95250dd3e8fbb13d4345a12d15f3bda384e715858ef7038a2e885d48bccb9b20e9b7f9bc3fbd1976bc3e3eb35c68997e212ab6fb6a1766d34e259a0dd5aae6b1041fe11031d55cf2cf8da7de6ae5b4b10d9785459a21843a64710e2676e596757cb1d9d7f44387177fd945e80af6860b93337c42897134fc92921aee6b8f1f4c5b0855fb3efa10ae4f87a7e9188a4dc544742d17a3806368ca8647f1dc62f15faf186f80665143f1e7180ba6977b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4d2f7d09770efb300fa2a113272dcc21280fb6c8826697957ea17294b20996b19928e38c82f8346146040ed0a84976bb6de11f932862206c362e15305ac5075d5cb60ec3a6b80ab195cec90459c43bbbd5736b5405d0af4209a01a2a3e311dd1c59c297e0955c9b0951662cec64d27a506fe8542a6b731263e0b8c9546b56ac7f8b38686b4df4656a6ed42de023cefff63dad7a9fc72cc2f2aca121b69ae87072f33ab626e9a043d34a9c3eea04446c7d9b789ac3a802e33c56d44783a0e0ec693a08b1266136bddafb0a991d95c79c0f92dec157981e6709124abf7bf8a91e1896702f0eba10e302e6626f7384840ab7adb4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he3024180aa396ad603b37484bb08242150bd4b579534b4062e163ab31c10c592e5de1055faea5d0b6503620552610a130eabb51811595de175ddbce0718e2ced471cb7f28d52d6be708fdc77cfeda423b98119cef200deecc1e959c6f4ced4f2544ad67e2c908f7f84895fd4613cc43f3e2b24be918c1dc69e722ac656872cc604df0cd24af472bf073d6c4c1150aaeed55204a0fbcb847f08815175d55e6c9609e4ae5e588a88abefe9e9ffb416998c8a9ad9b6085ab21687219db246eba6b4c2833575495fae1e7d2abba20ccd08b2370cb7024b5a6b9fa21211bc8c0688878216bade1b706859f4c932879f8f9c88af9d44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfae07ee84319763358e0f5265ce5154c0f2ccc1c76d8e780cb2cd743d9ed070aa7aa835cacee244fb05a3dd49f1c0bb78aa068038c6337a122ffe9c0bb162d8e92163db41df0f499a2afc08084d32ece5781b80f919fafd86373a50082884ced7cc8b3b2c4dc8cd65315981964afb610d99ef82e3292a99a8417ad5372004e7fda538f6084639ecba2e403803215eca3291a6ec113983796cf7c70fa316141756040f45ba5957d3af3fb72400a8a39ed3b64e5c1032728eb925ed422c2ee3677607e07b3b50522dbb637af2e46e9eae29c32a555ca878ae26a6d203bc8e2bdb8e398922b90287377bfc3ed7e4fcb09d46885c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc01d4e484630b55bb4e743a5f20a19f1dc34275246a738f54b97dce0e4c5f2143f462b9e8d8151328b06d6f401c52133eb98d94f23317ff2ef943b0ee764a7b775392dd5d1b9adb2cc3006b404733ffca42493dff573eda5d3dfe05a3dbb07217816a6afc19a5af8262d48093d21e550479c5f2a15d2205d2625c20c5d563c3862aee025219946f6415c3dea1855ea5d7d433cef08542a464570e25ddf4a16eabf504a27cb32bce7ce8d78d79537beb92265c88ec1257050545cf511a6a262d1eddfa6ca77ed54adfbdb1d5f5f6742a6aa5b434c18a9bda44be9c048dc9fbd66bfdcacfe49d7889f2f53975850566532d78ab3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfdeb7e44045cdf78241bc8a17269cd684a7a5f9b93efa08b3ce63010edd4c081cd7072429743b60279118642b56f1870938381ad88e0c86eafc62648a254d225803db4b8866e89fb739fef63de579b13f9b00cc3258f102780cb044b9fe69aac684bb69cfa11d444422dd37185fc2609d420567d1ee28de2c6c796ed3e399aa3ab7971cd5499d288dbf19ee4ef139865057630796a73e574cfb37dcdb4ea4d1d113e141501b0106b7763bc30566334e51f9f96a9d77b95aa03585839289931b8230f6ac56f2ec8d4ff9b984638a996f562d69f73e7e8d81d87000f99fd3346d2ca722965e661985c87396aefd2ab6caa1e8536;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h396e727cf6abe49dc0eeae300d160ce3ef718b6e627ab3977bbe05bcf9463ec43e2e28d6fa48ffbed80357089747d35a694a41ff60544f0eea1f7fcba72a21195714bb3a08d00cbe8487721e774bab2280ffcaffca5d41e39679c76631a87c4c167f455be5ea745909b749938167039794693c36ee2d466ed092e7e48aec12ba0d597a36bc3cb590a46d7d48e737bd03ca7772e496a338ad4538b9a49cb567c97c8d7d85a693273a84eb7de27d95d810c01d005268f2e4c9a1175c6633a2aaf844a882de519fd1a88a9d2afed5aea667c4dae03a12e9b9518f83563a5608188c8742b93b0e1344b9cb312bc4735d3a594a30f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hac04be22259ed6a3ea2783a5c5ba2fbad2b5d9e699ea8088bfb04e8a531169837755aeeec718d6fa1dbc9e43f251f3649255a8ef4494055036e81c388ffbbfdb9c6f2e068aee71db3f4c6f5c732de2306c7d4da735d7d6f444b05c389c4625335f045c99fe9733845b5f17ba645cd49b3cc78d2e640d89821c35cfc1bd1eabfdd0f034a64d38c39a5a7de5aba69cc96fb686308ebbd531d75fc802d473d1952778713fd4e5abf996c8aadbd189d48caeeaf835e6ee450b868367488859f05f1c063f1359db29cbff08737b792f12d0b03ea855fd4e0abc8b79f3a284d9e0ba815f115a0706ca9471679fcec61436ecc391a9db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4c17af159c51fe30caded2950be110f12222037560399f275d10f92d34faa8d40ea64dbcccf00708f4bcb975ba224105d41f3c435bcd867ec75546c0cd7568dba19ffba729e1f7165fc54bbe844ab34ba68c943e6586a3e1cf5581dfb9908a363e3a8e402cc935a207a1736b47b9d9920f654f9f22c84b45e6a614a1a4b884980420144f2aa71585535634a8fd1b7b784b18f231808cb36136a750fbaed7662b9cada6517280cf4d30441ec63297223f264b21128624d29717a2d27d35c1669b3bed5892e013a2628cf0d80cdc01005b224071865d65640f46eecf086b560543b189e71ee8082effcbc5122dcb546cc815279c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha6b899b4dfe6afcce5699878f23224eea2b4dcfc043a9f77bf00c664e1615baeeefe885a7fb7adf7cf9f8df0253bedc34a8500ad3072f4240137d616675926d206ab81990f74c1b2e4fd317fb09fbdce7188131e93c07e1c9310ee39697eaeb401870738bfc8f93649e076ddfb172cb9673d331c74dd139c1d62f51cf23d285665b75dbf9c4fc028639b582815f83b743e1435963fec80a49f47b33c28847698561d627aa2e170afd6da2d75f177840f0d67056336a6fa5be41acbf2a3f0611a997ed85113e873b6cf3fe175a98288c408da25a4c97289ccac9cfd596466e69fb9b6360e01cdab72c6ed02df64cc6d359214cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h17842c6de0ba6d618da835b6f15182c3d6064c62887175bd2396815599a9b15f8e1414e2d20b1eb73ff3a8d162b78e6d587588b76a86fd95762ddf210f149256dfd46ba899e9af3807074cc0b63cf1eb601621d9378920399978ab4f7677bba0a27dd9c18c988558d10a223a7cfc9debf8f28de2ac3763826b48919b9d2ae4e59ce642d4e57d803f54807f7b9d4163f7ab808797cd32289d81f7099a0a399605c7cfe8ae86d9f47c061850bd11730c0d7f347bed9e5d0010b187e46326d3d3a20a9fee646ad06a0e5cd58408991069be33bad5b7dca412806b18448935e57e0e46d61b6c95fb861bd410b8e65135691f77347c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h405731d003f23da1da908eadfdfd5e0dc90ff88bf07ce3ac8ab98b94f5043ce8ad6b749e9c3075ef0eb89c921c9050d8219712227b4f985d6d270ef4cea9356033fad839cc244f7f43bf3f252e5abd448bdaebb745c58cc0c584ede9d573330084a94288412882ae371ba6e56a083f4cedfd63dcaacf473f1d4320c4be5e7d0dbdbadb64068297fb14ab3ce244b8b5f6a54bbb53d96f297d305f2f58ca9f33f5f8c7dfeef6d82035317fdfdeef903d16aade38522b24c9b43f12e007b6a347ecb05f59d6050c20b5ac896af53e00c8337c06592cc75a5ef34c6cf1d1f9ae6ab8e4c316a83e8ad120e4f9d1f8efc5d106bbd1fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h731044229e62acb86a5b727ddd1430f4b4af38b13880bf67f5c84ab4caa8d77988cf29d141879047cfb0198fbc3d7e7a252f495906fc963bd7f77b0201db4bbc1a2d1262cc56da5f0510b6f25fbb61e44c4ccc19a2b4e1befb15790de874545919541e46beb9f22fe41f1e73b9e6b9cb9d9b18a499ad45a4709e85cd45c69d7041c7d020a187c9a5953388005dc49a04fcdf7d684dc9bf4ed9fb1f29622a3829aff87372b429ab70e1351824efecebc750d33c4a118bb51121a53dc5d4f821ecc03c6cb908c6583696d1463d3bde7055af45c7f71bb7ed207fba575838385c73b8584c851a6073cc208c5ba55dc707018c0ee7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5c1e8e95f1dd3a34d1af84542ab644514c8c3e9e0ba123bd734aa53d518e59598bf296addbb77b332378b40b967448b5b9847815d5037839ecf636766ed52089c48678323e9faebd4d8f462202b482a74be09984fa60e857241c6ed6ce5c54cbfdb035b15a3d3d3cb2b80bda40a6e02167986f6343d0c190a754d335d69204ee6a5a8f46ad41bf9ea11118d355928c0d4266482406b8aff404ec3b361b86c45901f3c7dcf4e77b64267604cd99747d60722a1b90ef9fdc5104cb73e6e59b97079d7b3f09efe6b92fea290d372760c9b7163875c251732649abd7c89b415e2a2dfd7643e7910f07020416c9bcf92ebf0bc98afa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2e36dcda701030b2b59c3699e266c1ad336e227c89a49970c8e00b5224544062e1ed2d663b6b228b9ca75a14cbd3362304a3524b7d7f9650554432e1dee30db60b817de8cff6de578bce4b7249ef9f63e06599cbe6a47cee64f3c1fe3c5b32bdbafe091fafb4e1d7552d3cd007162bc3a14584a51e81dd5049c8ca01dcffd6ce38cbcdfa6469420ed0778874927c3595dfe8c5cac73bf9022e794256a9aaf36300632b6e47cc437d00cda17c39ee122adfb602a64db10368cc41d6f4d0b2d87cc7af4642fa213a189093f2eb48b80c73814b70d4dfef884ea37a8b1921b29e2d08a9e24a59ccc6ee469759ead7153967ef402;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hdc50dbb596f2dad523a195a070f33ccde4e019ce658afca1b02dc28e31880c49eabd5b50ddee78f43fd321baeeb6a3bd7e280aba4a0ebc3533369f4aa04d4857eaeabe756fad656091d62d0eac09b471314fe615013bb49dfbecc558ec32080fb5b1b0ec0bd46d017f5e4aa0a68a3652e1b5d54b8865186b996ea163cfe517418191df96312bdbcd4d072ce3486facb48395dbf0f4fe727c294571c8d6c7f75c0d526edaa4df443c5bceff29761080a03663657c0021a78a24f9de5dcacb9043c28b7c386a9010c45ddbacf638b56c1f7b704ab5aaba05f71e937237a28353a639e16a05461f2c0eea614f2a72be82e04d4f34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hcae916c0fdbe70a471f72256fb6a89f19f4d3b7e311f6af903e568d87462ebd5e7c05be0bf43ab6f14bf5c73dcc53b158bf29590a243b9aa0a8d473cb1ef24ebec855e3c61e99992fdb1618e3cf69498222768ee48f039c8e2cd9804882ab864defda162dc442d0907b88bc9d31bbd4d0bd214104e340de38de4c97c98fd9e373d2f088168bf243a76eaef30f12d5f8ff5880db413648394f8d690f91eb6cfa8987664d1e4471c7b55d966e3ae43903f55701e1913b0de1c7bc4340c899fc637cfd05166669bd81a9cc0275ecf39dac6b98ebc6c506cbea6943d6398512b73da51684d3880ac7eb1dbd57e9cbff8402376ae65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h49c9fb05cfec9df6d07a8b4abc9f567f8447fef0a04ab2abcafae8908a69e7b538e9b49f66e025d6bbd4381bf4b436d6c49412ef1e6eed2e88046e4e31274df2d06ccdc801882f21bf4564301f3e7ae8a6aaf23042ff60f6bb6b146c7eea157656392313d1238b3c9973689bba43d1bac41c3f31f96bebc41cebbd89d6f4d7c8836438d7c08947a87c7b39737579584951b9312e8f48d104cec763d5d23b9b9ae263221fc8c9168ee28b03c494a388f6f22092477dc6f204c01f5a589ca9fcfbb61541e8aa2297c42d94f20864bb7d3b2b4a2ad094e39215f5a0caf42969a2b04d6058cfd790084602c9ed0612309e38d18e14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hcf41ddff22b7f8df764a90c91b39261bb99366a18f66084d2dbfc8d84a301bf786db55d4ef119ca87209105056486f607c4b4eb444bd0f917fd7b0ef0be6e6708f1f5d01fa24490912b59e2230e5712d7516136b3760faa310f9169232143b4d6e9c9d603b0d735fc111fff9d4b7bc2e83ec9504fa3cc36bde335cdf869108538cddef8ed17a92b7da2226b885fa2013397a76a3e08884dbb679820cacee24d18a737d36d706ca521e8c576e0ee311f4e9cbb7db970c0dcc1c16a7c32112b511218f96a8476d35573bb57a534b979b5026ebc2cebaef8ba41defd3f4dede9453a164e1cc71cbbc8d1a87af8d515b6703dc6192;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h85b5bd8696cd3cf88bf2772cdb25fdd50eb7415130fad1c9eee8bf5f8e7276590940d43f013bd2025b2dac5c40e0d5e57deb1cbe41d9bc8be67ae7ab273551e11ef7ccbf83eb6534fd0d1a9781d80eb1c0352f3de92102cba794f3505ec425192f300802b3f64f3bf24e1fdff3ff1899a53ae1d21d1d86f455ec76f9a722a300c1f79061dd67551ca5d46c1ea8e3684cbb8fb39dacac2c2f5d0bdd55b58aff1d7a64bc7fca7e9eadd714322ed7b69666f9d4d89adc7d06b54686dbb6f97b492035a5b0ad2e6f443b21f387a00990a87af24ea0377d66bbedbe1d003d43b893bc0494394f687908582e349206303565b02fec3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h949f27664abdf6d0f1c48e1400ab715f4bcdac29fbddae1e3702a1581e0e49a0f39282df37d824dc1429e8dcca9a651b91e867780617a6308cc8dbd24fb2c839c3c444c048b7d61953362848779bd7c3eac4c8d78cfeef6ac613b42b23994e093eb58f6f1dc633f867c1b582fd9c25324ea921baffd2949c091ffe3319644c40fc1cc61a8a0b00f90f63b1b1d4c788cc28cbaa175a64278d25fd322fe60e3655b21091f4d412fbb509f15d1219ddd6cc368b9a6588b59264a9a934cc33008baffa5071f3e2fa9c77316c8fdb5edd69976862ae78f13b1f892271bb49ac744b294df0ae53545972a09a74a2e526c5fb1d5108bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfba6e5d1efc1438dfd52b3161ec60770359079add98af1270eef195c7402823442dea33733d25ca3ec61f14c0e9bd477c01093d071ee11514edcda5a5693bd3d1e78cf4d56ad691def7c8c4d6527b42f505d9496aadd3ff16054e3f6d53c5005c1ec0364b4afd5fdac47157176879d7a98f3a00668b3bce16392d809db0e6cba06980d0b1a3b147dbf5c6cd68880794e46dd68c300cbb2ed20d5571a7ad97359780408dea973400e51694cb18fbea0482d19150ff9afcbe20d134a31f08717d0fb03e66309dcaf514c23b4c0b65dc173b755a29c36d98bb624c773ba99a519d7d92a8ad9492f52a39b938c8aaf32091f2c88d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc000557ea174e9476621b71dce8079b72ed873158d1ae5e764d766dfda523b0cb213844ee3347bbd92acd4657c62e5d1690573d8539c87c70a4fb622ce6fdbe9d69aa2d0b34b5e70cf5d2532394825332f0dc4903936830ec6bc19d71d58a4022ac7cc3912221426594f3bf0da219dfcfd32ea41deea892910ccbfd2903e03e3f7d73bddf7f2c6a482a16bec9c5622c03e3cf238ffb8bbce319f2ec7724f462d1533854f22deaf13b328b830a49c14a394f260726ac6f3454adb0b2e040b6996562142c21d4990307c6fb71204950141de989a6ba442815098f5a84d8d1126e52fe432ddac6e717bf5ee9ea7f9ebf0e3b09558;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1f704e5e657f8231b5b57c9f5492ffc94e6e0947e4e652ff94adaefbd09c891b19f875b5a64bcfaab04c0f6566a369e65036e38a8780456e95628508ab9a8b23eeaa1efc32bf96567ccb312575a0cb6b5b688c082ee393dabf98f7343c034900586ef8d44177d96e253a07c7d7457322d72a5650c60b087ef702b417d774312d40ffcdef797abdb30f24dac3d81d49a7c17769666a44b5e7e9400559dafad3e40408b025f19ef4b7f568ea14c59bd4032e7b7148178a747cee54be76e4c2a2e9e5f82761b18807035a9d1af30a519ed848b3852c646538f58f48f66e258ac2a2f1ec047f8d3dab389a6783146578f75d784740;
        #1
        $finish();
    end
endmodule
