module testbench();
    reg [25:0] src0;
    reg [25:0] src1;
    reg [25:0] src2;
    reg [25:0] src3;
    reg [25:0] src4;
    reg [25:0] src5;
    reg [25:0] src6;
    reg [25:0] src7;
    reg [25:0] src8;
    reg [25:0] src9;
    reg [25:0] src10;
    reg [25:0] src11;
    reg [25:0] src12;
    reg [25:0] src13;
    reg [25:0] src14;
    reg [25:0] src15;
    reg [25:0] src16;
    reg [25:0] src17;
    reg [25:0] src18;
    reg [25:0] src19;
    reg [25:0] src20;
    reg [25:0] src21;
    reg [25:0] src22;
    reg [25:0] src23;
    reg [25:0] src24;
    reg [25:0] src25;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [30:0] srcsum;
    wire [30:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e507f5f0baeb7423df906f21473b85666322603dc5db711e3524d05ed3ae9eeed1415ce03b670fced08c6fb1f48e16d86e4a88938c3e6d21aa24811c6bc224c0e457beff86e9cf5388420d7f5a6a983fac9bd070;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6267293f8f9a1572fed4913747f8c2d943165a4c99082fa6170dedeb885b3f11ed09bb0078fa2b49f71d654b5c698027ac08e7d02838bc56ce1498d0ef7470bc0ec3242729099f0ca2688388cf2e5697965fe157;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd11b9d35d7b2b22e78de61fbf49310dbd042315c6050eefd2468878eea87857b2b3198bda9b1a6d6aa33e2704fb1577ccf9f690133d3c15140b4481d47a4f518483b4fabfc59ddc66946497f2a0682ed440751c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6ff03fd25b43e6e7a27ba880202bc17c23f0208f596201ee29a0b183c3ad8e0790aab47b29e639d3cb538b243257c2444d1f212f81885ed5682edb39f5f63ab83737c7f8b3e47e149cab3b0cbc3b267f3aef8db6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3570e787f3270508a043163cfafe27f0a85d51506e539663c32a8c7832d1c324a637dd036ad1596c18613841daa82b88d833d53bf656df48ca8da90276106169827c859d9315b63d8d375b26e839be1fef585a4f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7a3cc29920d3daa92737b84daade8e0d4a37a83e576bef197a0fd9a23e8a7b11aaf53797b72326efe1e4c898a937b414ed712123aa95d6000531117476b86d38de27444fa904d3fc7b7416f2d87eb84bffb81c74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3004fc6c7d0d80cda36b36cd7b5cf99f51e56b3cbc655d073e9500f47be2f079e7585729095e52d82a4184cef0793e2f2bd71db552ac7546224d6c6d5ce74c4ba9eaf84c3e5493dcf2f741da4d9ae9531fc156c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde3fc1f94340a59a70982a1a73669adf6c71c070bbbcbcf926bd4c44f7b6edb598163e107d2153b05e8828dc498c592be485ca05ac766eceb5ea67a3130bc070d34186e17e98aff8884cd972a3aaffe6fb3fe58ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5f7a22ceed5ae2911efaee960269e822238056d3c5a1cfbbf12d95edcf89a1fdf709602336fa40813485beeb31a97e264cace32bcf5860efcd2ae8d60681cc2af5a42aaae6ba0d7072006271ca6eff4a461149b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2bde9f4abc57d72821fb079d57ccc8108b768e6be72401e11add59413737d409ece584b2530e53b2404881ca87379a59ef34a005f0931b54eb770de190ddbf346ca37cd4e1a4d60fe8315c634ddc3ea301c8fa22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe8145bb9aef4795acc53c1932ad77377920976eb1e10d481131a8e5cb109c1f1f6d45c3c24ae50998626bd8b0580043e2db762c1ac464a01caa6ed1490ca1f6212c5ce932569ef0a2473b5b7b6b6bcd3994716d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3edfad7b84a0736408f598b1a255de8fce69dadf93bbb5f7169e7bbd47327de3fce5ffd333e39853b1cbfed739047b156f24f14767c7729c588fc48b6bb5f3df7c23fc1b830ab1b2d100c1034a5ad1c3511358f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf80a9c00b271b26ae61a711315db3d02c240a906b6b6ce4128030a53a6ddd9dc947cb56b6af5fa56a5c2b79fb93c1ab6d3e3107ea6d436a6db9e8811a1ca33405ef91070495c0f64a86b90a7fbf6f9752ad9c4e32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha811e420226b80568142a102492dd49890506be077af2de85d0df75b09811dfe43471889a8a0fdcbd6555371ec9571807c1c1e450356491beb32ac4be9b1bd99c0498483337c23484418157db08e7097e179dd646;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ff01eec2f6f99698bb69fb1f821c7f7cb351a8f9f8487b87a62092cd66dfa0a37dd7839b01835002fc2540c50470291cbaa600ebc5db9b32478f31e4592f12821f5fa309414a440aa50ca1865cdff2b2e371d675;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2af686aea73cbd291db9540b48edc5337c63b13526fc5f2d972ca36be31a07679df190b25b5debbd8e6a8649d327f3c226c043d37609cd7552adb4d9a461cdd46c03a687dabf0db43fea1632b7f738e2166bc5645;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf52658d6879c532e9cac88e4bc80ee74872b685872a224ae48515bb8b5b2c0cb53ead27e30a3673da760f14e72c160c90de00e8ec42625d722a19e5fed554c1ee9faa6ce3a875e80cc7e073e7d8064d3128f124e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b223ba79c1fb0d737b71a6568a210012f4cea95e753f6a292e04175495a12753ad4465f72f209ef9655b8a3951a69e7cd60ca114c085d2a2b9338c7bdde86f445b05436a6fd668f13c87512baf6ecf5eaa0b4017;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ad8029c8364b1c9622e2f03d1034e964df9002c14f5ac44e85110c9af557c6e5e3d672ea695c367c7040e01500d7f2becb07956d466ae70b7e9ece9724416420ba0da5b43092e2ea325298c1a7a68cc49990c322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6784c20727b0136c1dcd8e435ab957e2468c6abf2a2d9031d49248d616dec3db9693a6c15cb35038e27e21a82f819e621190b6a20942400301bce8cf96e62a19a8be23d587c4d9e6e7affd30aa0293b2221f38bac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d94af280917b4484291ae5e600a8e96a6a17879a0a2cc971c73238a376cb91b4cc9df18bcbfb96f55993413237659fcc68ae5b22acad6d4efe983a331ec79c0f3ec9aece72a0ba0e0d74d4d50288e0bf9cf49809;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha611650cbf21d53e499c689b79ddf6392f52c0053a7c4d1f4352fdfd2b4fc9e3c9ba362db25769cceaf22fd42adfaeaa8fe3e02f5e8bf84c048ea0b9bb29a4166a9e9a0abd015b244b095bc062ef3a6f8d1d40a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h360519d52e75797502475a9cfce3254ed06e75332ed5807eab4b948abbb99d270d06ae27bc99ac1cc99c693d4cae0e846b7443f4901e50238257dd519fa9ec15588a8d50e4909099a51671a04477137d051a210e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb91533c6b15f9b859570683564c48edcd90a22d732e1fbc8d87274e3aeee4860d57df7914033dcb470fe70ed45fbaaabdfe47588a3a833f3e7640d8432ad46205578c7e5ec0d8736f1af35223d3a7b09b23a6fa83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h384dec577fbf9b858b94b8a90c87d9f767c085f3577ce7a27e4e8e4f6e03d479a4394c84d648db9e9c808d248a4ec9195071195764533dae4d7f0485953cbe676e57136d6fec0836a7884d7153f9669e0ade816ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d1650ffd24b0a94642aa208d13a4de4a953b3db8b97ceb560755f802aa5172c4c032459eb3c30f18022365dfa4f43c838f55c4f59fe6ffb8d682424b9ec9f84348ce52f943367babc8c5533332fdeb60c4e4cf7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37aee1849e2311f883758bdafc2a9d3e12b2d693d49195dad0530afa4ddf2d3fe4d4ad7dbc2307ffa91893e3eb01a78042eca5b0bd372bf5ff628085b7f4461c072a99d1616b591b2bce87c82aa8a6a05da4fe93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36202b4e0f47f9c9100ee053b9594abc5035af3e4f69323a51da34947bcd5797804cac246e186555d9516634051f28bebd359033d4b06c9604eb35abb6361ff26ba4196677d226e88c85c0c054c8ba682a08a842b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cef340a1c81792c6cf440949ea997ce384b77869ab043206e43fd0673813413100f8b790e518d60324c3ecbe4d4a6b2403177b1178fe90f5fa5f9d192635e0d4b661b1c398818707da1c284ec4b745ee53621c28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa792b00028578855832770848a0d9d977a558ddd05f19294992f365a5dbee6b0b46fddfa7b701c991a6a38c78dd365f9c35b18635ceca94233026fb3960b3e4b7987b0b7364309bc279dbedbcc5696b05e390fbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6799d83c899575496bda89af5f1abc77fbce3f4de8530fdceea027cb84033261ecf676e807bca6cad298b4a5fed7dedc1d948671ef4e3a83e34dc65e8595c5d901f800fd2aadfcd1beb66045d16a5a6d222eeb12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97f3f4924e1f6e2a892f5f20dabfb383ca9b41c0467b855c64f91e8cc008ffe8a51886d668abc0788ea6201d4fd31b25c1bcc6e51cab43c5b24d077ed24b242258716f64aca656e5221fa6c815734c1b04dc8c5ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hceb009b3a201ceaa0cfe915ff7d1b7584f4da5bafbf8e86f1c24dc52a8caafbb487c6069104676e697f57fc95c99a71af61f1c01d6e99c69171e9d17fa13e1497b93ce8c4258c4e5f33ec4d77e57c1b31381b2931;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb35384c30c200b148b048472497f5dc5a0dab1cd1e8c1f059ae48dc06074f56a606f047854a4646081500561c87a9f69893d99fd8cc9dff9ad7b1b0aaed0bf0420650556342b4fc2d48d255c8b40db8dcc762ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e88deec1f02e6cc1bdb17a8c028c7e8bf058313561dc0cee5a8e58c86c24a20e93b6b54797267dbd7333452c4e0457ad7794f3d5527be59dbbe40b3d028e5e05a5b2e04295070384e2be8e9dafa9170ae9648eec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7920401e3731536b1ff2edef0f197c1f278911682c05a75f8d3568b433e1d8efdfd33773cfd7bda43d4d79012284109c8531287f674b9c9f4f8bc2fb353c50b2aa0863eb29f10dac8594a5cbd0fbf009fa279eb4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f0e4ed489615cf1e258a7195a0c3a62720c21884f166fa651371f7f0fbdc60d7701e42fed32d3111d9f29773c9b3726eef67acf389191292fcf10026c9e122f9dede3b60839312bd84fdad4446a05b0de3bc92d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66c14ec58630e7bf7daee6c674c2390edaa20c9dfcabad95fee8a6b41a72a935d545af18cd169c0dda425d1914106ad1e59a1f30d01c87ccf1bb473c1c27ad7b3ad11db47d5898ef7c87e164e52d3bdc4411a5f57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb6e9ffab893d33fab91a6f25da010d2318803ad0d729d7d35808e991f34a9a9ed3baf9acc2d50df89cf84f4a576b46150525a8e2de996ef15474fe7350480281ddb93f1a9194e081168014dfa604978ab5c4c289;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37aee691ec379b0ca85337d0c4140900add8fbebc0fc3f1eb1a1972e268504833567bd532a001d7bedd181a3b86e153179fc9d1a13eabef6bde68df54496078d356a4f86a8a9d006adfffd68500aa62112939a450;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a5c7d6b2df575d8478a7f150238a580b120eab8a99ae0388dd46856b31e9d3060ccb59cd67d4cbb4a569901ad5c49125ca074d456d35432d4038b67f9fc95eb66b5f83bb3fcf7ce7b560efa0c3962476326c10bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b8ad159ff8098f3d7f37b03f9bcb6f4540a0c02c70f08344afe12cb0b8030f6143d0829150f0181dac0881aa49bf4c83629231219bc8252edd8cb187191a9293ade446ab3d080201a0e92cb4fe9de41d9c4062fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95f4921f1c1632e9f66471d17662380b3ea39354b6e9acfd3a2cba2a40a7dd8fcab4619c7e0d999d54b3ae4ebbe3866a80a08bdaea2f894765548d38ae39479d11779fc56c5413fff7822e9795ce8b28042d3df2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h115f6b2608f59a9eef4aae6927294365060345f991b3b477813c36b51955cbb68d7052c8d4aab00d0347b1c3e688b5bf34978df365cf44dcc68a66a0fe2b9a3bb7dbbc89c3eef3b51763c3fbdd073a8a9205e2438;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79aebe628d4643ac4fef1feb29af9274054b61670aa682c543912480681077c00fa6b33c7bacc23ef20abc674d1450ac41cdf6ff852f96de653cbad444a988d0b3acc8c8ca563f7d0513e13e8e32be19622708f77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1ac46a27fc9fc032877a1a713750f6e734117f70e009594353abef11c3826bc9b474bb6224602ec889328ab29833fd1ec3af24416f54191cdfb2f451eeb3d4d48144194d269fd31144cff10b78b4bd23136e110e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h306f374408a0c25fa004390a1e391d89570b1d7e5836bc75a0738609a6e0bd82306927a54639801d48590c4b9eb766bc0ed5e89d9630bc1eb61dbe217381d00d83cfede2bed199620cbdb4e7edad722ae665f3364;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he40102e27ac17324170bec3d1712d54afd34548d5babfa6c726cdc76dc3276dd2e65d2dd01f21c86659e7055c13b3abc941530f776851149f3235b644c5d08f93ef8cb32436fedf2ac916ae7dcd14f1138e3fec88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb3b004eb14d536ecd3c234d3c7ee8fd6fadcf748a9bbc6b7faa7414db08c07ec2b432031cf32c43174764b4612d70ae542a1ec140058a9803b91bb63ea2ebf1da90f4cae7839ddd07b2e3e11c46cc8e3f7c312d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5518f89bfbbf14befcd1f149b11bad775d96629a06c68f6bfd1d9f27b2de6dfb542a9eb646d208f24d82b29b5759399983fc9a356b32eed789c20301eb5e5e5ba939a18450cb7e7ed398fe65aa121d0a342d0d86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6305f075b6ab79ea60b5d67517c4f9ea18cc2264ee6b68b15161b096c8ba158b5d25cea84d4ba020c1aa2b5f9891ac5fac84f0f307ae349fd505d7cfdb51c539ca13f44452a43efc443186a555e5b8c76e84763cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h570e4790dac05ad4ebcc787e62ed64becf0828a3a471064940e3ab265c9da9773778c6a53f99cf45308232aa8159fd02d8cbc490dc5ebc8abe917b20fa333335bf08c6d94212121625ce4677ed01d25c8a6944b43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48f782f01a465e58d644fcdca61767f41a2d686647b6db43b6c76caa8bda741e33269d445ce8746e7c2f38b4758b119421e9807058d6a74ade1b52b3a957d97500314c66b09a5c484a203fc417222afbcf8df13f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29671b140a752b043425e757ba56738f4826157e10c899eee583040044a5d8d2b8ac634e931bbc798ed03f269a066cc0e4bf592daf31a39605554baa39be94e95fd93d7e81ee2c4103f22ad1b89515919a7d37b70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5c0968e7664a88c30ef4f22e4ab413e5300cddbf9d1247d77846ae7d893537d6321d583066e1bf71a64cb105a053db18545841b45cde5ca2aec2266e0510d7a1035f183bca1d39937b31fec8c02a85fbd667c2fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c5f2cc5400a84f1b7044d7741e28c7684bd57a5b6b044aff39aefc16b006ba9c4d341c92d39104c3279118f7ba5705d90381cd85d57c3a976f9052d8d2fdbd17fba48297070f0cc661d2555dd0f6bedd186c5a4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf14325bc5f38aa74de1e8e9880b3eaa005b0af6c7b1cbb9364a48ef3ce62b897a5a0339bd66fc329e59df159edf1faec80ec3f8920b64de8db728150e3bc5bbf11dc23c5f01ad30640892f40280f879f2c2e020cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53d88044034f4420bbd84f391b45bbba34b514e1c4fcec9d5b7afa49d2621a6e765f24327c0a7361182ff5a246c8bf3f6aae8d4db23c2713ac554de7d221a4cde23fd362f7b6435a2176209f63e7feeaf08368373;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a6bba70ed34ecad81410f2ffcc1da1bed0d0870163d9c2c6737b6165742b58cdfd2a3110d41b65b2df3cef62b017c58491370e8f2e30e73e30afdbcdaae830a5c6fdf723d4d2760ecaa48445b0520bb2f72016f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a4273c93de7a7e637214de67e9384d42afdf173c1c19c8268e240856a0a0eb46a752cc8a7cbf4edc2c81b2c790f819b99346405e1818246bb1f2a3e8bcee199656d2742acb88be5719883b79eeb6f329c52901b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95f7c1d64feb2aea20427c56effc76b232c5cc6278c3942806bce34f1ffb7c99b0df343711c810fae8555e639a11fb173a0fba0d855c6dc5c7b6a66dafb4b79cc7189dc7a060318b92f29d7cdd167858b9555f21a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4d481ecec96ba84812e771c4c6f7425a32776b1b2bb722482d4c8e7d0bac12ce168a01edbb1fd05d8759dd1476dc3be742d426254a05502932bcabf7827d7fcf082cd8e2b4b40766c450ff62c8bc325393f77c72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha57b3c130e8fbf24b0569b167f70642f966e4a9052967a2042aa00bb02359d00354fe3b346170e7605571d8cf7f3434add2cb31d786f7be2dd3ce828b66f569882d9aadec40dfce73a4097a75c1dffebf5050a081;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd887b2d4241ed08062ed98ccd0bbb35577b67dc9ff0fb83f4b3abd590943948dfb4d1a3497699700e5db7344ecc52a9169857a2517042d365022d58480e6a1528262138d222544796a113df70c3b2de4ffbfd501;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h451e41a3ab9e0ab07f6c3c483ab286652cb2382f4dad45101c97a22e37daa5eb60953c7b552eadc9a24d2740780dd60d280d1839d2224b4672ab55a7948825806b693a41071c5c5338c67814e3235e40e73ce4b05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heac2e97cb78a176439b20aee133ff53756703eb364612544b67d4934b50209ff3f0e6fc6aaa86fba9703e44a6e1337cec71aba46343ce00c76012667f0fd2c0d2b7e917504c71120bfc67fa2957c73687852a380f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97942ff78e5a01fec4cb11ebb0839d69ef777a6f2eb0ca8ad38da690084da9a2885ee2822a83359f5fa24d9959aa5208d603590a57b1fb4fd3e926945b53e1925a8312f29b1d1ad43d14bfa26948f8a1eb07aa662;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb61e3ddcce58efbff48efa7e61af67d81d72816db4468712484ad40ae789467c9e5a26334ecba9e2dc24620f4c212e560410878b73fe1050d96007d4409eebf8472d383a7cdeea016e3680ff32fce7a4916990941;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b7a7c1d1215ff717aabfdc7f5a42698150996f14c09f0bce71bb9ad61b4a482df6b123996b71ae2a1191cf661c4b4443bd0a0482c08fdc25162aa19ddff4b8524fa8ebc9d3235399528b3be86c9ddd99f5a7a66f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0f9c969028ccbb709dbaa89d2edf70933c8bc93fe5908e9161d6408cbe4e9802bd1e66de5992245761f9fa5d54d73a7593b166349d21efb073bccbac175c928d9eb4e829f4c99620f00218bca4530a18fc3c80ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e6ba7d0324bae899cfb41ed30af716a3224e51f857a2a796680bc263f68e0756436562537688430af0e30b7831ea2dbe7904b7b482349d4ec94b1ac7593b387ce722fa5ae7f7da7c194fb6b086bde9f7bb7283b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d646132f9fca76f5cc35078317c682eaa8fe3a2425707cb709613b24658e68a0641efffe40f0680d24bb180f82360df73172ef86acb2a882b356689ad5b672c6f9ef6ac502f64ae2630c3ba4c4c6a84763a87c03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aa2cf31417b7869f8acd26a1563eafb47ffc6febb514a2246cbf4ccad2b6ec32907b02e6b68fb048a1f7b3e75665e9deef1ec721bdbbd2c9b8372bccf9e4e4d592059019c2290fe16389ea4bd087078de34826a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50b251b2ffdbeba523d45b27e7f7044722715e7ef7f78cf3f04b550f9be2cc75cdfc5968737ebbc5fc6ba2688e97811752a47404cd4c297ca76041737e046d364cdb73f7b8b4b6f52cea768485dfa89abe8721c22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h983461dbfe742e530b91d2ee90367929f32f396942d8e93b285009d590a60b431cab3f0e2b01d8190e6eb9a9e201a760421f591280ea29485cb22a9749467e4ec8b6c690c219bf6b999d266f3759fc11a14f182c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97510977da59efeb902c9f26dcd1bb2a2f6483d19c27a8348b4712269217807232abf401fbe35d43518e007d9353ec109c790b4aa25add1dff64ab6003a962186437248dceb5800e2f1c125825cee2db876926c41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f5b0889fe60c7ebb43d96a35e0c0a6a23e731c58af63dfe73f2db966733f9b78b7432b697dd4fe5cfe58502e7f158b8aaeb535aa0e63ce7fa548f68c47564dbfbb50966ba53a5339bfc6b9306981d7d151aef41f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b769120abc45a3b1e23d03fd1226bd1fd4db645aa8bb1f09b4047da47954845dfc615d47624db07510e5b13a912cab138ff25d90fd6a4f6467ef8e9b63641848fb1472ec963020058d2b5e2dacc7e7700e7bac05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4428588c66da982a1634d1a1631070bc29db7ffc1a5140b1f77cfda28b190afe819dbd1c2a2274de2aac6ef94242e4f8e8e77f651fe2e6d3ad4193dfd6d533f3f9f46b167e3f432f712cc88f65e91aa4c341a43c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97edde2f2954a8e790dbbaef9a1cc7636d3c5b011767d8aa82eb0bf2833de98564aa8879fc0cc025590ccc3f25cad2163cc66f284d281680fd4a7221a9c437cae8004445e9f141ee8154aeabcc67165a30dac4f48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e5177cfe01428fbd39b92b15cb6583b50023e6d1aa69eaa5e309b34d32f68a09dc7769b9703d913104a6e3c7aaf0e1104065c047a05b43a69829ad39360d8d155e39c0413c5b6526788e490c00cdab2c741b1bf4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ea0afd5ddd5280dd7a8b35888343ff30548280111e202d95c58793b16efa2b60dff16fb50f39999428ed6471dacd6cf7daa0f08d0c58c8eb39dcd7aecd4aa9f49619cd1e6b9d7a059af836ad95f612e98611c546;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a1c9c6e7e8e40ba1a1dc60580efcd4c8b4ba79f6ef18eef57f44897f8943ba847e2ef408f62b6d9a0870ad8ad2c6dea45c49ad3600f72cfb81a5b01f4c39c55dedc2ad4039b92daf4ae5163a17bf0033da41e518;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc92cbd787df230f6c9e35ad9226d5722ec931ece029d85d00b2ab068811f6e4477958e8253d8af83afadc819a8a98d608010cd2501267e77b92e8842049a4425db84ce601c20ead73f9303428e82cbff10251dc4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3ce98322d478c22b552bcc6c235f1a99cd0373aeafecaa2d43c9b955586f1d629a2c2d327d98dcfb6cd39ca32424e80e3b931cef6efaedc775260ebf7c346b740484c8e2442c33a6cbcc548291932eb1e48d4114;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4c8a37bafa34963191720c35a4c2dd159b23b0a05096a92368b4200990c8f5d3e785cca03455594274446822927a709f12aaff6364c3f6ab03bb96e27c1fccc0eb10674c4ebae7ab89334e07ce643a352230169e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9702bdc702e2896769d6f56db928e5eb4a323c8c6af53bbf68112070c2b6792b6784ce0c43f818dcca49c15bb3653b8a00a47e36622df6c585b8d62a156c91357a5cea6ba8bc26b5c046ff5d92b3a98708ca2b327;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43799b4ac66b0eabc09f973cb9032e144f8ebff9701e83a1831fc03133e2d254571581863c845d8bf97e67e16db7385cd641dce9268c60cc085bb61610a39fba73b3d94014be11ce53448508a245f7c12ef835363;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61fac69ca19caaa542940e5dc414121e885fcfb7f900d58d36e8d4772449c7e9ba3d54e74ebaba367c154ad5e93c4a0fc8365daf23933bfac49dc9f6825c6772ee3ac7b63579635e5affe7d9298f8df14c22a1c9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2eeb8adf47c8582c682c749ddbf6be192cb5a999cbedc41d8e58fa15476471ee474627569fa749c6c66b7dd116980de4378f553fdfef6437f0a3dcf5bbb6414dc725906a95a2218edab76ff30206858d7b127848;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4d88b3d75413d0666be8a391e10deb83d4dadad510809855bcd53957802ce5ea63c5a557094b3ba8d65ae8df9616232a31977d0d51196e083a4d970892a1ef4c0a8ae8df4fe0e9a9854e97bec91023cc4624388e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97de148f6ed425cc1e641e46cba493acbde099305c603d53d4d42755d834dbae8441cb82f92506ed44572836f27ef5f2f2cdd27117fb321ad613eb807c722a7d91141d451b47ebdb2adf9062d77830f3d97a72ebc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d366ac9afe14d7e69111a5f20d471be070adc546f6c4c4e242b2b72dd69f046448bb2d497639ae35738f2cc4bbb8b6dfe557f618d9f477f4d5f0ca091af5cc385416a30f946536444fc6b32b98ae576f42c76068;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf32e59fb7616f771e35437129126702a3900db923e3207733e477f368ed7323ba47f63439236af6dbd06cf6e3438c44c08ee33ac5cea02e76e1a4279faa16e12913759fd0641122eafff802d9895813ed09adf4b0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h702b5374aca6d60e5efa710ef8f8427caec5931b513e4b386dbe6cdde255f0acbb23e243e5dff8fa44791ed7863ebd24231bd88b78cb762bc923b2a619d9e60c88dbe92d65a867535d4edde946d991eeee0b9c0f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf638749ba2cabf9d5cbafc4d1266b957a0cbd197d9d11caf5b04bd9a4464cadb2459e43215277764cf7594f8cfa69631a8269d231f17c70119dfd5fb85a4041975958848337bb8c04b700ab09e76738176f726e38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76262479e2f89c0d6d614b32394d379b6f05138979f65ded910e99e57a1dfa86ce9c1d39c168d8c373c64ba656fd9e96027d97ffac689fedb915f84280c36d78e0efec7194f32e36761ff76a8a66722ff8ce7c76b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c76a89460840dafaebdce302467b3b34dba09aecc288dbfcd78fff4fbefbcb1774a49f29fd73eaae4e18b502bb9f82632872a2df6f66a54226589cde7a261b37af4941864c0199b062aeecf98d723b112217c53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h997e394cabb3e4cf24e13c229a8a60b4e371edf7a279e881af05ba8b96584725a5dd9f9c00b2df94ff9803776f6fcc9e3bd8df5ecee54c2ea313fd9c4ce8ec0a15ed71201b7f6d938961540964e4f650d337b3d7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4da8df064a64d073051cda052ad6f62154940ec3f198d0420d71f261fe48ac678cc6e66856afc4ea13fe41525d9e0adca17a30881a82550696eec5864972d221f974dffc4792e82fdbc7bd029b09677532106e4c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he40db40d87c5bf4f726e5496d9643534ea6e91b45d3ddc75ce0e98b5587f2269dd104d512569dba4729115601118acf4e232c1ff496f589c5fd8285e7a9107ac804896df28e093f20faafd7538983eb94b01f58f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he68e52bdcaf94a31a34e4ae72d0c7c62b6b278dd3cbcae8e1fccab3f4da311501e73d156b37be9cd6d1bdd0aacf6b44bf2c4949995bf114136f9332351a51f805b96181934cbd4833506ebe80e515488158c5ec66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bc3f597b8ff7bcc09108447371cede1b3a11f198ee535420f2fa8fa2765a61b6e1064dffd0a49f9bdf5b5fa11ca7ba2e089652705e293778beb300827f1fae907a5e18d88e6f5ed41ba6971527e13972965a6a9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45c98b15cd4b6ab776e7d4f67b5421cc79fdbcdecbffc9392a19f1e774eade05af74bcab0742fc70b8c785a18d27e29bf5ff3efcc8948513c7980c3e48fa9718594f600964fde33b81b59d0ac7b7652dca363ee00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf25e75c378f66c25dd6f196b6bf625a4b8b11f38efa0d5ac91486dd6852c71db74dafab475af4ec1653e1fca70f4999c8db2b3a62019c74cb6adbc331e4e97efa7abf3c87fa9b8d648081e8c459d030fb3f3a886;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he60dfa54041c8deb38adfa6c2048cebaa81f8eeb6228b40a2411c327473f989c86de1a3bff80325371b109f50164fae7895ef601999e4dfd833c28a0cd8b60b47e50f9b82c5022f7701d301bfe18897789516f6a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d95df9171282038090cd1ece219830b98960892c06b3553c74a8049f4aca7f86f0718892246a3e4f7c2eff479b98abf3b0458c477b5f134da21e4843904e85f4391a426265f33a884cb0021bf61ce6408003fe36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h319ba86fa982b320db7a6ccb1d7daa9d739e262944cb2757b6c142e4db116a837d138809ca15f0eff9427132912eefd047e579f361bd5bf500c858bbe665a8b99e5c759ea5191e06d9ef147f08008d3d1fada7244;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8142ef88da6b70178a74af9df34f80d711cdf3c190ddc51bcb205d05a0114f193bf4c609a3438e564589b48837e585236b846228b329166cfc393445d472b085c452fd02626c81a40a881d6747de1d832e24629e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha52459770025f01bd715b596429891c4c97bf6d26db7ddc3f8cec8582fdf5325082519db4d919ce73d7ab63f84295dd2f9fa4cbcdff759937b21046617b20fa286e0ccd8dd3003eebd13423c9826ed65840e658fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44234a4c9178cbfbb799a23906917c6d81cc17f53a4835743f65a14bac203254793b2e4ab9fe56f339652a339dc9fc2e1585e2fd1ffc515a13f8a6841a97b3ee91e672c114547c78bfc13334dad123734c85635bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeea9e332467ddb0c7f65c17023e8f739bb65d40ab2316a247378fda01390778a4910fd1145c3d8122095615fe209924b0c2cfcdd93db940bf45d103ea18d00315a5ba5b6bfa79b7242a6e2958acdae500cf9ec73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c84a5dbc23c5f700b2c3b9aa9b6c683b48cd9c34ef6a5e1601f697c50815a473fa00b2bc0121fb2a5facf3438f1b630f413034ac2ea7863e95dbca5e929714bf37c4dd39af53a787020f93c2c56d2bbe900c6881;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11d781bb3de8d2e77b81f27710e0a390ab10c5d4624d8c2e9a975dac767a49b68fd4c66c503304eb27612226a1051932d2a909f2ab6dee31ff8cb63db4a5639f018da0620b3dae869650d00aa84b7e4e59409d0fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62ea535e34ad31970092fa9dc0b027b774f625924a501efe658e25da39c7ec418521a9369ce5b623aaa335dd3711d98c51bb18becf09a344db71d8496f3964e916d3fdc492cd55084dd79ce7e7cee2e0c46fcd4bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9c8e61fa93409bc89c073066609e17c4dabae9131cee950ca5ad1bd12c8c88f57de32dd2d730f1bb327c3995f0e3e8197aa780d496165f0b398060b229f0aac3a3961e4b57980975771fe99ec9b6c503381fece4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha638d7e22d857aabbe287e53be904159534a8379c1ab7407411f71f811b535e8014d65dc6f777949f358d1bc12c836066edf76d6031f5b18c224c7bf4729b92f3e53ba217ca3ee3cbb4338c4055e8750b2fa4bb26;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8e57205b99cadc36111bc76df0cba59954ae1372257fdda773cd241ace10d36e309d7983a9c875e65a65bb2db8489fa7c2cbf95e1a399d601322d28909875c3e7b8be81c088fab69e8b244da3a3dba8dea04af15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5e463137fca68f1b2c5515618ac7d0ec3e18f49f00b6ad779c35ff0b2ee76fa6dd2fe8204d273b3eb60426067d5f9e990e34eaf65e34ba18d48c125e8ac45ea9e4fff8a2006e0f04b0d1a5ad67177d1c9cdeecc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he10b69d1786f08015bcc140c0caa1107602fcb75d257880c5bc9551da7fede2573515ce9a80fecec2d2d761e4275831580ababf0d4d3f6b76cff7c3cc7b4c91e226bb55a788d91ede151a6679839603817d45d123;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d991d37bf1bf8cd9f635998d0dcf1e725444b5888fb941ed5a79673cf7712cdd2ac12ee17e1794da4839ca9916d5c53b92e6e822f39993b85fca772dbe49db4714c4e177556941d723efae10093799b5dba87b0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34531bfb88b3004370ca79d8d612b7202ded7fa5ab43559c77c16cb4f698b98c1671fec00248801f2cfcb01ad45d8f4d44c3c3d2fdc0cd27340f6d59127dbbb867c1fecda95818fdf1b5debc833d5d1e53690abfe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9406cd2f829d6dcb67681d851019415c77fecbfc29c9968f14227c4a593f47984f26a91bc7c8d8afb266c728569c41955970e702020bc13a3accfc1d4af896eb27541b0f3b9dd75707cb18f3fc90659642951bd9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9497df16f90b9cad3bee33e256bc3f79a07c0e3d4b6dea3886dd326a76c1e0acb52bd4d5ed5a499f4b39446b44a54123a70b970c1f61fc531b84ff844db0affb81fca50dea9e88ceb49ea8105910309f1c1a36e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48bab24caae401dc0ef97fb09116cf90861ceae77607a28f69152ae8f6945ad86b60dec8788aaeaaef747821d358b02d342644b73426f8509d94f9e23ba27f9b8d6c6835125919ad9f5fdc4094f1368d8b78130f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe2115e4d38133651b2ed0d3415b8bc4a870b68c9adea8b16e21f8082920a0f287072d3c747771191efef280d7cd175d0241967a5e83eb3b4cd88b0a2efcc6b8f6a2f1e4a0ace1ffcaf66969cb7b1576664008333;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf6d26e9d9944fb75578105e1f920c608d657536e2117360cfb137b4d75a8b16fa8707e321025cd21bc40d3898807e81e08ead5f156eb80220e61dcf9e8bfedf0b31e8e6df9c4b8d9796bd857979920b2519ca0cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h262108b9c0bb031332679447ef54aa02c0d3da6e102f1815185f121decb6032baa01735079c227cba7a648627c6108839c949bb4167483362aea67ed5a67af530e4098e334f592007d83285768b565e5670873521;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48649b9d66d5c368cbce49cda7d37936b732f31ba5b8288b73c4212a641283fa37cc52cac25e70393aa0d738b6eeeb751b92d556043331ab80659e122ffe24f56733cb67d9800f0c6c4b878d14c743bfce8681a23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf123c960fe0e7c75b482e9666d8c6535fe5dc62f9d267d47416ca0eb1fbe7fd4adb3e94d9f20481ac9268007790de18d49f415122619bcbf2d49c16600e4994dcdb6a063317b45ed9632c7966354931e5698dc1b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78f2c073427d1bb9d24ae7a6e8de7aad673d7b6e20fe84217be60a4798f15583b68fe69b10538228d056556ccb4812856aa4608139344e1402d1cf67dc193241f488f8d1dfae9b66786ef49600894c30d6a9ed476;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb458cc5cccf26538b3bf6e722838bfc2648afdebef1ad94d461686eb860f80be554912493d988d2efdf1062bdb136bd9f7000b067d3617ff7b60696bd2a381ff7cc5ae93e7b741bbead34366cbe75c57a5d6e6d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf92d24503941701fb0ef6509418215020a647b18e813ea069b6c36fb7ba888ef15c2945d4b49f2b68d3e54090646fffef149382f007d0a890eb9be0598f9312c83da67cbe30cf10f0e855a0db618d3456bbc8b6fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56d67532911d5ee5f1a181955cf8feca4a731f37a74b8ae280f96df4412cdb055bc042df3e053d07787e8a7b5ace43c23c1ea03cef03790f6ab7b35516dcc4573a101b1465d6d38710a50d9b94f33ebc05598040d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61be20cda89682b6ff976b318225880944e7a352c8bc29e5bfca9c20642663808b79faad8c3f0acbb7fac49097d7238f7089d941831a99012fde655c71ad5beca9a43c215e117c0c08ca6e48349622f553f7f9e38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5807e8fc4dec419722da3126c49ee75792e194daa87b9f9e35f2baeba40c44d95a10c6cf99467f190a4efc5d55d4249ad66482bd328a73033f0ca7faa5fe9368863c1815951e32ae6fdca7fdd2aee98ac2bbbce60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h210477d1440b30ec068634bc65115a5e2441a150f2977d53e1585d5643600f9cac72246ab19d0bb650933b6b18eecac4573511e496234a74069e5481211676aa070cbd841667a0cf531d014d6235fd3fd73203dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38b581932d53ad4d1ebdd91b5d87a1e89bc1042046f6fd550d7f0473d199567105a19b69ad24b3b72b72a061d592d348ef74e0137a6c7285e1f7251217325e33801510c55e9d62c00b8e5cd5e1ca3d91ed8ee9985;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e25f0a90be6c2d4f22e32f179f58940421deaaa81bb38270deb6112872b1764da04bd9aceedbf82719744eab671d23b84cf42b9b05f3069b11a530437267359f4de18e3d85d9cdd8c8aa91e1e7ec491d6b49d1ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4738943311c6976fb0247e50bb992028a2e9eecc3cbaf4ab8f9480ce62d6b235dc0573645258b417b1be5952877ba1802eea3d10f373e3b35e74c36a333533a27d223b7c661fcc5fa306cb96745d020d47f66bd83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafe797ff7a32da133a58accadbbfa517d043815f21c83e4a81c46a2be288a9295bf227f25183fad1c415a2b67d2cc9d0201fb93e0574508b9c7353a559b8e272dce16520a265708631f5df16aa8fbaa6bc9750d64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h717344f58d7fd7ec8708ac8e4e4cc03479ca4c9494ebcf27e6d562e384a486da149bf142793b4725666a3b509e1e11f64818398c83d7e2437f275d6c0a1e03d1a05d6fe8fef7cd0e0e1a4528e1a00b0e178e4ec80;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36ee5dce08ddc6e0ab7f191c9fa64ebba1570e01d419cf7733e2678e0adebb5b8fdf10fd98009c072ad3d9a7b8f76cf044ef68d9a4093e8f63286d7368bb67e8413d7619c29c46393cf32ff5660d9d7cb860f1cae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0f37c94387d35f77c58ef100cf915f7e2d1fd994c361c552cfae57e2331eee3022660ce581198b364c294bb038077ca1237c30c992cde1e40b22df9e9a7954674d0c7fade80ef77f0b097f1af5189192a38f8a05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3024354d6ad53f25f0476be1043f44aa30b100b69a214814eca837f3f38ffcf732ebc7e93a72f7293c79f54126cb3bd0053297b58a15c74d84f4b80332f30921035ebfff326004bea4517ec01788fb8fafc99250d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19ce4a43247d1513370ae2cfa1bd385d7e394c6f9bbd6eb522fb12b7aaf448e26a18f2ddfc01da9541ffdc631ace3a5bea924756a70869f88e1c5bed4e7fc283039a8a2ed6037ba72d66b0e1fdff0d9213a9a544e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb840133b10031a5397ae2eaff6bfe8c76699826a85130ab13e92c642f2625888932b56ac5d96b7e62428b49df910dfe1eb42fce764b0fb448d967345da93ab20c73acc39fa96f9084203aeac1eea0fd3dd50b0360;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b0d9cf17215eef4502672f30e75d4e26e7d0d512a3178487a207ceba201973aefc63369b5facc3503d7e3b8219f2eb38223e8a6b0e1446bd3d4e49a1e4a2fb59850ff1752ebbecccaf5c4b58c26f5328a029b221;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4804e04dfa8a5a5ea5cfa5463c27227c5bfc62ba075a3f79656b0c02c3f111e55ec8e3b5166b1e0a9c2e2128f7c9b5bf57e0b27071987ad2db0f91e5bc4e301e27e085f8719e15c8b2ad73d06035bf134a1ce9bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1d6d10ff9647c49486582609139b9465b8e7c2ebd6ed72b9971326750f2e4bc652d37bf416ec4a10b2efbb665fbc6028da87cb5ed994ea4adf9e4b822f82443625fd61f338c376549acad4261db33612d8d17943;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb01eb36084e8cd68f76378a5158c55eb493ce5cc700b3159092ab1df7beac94ef3bc47896bab362f3aa14181f30438507f6f1334312a8da8ebf8945a9d4ff8ac68d82971cede84bb27f5edb0ca971a61836e19dec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha10b1577b798053baef10f71a25dbd3b8ddbd8bb52d3750f8a60ee16640a7f8a97431be6372221c4db88b7dff4eef47cdcbc1257eaa00c5e1251eceb889b02f68000057ef9a7bba538f8ff606ab28fe7ca0d68b66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h896ea429687519054c7202b704e11c8ac903986d00fbb0a5e63ba6dc93f90cb21e10b793aba766dc51927814fef4446b621d084dc9c8e8397e505a042403c72d3a7b22dd9e675b82a1691ca2a115cea0282179c9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha617b5e5a1866eb15cd41b3bb877892f7b04a38d0e56c12a2e7cca5ae949b6d8451082a8d70d4e8f8b7c3509a09f7e867984de0818191dfb0244a1c6e5bb9988f77bf903733d9ef5787a8178e3b87a16594b4ce8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h209b09364f510203a997fc4cdc8a2aded3ecb5bb30e8bd3492562a8a600e4cfab0db8af9a9c8bde1d6de889eebe3e135c8a154e9fdbe244a02531434926c132834041ad42bc5b91a700ff1d7fb343121729e3d7dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dd5f4463d0a6fef78b827159187b0d75121b930c356bc00d348bc921b9ed0fb552f11a4f93356c87b360b997fc8258cd60f588b927799edd9374b64ade3228ac490d0be5007d16f3e9b0e86484512203981bcfcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab56db6b4724ba82386076057d4ef4ce94aaf57345583b989ee8eeca9e7fc4e9688f842d895ad3bfebc6c6c94d22087eaf8e8f270463d22edbd6829e53d407c846a71a2cc42dea43c5501ce1fc44e2ed23310733b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4788460762679b07017150c512a0fc0e5bdc24b5e79bd9fcee931efd0bab787119c5e81f05af7cf43bc49e6ace32e045025320154a5b504b36326615c8b78a1207cf83ee1bd2926920980098759fcea0b9c42d5d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7840e04ed72643711d3f43d65704902aece41d3ca639548c7e44107e91d418c78e95d1549d2f64eb6260794f23b7600b027c150d85d26fa5d0535ec36e1c9741e3b24d3f21719a8de1247711fffe5170bfcd47005;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3f65b3658ce3f71f0318335f776d566fdd9deaff354661638a09894c659712f3c1c487ae00ee6ea5024d8bbac10cfee875c3f2d61b81074dff12d6c6ccb1d1c07ac066656c9c52d84009db4780303f1f8d5a9f66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b43fc46bfa7721a300f0567cef452f382c36fedda07d1edd4fa5d6edd6e7e0b8d350f38f549e9212245cf6dd645a2b6b0488e8df6104fce5f3ae6784e595860d7783356762906c7b0698b194183578be79924666;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51509f43ba2afdb699e0b1e8aea28725c6342a87560bb2030e900449639ea1de22b6ffe77a5cb4716a49850bb593734e873e1b500afe9f4506208f7d1a0ef10eff33fe194c0e72e513ebb34664c3db8845ee0787c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d518da81021e5807046057f6667d6b56868ef5d8273b83af58f3d4afb2878523ce46461342d6e1c39f41b37d78e8115fd32edb15c4cadbd71ba81db217cdd79b613e92b5febe3a1413d3e783554fe482176a1d7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb83f5de07304e4d71655585da00b23bfc1da1697428c1ae0517224019d4d7003416047e2381c835bef212a234b31594faed8835de4869f7fa2a91cf7a3561465c3cb07da8d4e3d72f5cec312847756958394a8f1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h393adaffd8e863f4aaec5ed339f8f7d3452ad026ee3e68ee8e4ceeb1b38bfb266ef5950d205be9e497fec9eab13cdaf1175756444ed1f14e69b660dbf39f5df0bd51e27cca3d90ea293774b33e73242df98ef3dd4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80217afb228f75c931ae91764a1d9c8d6ce6d3d3fcfde6646167c58ccea65e0cfbe9e54d7d87e737168fbea9f5a0b6d077814ea5987d1b3b6ee764276f1a9ed8e0767c8f3b1d67214ffa3c6cef67b5233e156b140;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b78af0e907c84535124bfea0d297bcf381847b470ead54f2da664633fae48c2158fb117bef9efd6cb88bc2c9d39036f2625c7cea7954072db299f58496b5242abaecaabb5ce5ac14bd010e0e550dc891750676d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9078f2b8c98630b097e99f07e68ae2a21603a3e887a3b23a6dbe1a6119e6b2985b45bdac8ca478ce7687d7ad1b6dba2609571461976ee7e35e974d8df455be8724de93aa7fbe0ca4fecaae8e8d48bfd7ef7b7d7a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda23eaa0724a3043cd337050987f37833ebf85880b04cb20a65a49107811ae26b69d46057ef5aff2ba76100f35d6b67b1127c53e9a696c8fb305d750e514228693fea592b9d8256a6bd5156246d573a9e8fcba53a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaa534453cf1174ec7602319607f585919519de65095dcd6f0d3dcb64045d583f28edb7065f8e428c5c958f9a50fd6256a800b788b1d344c288de7609bdfe9a853f639011d0f38faab30a30b0feb8caf380b4e169;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27b14719667d9a55de2b70ac7b3005650b500c80efe4f7590a98310e4abe0a94342af0f829e5194f6b4bc9fb41ccde4f276a50eb5d6802358194e3eae614644f8fcb5823b9049bd2749a69c3b7f802ba7ab83d6f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc19b68e2540472f0e9c2f011a563560ecd3dd05c4d231f8dc00b066cdce564a394471bd812ad16ae95be8fb71c0ef6b2b927bfe2b0c7666d38e95ded7f155a81cc5c11148a6ba4c1ee8afdc0cc407b6f2a56c5a6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84d04ae1a75ef53f8c00a0bd616adf8d8442e21c58a217e661cb1d745dcfe1a3096b52be6f7f12b9cab9d33cc08df440f3c3d2722fb8f3ff56bcb2b47eda6d86ba5151eb1a456e45490532b67675d151b44026de4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdff9c555d93b4e0e361136b1cd34e308f936c3f8e147e7264ff1e555aaa5c3e77a37f3b4d3d88df3134459a1f2768864e6fa037fa22bc2e9f2ba4d6adfc82312678bb5e1666ca586d3512567ad0b3c64b7767336d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeeb9b4f6016c295fb551d6014c87ec2faab3dbec9ae253b4bb425ecd8e203a1afa4367d43d8ecbfd223676c5fddfad9877f0090dabf1cdbcf2ea8d3a4443bf4dc37af010a3167c51239f949a9f035a0916e53d8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23a53a17522eaa1ce382464c6a58dac8f2a51e26d310526827dbfac2d343f777ffd1d7f5dfd93f3d8a47bcfecd6bea13bce945222ab0f3fa02f7cdaac94a53656138a4e8e4f59204646927a747a13ff7cab0e9cb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96d0a95c1c8b2f01d0ea1cb926b0127468748bbae95b0fe4866abe2ddc7a0dcc359e1e89d319f0fbf575d41b6abef727d67443fb6eef5dbd0921192012301dbfdeea36a944e272b80ff8877c6e847dc343041decf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a0d33ebdb81dc0e6a8c4242dc17cd80ad0bef4456c467f3fa7cccbd3386a29daab7d4e6b5e31903fce847c97c878a0de45c027d0e150f71891d931610471eb51f687f39ed19cf312439fb39975fc918e411d623e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8abc7e71cd8bac0f252d0849b6fdee0237b17ee6e9e2bff503b88071e93d855618a1492b16e8042656b09316f45ab7b36a3abd6f82d327de914819f9b8c93f198fc368d499c4add37bd3614705452a193e2b79a1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0127df223e3bdfcb244020dddaf65cd2b659969d6dff42f1c64ff237931855e4683bb4f896ce47997f6a1a963f22ccec36727ffbbd96a99f168815b7be724281fa581e12868864faa2fdb00b6a9e0306fcd7b76b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78d4c6d0855f1552fa45105ac9d907a7d0d44c2dc806351f3c892787dfbc89b71830cd6c82e9c7233183e111b7927898e974479e06bfe9ed559f0c405cd279f9b788772178acdd1c089901261892499380482d6df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef2f3cf3d4b50ff3249e62af3b8894f07ad4f623cc880d976aee8ec1cd5efd619c00a9375c5c9d0fb7c990a4547415400286abfe442c20580f3f6470eb9300422155dca223263a946343a1f366540e6eef58bf3a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae720cebb0b66a342edd9f7f2b3a4e44dfdd641ca4604c4f7a5ecbc536ab7f23281348714828f73784458c99413259c88544b1fde53b7cc1f9348b199efbb77d68c29ade7418ef55d7b721c7e88c0d71eaa91e063;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72a399b29c00f827a14781b7ef02691a6e7fd2421841797a84f4b59d4544e3a511c588584dfc3eab7ec9b09a080e5e13edf0fe8b0267bb517d6d623346646549a81a3ce26a89e856d2b081ed14d2545a8e777d4aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc098eb9aa8160abc990efa38b4feedd35a2595f4a0848f0d80f5732b2872f181f42c074d152fd86515cba2e8d5fe16dd8a305878404e10cd5abbcbda582ccd4b03e137f9d4e4c56c91b6785d3b865aa020adad8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34a4b0920c39171c2a5c04c220d80c9cbf511bc4a836814277ac648ebd09f49f520cb635896568d32293117ea6889c0a01f3975cdb9d47eea22fca92060e8a83a34ac233bb019faa5a1ae8bb5910640b35455be40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b82bfd262e3b129d4ba936b9cdf6d264874698a0a17fe76e659c5a9631571c937551414865700a6b429696546d9dade3689c61a91f7588f15a09e16b6876d4fcd878003c1a03401e7b93aff9ee57fb4c223c79a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0c0ae28548f6ae1d53a0c58e4dd74345e9b483df73c954f9bb1e415f533d41eb7e049bb5e4c71f65a1ece1bbf1ebafb646a42ea263e26908217f3a1223a048cb321ba25c1e8fd354ad89369f87f293c29688c03c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31991d3f46ee425c970ba1c62da0122f9a45486f02f8d572023f46a70c4658452dbbb97f9091e64750b08557a94a2f628cf71d9e43882786d77c85f84355feaa1cc0243728ef5fc74d1416c7d810d0cc1486da6b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d9953b8cd9fbb615e31f9173f8b29c2efa3cce95391ebc9b5cbe5242fda6e4e75d10bb3c0badd8126fe394368f30501e0534f825aaafd808c466b4a0b6fc44b4718bec7ca8d8592618bde6cf9a929de654c0e7f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb55133f403f1d46be4265cd5aaa9c517b4a15e8916307765e1983f901116bcffd7d0b2b3891f4ad99ebdc27ef42a583c1e1993c7a91d2ba3b78833b17b30567705c04ee821839c2b7c59b4b8b92bfd63deee57543;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd3379be3885dac19c3c88fe61b0b70f6d0cf6cf735df4ab110c6241df4407f81fb6b397ee95800fbaf9260620f2e44fdac8cf51a9c09617e8d87d35c2635921846fc732ff41a4fd40847599719eea1aeab9a798f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6886bb20f164d9050bba16110b59a6e6c3f5d221d36f1370a8948a6fba47a89dccec17fa6a9b4761f6cf6b04dfce7942d45e4e033445c16c332919a119899dd1acbd64e9bb9e7b1c9a0447ea99cee69593e6197c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce3978d4a5a6ba2a007bdd2b2c2415b76f9a091d4f7f65386e4b4a6a6550f223722a37e3742642507048fc7bb7c7e701e45c813c706cf36ea31c616bfe41beb4d99e056ed33169dfd71b59e9da89adf4e4a0d02f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba4e842f54db37c7ea982a44e7f771017953bd55a2b01f3ead6d04ab586882dfa66c40c64337537d631042837b8ffeb137bda24c469ff0bdc2251f151daeb93760fbb39f5907ba71231c849d5df32c934db72e2fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95cce01be7ecc01d363ba019dce9115fda311d9aabcb824a1709f3cfcb12e436abc9f990062846919cdb1e969ae5c206c30099cec78506bfd7b59b94bda29143aa5c00663bc9f84bc7001dcc72dab6a5930dec36f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5178fb3f2532cf93fa474a5826258d1981054f493b906bd7f2c7720748570d47acd91fd2bc8cdddfc603ca26fada6d8a4531058008616d089f9e08e264e37818b58f7732f6897d9aa66887033fcff7d710b64393;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h478bebc90252d4eaee5790f4adfd249556310459da2b83ae347ac7226e15b52d0cfd0c061c55da4dec24f4e292cf5192bb580640fcf2127d8b5ec049caa70d2a8eef5b3809d15e88df54d0bddab01e24bfb78677a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf89fd9c480b909f153210290bcd5e9cf5df43d2a928d4690dbe3ef2824cd41cff0e75409a16367d830d541e90903af78374cf081d7a2f387495e6667b87d9ec52fc5d11fde3c0c6f44437aa3c43be22b7d7f9732;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb87bb0a0185bf1a7b991d2e4fe6dace09e5e33b7d2e5add3b44c104ffa69cf172210ffc3cbf84026e586d0bbeb3404473250a6ea3eb490636852306f3eb362bcb4869b7ec6e9f436fc8ddbb635d4b14bea873c2bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1c064646e8fb9552b17c933f14b7eb2b5b8036bd04018277dd2d006eaacb0a608dba21a98dc46b644fcd88709320505a6f199891c72d97ffb4e8f82a4c3d3d94c8b1d8fb188e62677923f605a7b80b682dc416ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda67cff5d86203ca1e2612d7b717e99623f1c2b37ad2ce7e280c9db4d31450878f08061a0e923d3830cecfb261eeaaffafe837ff6a15e63901e18d81c6ef9bcd23509a677f8d149cb8f5120e438b055706d611cfa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d1907fe32c2c874b0397897fc9e3ec3eb4fcfbd8b5c801c91bd5a89789f0ac388787394157e2130f5d7aeea0c2953565f22ae5944ce5df64f9175537d72d25e3b923ce4f36836479f686567108a044094663e36d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had5b0086906a9248dd848150295329fef5d27adcbf3e2b4ae69c73bf0bbe7d5108369f7bb2fb6e5295c9579e9ef7daf76e874d21bbfb76a63b98c7d3920f2f602577f46f6c7ae85ef3024f3ab24cd97110ed0f873;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2566567afb13b6ddc7976cd314fc425f33a81fb15b7f8155a578465a2d103fc98a775a8d3bfd35f9ce8960c473e9ea01f18f23d7e27ee65d9539b07a1d525ebff1c00f8d520247e20afdada1f6272504f94af9aea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f6649d50f99c984040c230683d219e1c1a9f88ebd2cfce021ff2a476cb5ac102646bd94f6ef88ab8daa13ae423dc4fadb6ba5c73de27b6e8ed009102106a97a619f41788b4d02a13c4323efc69947765a7896a23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e37149b8d6a5d986c3b114aa3ec548c927caf87966252e3fe23969b39bda1abb40a82be799490e857c9751aa85c958e798e6a7a47762b71aa46d016271626fab2cb2c1753d606305d6942569fd28bcd682aadce8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8096b7cfaba673f4b8925bdb4b69f87b236ae23d3a550f6b053e290cae578f3b408c1300e0fb22dae4394263a1420419ef3868b85a702a643bc75d751e01ae91bbabc2f168ce6b03babb79fbcccec750e11cf35e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53e898515f60d5f46929f532bd5f23c6a2fc956e0c0974a6ef67244873fce3311a55789b53c64c17760eec3db2f1fb395794c8a1447ebff76cc517b308271307d55fc4eceb576e0d3dcb0cd3a66646d4c202daad8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff6f4cefe40643928391d2ea320cf3bd879745274848436774e2485d0fb16def5f449497ce45b0a2a0c8722959c713ae119f2f4646d193ba51fea40fa4a550853cd8f9f3782a08eeecc3cbe3c6ba93405e12ad0d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b4960f72bcceb12e0b94eca95b92a5960fe7978dc7eb6fea60687fe9d31475a5d40e19fa07e408b6f983b9a56c6701b6f0ac728a92e098f94bf8a016464b4ab533278c31d13b850726e5b5fb18ca2cab2d402d00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h505eea942474a3357cbc8a56a2e4b34483a4231a2e2e7fe9768fd00f798def36adbc18d917838c66ca0de288f6dd4edc064df6e55693789ab35a52ac16d576d0e51e4f7d9068b3838c0223cb1977cd77616e45f8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf7844a06b8983cc0225261aa9da0a89992754f5cde45aca28fc8ddbe546a222ecfee44c567a3a83a9dfac74f19db1d6a40cc58cda8f798d670c2e975193aa7a19f0b2120d126dbcd2854d22516578adaf3f07256;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85dec079b009072097b6556a035a64dcd8803d71b6b4ded4e9bbe1508e4e1fa783ffdf99a8582cf674674eb7a4b1102af92ce9a26c869bcbcafff791f9111d981dfe9a76e9cee83ebc6cd8885813465da0be1dd1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he649609d681d55240c7737711ee41bcb272b51344a583457849bbeb94a19bf5f878ede45150fb5fabb9c4daadb83bafbaf81354df88cc17178077b1d5d13371815c375296d1a0551952ac87fafaaba2a0e0626786;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5deca6e683e261fd7757d046631cd80efe6a39877ef456cdc7d17911655edfde1538496cb0794b460b7a1b54c3dcd796dfd8da9afc4a105e1c3c106bbf0b9997d0781f05c42a77e765499eb30e41a827fb698c4f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h290476de647bb73e3413119a103a89d0d79c69c62b198c97a988af44f3834dffbd977e87ff8373ef2319997021e0d16f0dff72f1d593a37eb9f26246ecb1bfc1d00e27348cd8c9bcc7c6dca585e45f10ba7570152;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc8114ca7a04107559f2611633ed6b629c8093a826cb2ac90387619baf092338e2874197f186d3359f4e149e4a30ff56d772f07d85780fd451188e752f4e98379250a06e2e63e057180d889e65bb853253047f010;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf88a3366ebd710dec1780690d08e01cdc9d0ef3d1322d9e21a044abc65b4ec42d4887fa9b4131c6d0d4cd0ebf8112401b42771f17cc70be4e83cb9ec95827792b110a587591daecce5c62d7647c4a17c88d538562;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h931f2595e1d57bce9687f83624863e86b0ed95080e07150759010c3681d767bb36c0c8649b74d24d49eac9a921c54efe59bd8b4a60771a20b78b46ef53473fbb6cebd2905b2f58f71f795a8375eac9ec9577768d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h866086e98eb4af6c5dc5ba27a30a1ea56d0df6d0e71d4fc3fb7557e59b36cae9f8a908dfd9a92003195846432c5c85603df73631b4a7c3cffdba7023a37b90d39eac1ff7449150ced13791cf880c8ff3e06c6ecf1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68cd6d41e6cb94d83e3df278e15c430b87124697ae9051bae7c925a90256cece961b7bec97557e4deeb15ec39718372be76e45557c1a20eef735811a42f1084c5970eb581b540a89531fbb0db2ac00043ccd12f80;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf98cf3736eca83b19cc85056061e16571672c690a95713a73bade6839dbeb7c92e40eb5f06f0445be8610aedd24a2bbb1373a85b7eb16c895870235d6797c78c1131b3c0f9005fcc39323303a769ff3546fc0ecd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9474a073ceb392dc4f0ed838f23c219fcb663b7c0147718dc2f2ef1e3600dab374e587ab3203d7830dad36b7b66590e8b2c3ba5a9f22d9f056ae0ef9feb7d838caee2cc435170577d07a421297be99971bf3082b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1bc15da449d16d302f53943ae86770af4b9c919cdeab6b4ac55ac20b71b9ebbf31d040c8fa61dffbdfe281dddfca4c2445e2698ce7abee21c948c11759b9a76dfe6a8fb67c97a378a17d64731aa5d5d79e63583e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5983dbce86038fc6ebf72226edf6f52915bddcc1ff3963476e0be3f96da042e59855f1e51ee807e36cbd69abab71e19c939d76cbc83b5fa239e4d725d7ca6bf96e1fdc80b66e5a83f6aeaadcaaa275a7bce24486;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha521bab00cdc19b293058c587b79422847a1957a41dfdcac9fcd6f4eaa9a684d9aaddafcdde7b3a4fba5f21b44e6181ac2206f49b395a4dd5c8459ee2e8d44324fe15b065ef2b89e78e8ab54e2b338492bf99b6d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h887bb5d704adcbbbee7a33801d705cc8a4bd511b045821d70665b488663e353599c996583b2857a80dad413599d8883ef1d8dcfd1e022d8a88606c181e7c0fa76b0c5f18ccf06a582181cf411cdbd92a09477b217;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e08f642a37f79398a62b3251227e9f494555b1d30fd57ef63943e9d84b5c606eb5750076f84db9836e5d1b69390ab6f7381970f597c14f2101803fb8f66e7276823ecb91efc4c37053b80000f373b55a2c6b30bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ce1de2f090e9a0af62b6eaeacef9d4499439fdbdf287baf0c6a6980d288a73f4ede255bbc674c19f3e85951a6b3ec9d9818b4e96aa10bc35ea50891eb2976c2f11d5b79c1ec02afe4e98ebf5912978cb2e929deb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0975e13e9003984cb80e5358cb1164c733683a9a016ad3d1f18e10ce52196e792a7b2a0cb6e045275f8384681b919ef88be1e016f647fd162c038b776713f04942844fc21aa9bb526f27147aa938bde7355e8d12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e21572a3eaae156e45f68394f13b4cd0666380aeccf7fd3b5e27417ee1a62b9b9b1c15b4672a48144d4829015eb526b7e721dfbcaf909f63f755e88d1ad675c732f04d0b0a6063f379e592b2cb086814372897dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3022c9994fd6ab69361ef7e50fcb4281d3d3336f070da5ce57f40ae1200ef391ee031285f44e16950f26d0a3ea01db131b01e44b02bd09775e188cfc1a3019a6a536768cb59873b02403250ed38e5502840cd927e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf40290c9ad61c28765d2c5df27c54b6a26c341d28c7659f6f18bf521807bb2afbb0ab3d939229c0c1851825229bb4f03f97f40988fb8adf0b0507f0e4b26c5c849bf311e6d8b4ef4c9e7bf356b6bc1f471cfb26d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3ad3e232001b59d4d9252a2a718456c89d8b8a301e5248b6a045c611aa1fb0da3344f64f100ac751959acc806c892fd69121d093b16e7469101b0ee1eb4d843bf7e5aa79f68169e69c2f49f94f531322dd42d76f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c6a3e4f1a18cfff42bd353920fb5a02c960221edbbabf52ade9fd3a1d9f5f0b9921411fcdf219ec14861a79dd388298533fcebd4c61099bd0208dd8ce414b41be72cb5cab00dfbaa9c4c62025f44967e8662abf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd5c88527fcde0360c168af78b53406d0b49829032841917deeb2b44d21f6e510fdec4ba4b401a8f0f764791743f3dbccb76bb48633f6a772b0ac4f0872212117db5af4bb2ea756eb0419bcf10666151ea4ae3d59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb724dbdddf88c087e8d01437fe1cb043ccbb3378fa50a63af13a493df2ba7f252846a159b897dcce9dc145d0555490bc1c57d80ab3a96e81d308690fbe5be90c505523a9c44864a88b4de8ba6be330085ad8aeea7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc6ea188faf26d77ad16b90255342f01462bc52a481240367d7a797d38dfc163f2b851e78dcf5624c0b84953cfdc0539e4d427c4f2e331dce127b5d85e68fde330ec6aab1838506a886639b4a0e632ba3dc11022c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb877874efb9b39f81c2a4bfa5fc52e3abdc46e5c3cfca57c0c1187caa7d40ce1334813f32c30d8bc0aa9c9c26251240c3d1426692611c7aa663ceedceec513e9615770d3f33815fdea2d0d0ec6a135d464e4ffcf8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bdca30b1754ca907b2f6242dbdd4259ccfdd5ef1bbf14440c6f9481ca9bfb7689e85ae8d50f721df9e465ab3eb79f77f163fd652a2244623adc88dde75bcae8b36226b9819099fa90a7b9476eca9a23f922992a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h140665fc8f431b459b1cf46e5f48d53323c8df47fa9419eae945ebe1a97968d981a3a1b3ed6294ad511796428417c0db4603e606fe195b792fccf4d4ddc7da79895f699cf4806b362e8ed7ad02d6d6668afec23b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a21acdf38d0d26ac0710f4e40ec982d91285dbdd44f1b57de0c4174dd351993b93c7dbe3785367c6bb46b76fe50933c2d767d9949d74147ae4b31ed3c69823bd63c4697fad2d59a16fbd17a1497fdd3318e3f9b3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda7756a9b9013418164260178bb740e3e964fcc01082449b881c1ae08aafbe1e0222643a44a3268496eb79e691ea5c18de148acd43ef837a3b3c71f714c75dfc529394ad5c16e0b2135e7690c5b7ce7ac190ffe0e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1092e5258e048a824985f99683e7f629a999a49bee9f2acb179fcb11157b62e695056b6af891c3535ad1f3187a014e317c631e1448ca076b9ecad4cf2e613e3f89e875bce7fd8944bee2024c5db0dd49847d82455;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f64d8e424dfa19673d18026083df231b869b3984c0c00473e10b1e2df35b7ebec2a366442d1d83deaed848aaf2ff7b6baf1f9e1ca415122bb4d8dfbf24b28bb33e27129a21a4df4be1bec85356eb062cdfbbba71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9e024dae878409af8987322320577e4fb385b107ba99918eda237d34e12277821661c93e13cef15a17220a8ef95206aa6d9c945c094c86e33d397dabbf3892eb8fffc9ead63f9e735142877e05dfeac7f9a5faf9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fb91692b706656683144aad466206ffc4e6889aa70e71ae45a1ea090c4e1153b06db2dad3e6a6eba28bceb1cc11d1b17ae3834030139bfef3d66b9ccf569d7340a9b2d3d2531ffd29593a1e8f02d0bc143ae59c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6608e8800b4f05bba00fac3c580905c3e3bacbaa971a370888d7007901c41190c64df01e759afa05936cbef8ebc6f15aea7b058eac1f0500c664e3dc011b67d2049d232058001b03a986ab52e4ef581a7650c33d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3019f7f8c00a46989850b0bdffa60e0191006ba51425b1bdb9b57ace98fa71721982676f0967253d970159a15180b6e7cb711658c038eb2af26600dbc5f0de2d5c4ae5bd5387a8b3768f253a6555be8fb589c628a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c21d6c1aae01b8fc9d5e92c2c4937f1e20ec3a1dcae9f312c707be1ce05bab955e2093dfd7a7d0240c1bf1451be7bb92b69e7984ceeb8344fd410632e41e04f8c1c59cbb449daa3c67ddfa4ed6f3b70d3bea38b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea1816642aa2bb4ce4e3ff2009f746053d0e94965a09a5ec89b57b7d39992a3968081b74130202c0cbf26b9573012aeac402e4ea093460bd4dd340d28409e223b7a0e540d0416d9af36c64656f8f6eeeb94a93b29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ddefae58f0106dde0e04e2bbd6d758c6ed49105ad82a39051971259291bfb3c3f0e4a78c7e6f1886b343ee80f979f34126eb265ed55fed04447450d97cc14fc6634498c210f96d69a9ebeca750e92c9db70c4c81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9203ca9159761083d16c6e5f32ed15b9a3bc9a58c26c545dd198116726b3675a14e5888b1fb014377d372d5d1f261b3d9da304463cf0bec0124ed28df5cf16eb0166b64173dc4c50901ea80722a2ab4e5743b550;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a574250eb5880ea677ce9323c56000330595303eb7c4c7a911c60045866c931396e4fb06e6a082940f2614582398c190cf172997606b70dc690740674a5bd624eb6226dcdea84be0e4cb265d13eedfec18211e3e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55ff124ba58ace467f5462234d494008dad692945ca214f10b337990a1facfd33a587797e1158eeca3fe39bc4f951048152c39555e6d2d92f9ca8d5b24d404c8c5e2a15e65527b53161a8fef46c0381351aeeb98;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ca31362317983326bf07beecb8b73020244692bb3d9745dc0dd1f3b413faa11279fe5cd50389518ca901c3848054253e9187c3817b9a2e8467e343f3d0fbbd96d78f6b354590f02a77448c73d2224ee2b6360bc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67f8a4180b63cf073dceb7b10e6e1ca7f2b87d78bb3627fc2596815dab59a6328f676faf55b9eda4db3ae89fe4e5e941e112af307662d8bc78a7780a9ed0757c91873bef43769457ecb48be95d9eb69bf90e308;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha67a76e3a00d20e7fa7224d0bda1f6f6c36e6820128715ebbd7c2c4132f9be945de74683150d3a484de0ec8ca703eb9aa56606b996be1a9fd1b28e46189066017de3c7c78ed62bdc58a2cf9d3374b4d8f3cdc77cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5846589abde7cbf84c221eca4aa8d326ce7bd6d064221155623d10d8faec452fbf2baa4e2a335f9277783b035449dfdb3efa78fc4d13af883a8345bc1f24cee5057bbc0894e44225072273cc7251e237cef97bd88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bb4fefe6208da63fa8e6310c1b759747088f4962069f0627aa5f119f33fa6b4fb5b6ea84727ec3d577263c424bf9d72a6d610fe72060aef898231d45570a73b357177c2224f60c63ada6a06b7265a937497cc380;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb0c7dcb73304d2a4fe113fae25c1a83dfcd82d0d6c09e1eda1c6e1dccc60b14b909a9f7cd23f46dbf90fd34649a62db040bbc66072bdfba2f8b5fa745393223739e064681bbad284969554a8d27c315418be6d39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65cf5408db63a48271431d166b410f58526ccde4f59ffa418e26fb51492a5f67232b724a1ebb9237a4081696a5ab5e376f67ca37dd6c138980d819aad1ed9f22ff893b6472869375598eebd1c0e835e675bc7deb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cc7e98a5651c903b4d466f07acd60762396d5af07d30865b6b16d1528a0093c09646fffb18bb5f7053bdccf3059a2e15c40d71435ae6a5117e5bc3019e9b147190daa329dd8c6deea2ee6e916f6175aec4dec84f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e8c611b35a938f1ec8f7e75887f4baacbac8269c0f5a48954da46bee0de9d2971083f5df3b8974403f5698d63c4e76bb3bcca26042dbe9816c895bf53e99a97a259cd7bdc0c1f79a222e203df1d44c974b4a1d28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbc7adcafe601dedc158989a5c49c01fa51b1cb82cab75e97285fe3241d71cd569f82d1a6b53b726c9e4ce288c21583823c01d80188a65404db174083bd392ced86d50e49cb352cafc1d78880093bcba3f3857f56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h758c39eb0379243410fd0253baf9bc94926cab057a04efc37a8d8dfa2ee486294145f28d32ef57cde0b706cb3d794287e7c71cbc257c284fa6759f3b391cc270dfe6311a0681ea5082893b5eb399735438c4ab588;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h231436c6816c5b7464b3b4bd44bcca4cb004e3c21cc9ecfd331a36dbb93539abf7246c1b753235ee14deea104e8caa5ba29da492a3a0c2f044d48494976b763e9ba3e878b12e8120852aeae96500e2e41db5f3ee1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b13b3b07914a9b1f6352b4ce0dac8fcae7477a0734dbf2c2b4f0dec01aec96dcfbad6538fab85fcbeae8ded9c94ed52c30b73e445ef15fa831cbf18dec05c4dd13c2982e4197832afb877cec9d97d4c98ae7191a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a1228b65a326efa93038d761371ebbe6da5aa57c48253754a6083a2abdc5bf405dcfc15ed1b7146faa1e9c125915ca639d62286bddcd6fddabf8146f7717cacc5feb2e78082155011ba383297ae0d1b65a63cbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85956fd0fa110ebe2e12ea1770ecf52ffa587ed56c5b9ce50909af228f9cac8e0bfdd0c02ca87b8544fba6674229f807778c9e3ba2f233e08f8da9e3a8b2b129bf0e79f11fbad7dbc309bbf13081b7078dea72946;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23bc54dfcd78559267092db84f8e0aa4be6f6b303c099cd95cdfc21514ac176fc60ba1a491912225bf935ef449943d2cf2c7afb90ebec3ee0e58c442847b103f55c2ca29c3b3aeb5184c209dbc5c57fc97cf02843;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31641bb7192df26d07fc1d85562bd243b47725d0496261a2cc6bfa20cd84ce7c7f831e2e44f54b4580c9d060cccf8b33ecd8b1fc21989cf8ed783770f04e4151ded314dc54527e48377b0cb1833ce09a1fa6afc5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27ad8aabf13b92a1a1c72245011faeb54619ff547427b1f79eb9672e62f8fdb033d12db17d83eb1f6293bc9b0db95d99048d9f5d18b6c7d74934c36928a32bf3a572186f5008ecbf1e12fcc2ea8e46314c5f42789;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha05f1688a9b2bee865845832c704df79408d0fed9ea12c2e41138f498f50fb929b353e7a3ac3c1aa30e3c0387bb3080244fb7752f3b78e0c9abb0fba379e8228d2e5e7d254ba318d6e34421cc77eacd898fb5d970;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd76d9192c9a080ac6e7c85dc38ec6714f1303e5f756f89b8dc5205320c69a7c7efc454078b5afee4faa33b0f65018a7cc57fc25d8f5557c31d5e59ee66314e0a5336e513ab03ba2b5b5ce80aea735948ece0dbaad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeafb2766f94a8fb8bb2261bbb430d7c27564ed9f4b4fcb84d6379bd8651cfcd3566a0d621ee34957799467cb66251ca25aa4d222b966a6778d232c0d6f8da8325f46892902f489b023686fddb5251bde51739fd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d8c62b3a042df449f9a2fddf1ea4189a07135c7ce2371347d7992953a80e0ff22547ddd97f6304cb782d3d93cfa29ffa16788bdada391c1da140a26f4b784f90a30f048802142bf7f319f134c68860697f2716b4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed7a16fc1c4cc171e9f1000ab134d740949d242f33e8e6f725cccdc28586d65a0c6e837fa73eb0cc866727b1b889abd4c056270d44863d30599a48f35955050e801e07766d35995c98741c3123353cfd689e47055;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb27dcc0a9ccf497b3e92abd9e26713d0a42a067f1a1f32cc0d65a95c118960864d261c99f3de11a8988ba7496cac3bed1e60d71afe796b37bd81bd3673dd7827a2c39718dd59f0ae6258af8002daef6fd04e10c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7be017b820c70fbf4cca9b48209316b250de8a1173024f670b656a60c4d7a3a5e587dc1bf1cae85c6b2b16af0e0cca0ce5a5d02c316bed9c362fed7f1f30218ff7185ecad71b6e8e11046555d02ee573986699621;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4562db7c5320e85d172331754077009d83a29bfc9d585e852c41de87d9c15f1e631a44faec874b30aaeeccada231ea38ad7f1020c0f261fd89f19218175c367146ac1f4616ed948176ef99d1cf55ba06b74a51ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce92706eca9b2038da85677032264cf4f6a93354a0665dba2274a9477225e19755eee5a9a20a8924ebf9caea7569d7cd65fb3d04d117067a14c860cb7c31b3ec0f66486cdf4bdf5b6a36fb10a3be49290759f693a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c9966c90cfbc1b6d28f7651811da4331da73aa130f5d9de6890478ddfce78a4eda698645bcf00bf06b9b1d0bbb79486b502741ccf0c507877f0cfd6fee2d1dce9c96bd9f8acc3f95cca5b751789da44dd444d079;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1222709e57b504c0aef989e611075385d16a0540764cb768e6007839c82ed7af7cf88cdecb54ab2d0f1e5538dbd951e9df95c6a3190af8c1727408ff828e058c272ab0b7ea5ec5b39f9f1f74c8f819bcbac0fef26;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2e8db405a0174c28dd572c2497ec105a8072be67a35bc8e3e727164907e8d683dd6145412f5f182c8ad5fecf66f0c8d24f9bfcb2ce154edfebaa325a8e0dc55a0e0063b8c25c176f3f89ae27db8e0dff732281d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he700557247d0a1171f249512f41afc000935c7ecd2d2aa1bb399d13bcfc9891d38a1c917eb9948b3f38145183cf540f2899664f6aea103066e58204e178d4e4aafdd7da6f155099b2567a5211e599f1aa4510957;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h863401183d64eae67a0450460418c0112b94f5e0c45205b84f1446cd0bf163d5f273740340b47d801327ec2d7eedfe6a5dd5db49496df495442da9c32824683639263a109b88473a05ca79a4d6a691ec0f5a244b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he56c5014c8d94471ce51e05cb6d14529b10f95df0cd746c95e258992706e929805a956d095f6d2bb4045026077f39e4e5e6dd375e166eb5e68e09b3faa0ba6bbd5fb70cd3b234d65df4524292b431526ac180dff0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h316223e0a42ad5e2a83e1f87b4b8ef00141fa2ee699d82cdaafd656cf084c2278487390c3e1a94037a6a1a646898fa5a7feb5181f0fb027cbd7fe0ff6f70175f021c9d0f5d2b614db8b4cffb91993c33fee007080;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c2244f613c6b07815a2de4a05de56245bfcb9ff4d0de9a29cb47ec8d1c4d79ec2b8f90d3c95755fcda1d8cbbfaa610b1c2967c95b1cc8c90a345216801de406380e534dba346691c824465907206c313cee8faed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2deb83d8717637750c10a99092f0e8f01145eb05b7aba86574d3b9cb99451604bc2b6cee57a2fa410ce860714b2c8d9c8be1cf8c0e3ac6e54d854ee8b9f2996dd17c0274a0a8ecda83723520ac9c4ec0e55a538c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2459233f666b090446babce8175636bf1692c7b4e3f4b4da65b227251c679773d52bbdc2f02366fff681d032e815993aa5cbbacb99c185cbf1e1d8a4085858a1a23f42e2cb390c570cc25de7de619ab5273aa6cdc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a8342263d97e8b9a8ccb4e8d1107c698eb0103979fc570de11fa31cd9f636347d53f21028c859359e2e5772627bab78933ff07d1fbfc2430cf6d22f7c66e83c46520289df8413e7a2888780a5868a49905c1aed9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb44a24c73d2b460c10de1524b7115d823b5dc3416ec87709ba4a8c48b399ed85388d92c8cd3321021cac39eae18cf871d0f6ab70423fe1f890d429633ed1faaeeb7e373d7b358af64f2d6f98698768319938f5f03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b912c3b1389be801a52275be67e215be5b326bf258fde31aa6f78709ef24555c81a2246e1f95cf2a209cbaf6720a8bfb6107ac6e32eb6b9efc87f05d81a1f39e1f593a60ae7db7dacd9945935acc8bc035b1303c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81d5285a59ccfcd04907de3622cf6edb1a36f8ddd311a62018687226f125d5b03cb7eb152ed1c2a6ac22c40454f8852fca0defb8a860b4354074a6d3d4be5c0e1e8f93912eb13ef2563e41050c4b6b40f3d1dae89;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55c8fbe6c6fb733bf3b99f455da2cc3dbdd98ef4f30d7d8598ba4640b33ac36c93a3c28be8337546b42a6b8b2ca18d90383fcd229003aa49b0ad17204858d971c888c036923d6e4885cfdc5c49a580bc8d8c2d5c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h462a2d146154419b144dcfa9e28f0625b0f1cffeda6ad66265e6955ac35974f06cf31971182cc7cd81d58dc0027efa1329b77ab52073cc36298b11521120d1b83cf50fe41bd15157ddb62e4d5f66eca8d924c7bbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a670be8ba64b0d70875035260bb6524fb68c778ff3e090fdd581a9956f617fb32b9dc8b3057465d19fe300d0655574006c548c44be934323d7e4a909e9f130fa853ff3a9a1457f3cc5ce6f5670c0ae89f1faff4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75a38f53c8a560ad66cf4f0183066636499e956d169be2f283f646158b955dce744f9d6db11862cee462a38837a2abebb0b0473364424aedc9bafd0d488cc18989732c23969125768e3b2dcea8c6a3f9ded9a9791;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81d7c2a815d80ac1d06eb75684cb2498a6a86155a2f118ef1ecf1a0cd68b242c4c69f60f4129019f260cc9bb271304f15a287883881e4e845fdcb5b08a2c073f7f802c8d85df8c300b6c6451d8946e64003476101;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bee05f0136710e67698f74ca9904412cc2b4defc53878ea19bd16557015e2251557fb69524c6761c70fcb3fafbaf680dde00dbf53fbdf7a276db0839b19a337a1baa60a7113bda4c446d63927dc061edafd722c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc61f521b3a1f1b02f5de69ec3d668613f710cebe3dc763eb50beda67927d2e528ea7a6a2f99f5404f050ce0ccf801821cea097a1d0ec81f3fef66bce02c98532b24bfb9572a729397906cad0bda5e1db296efb9d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha681717486d759557aefbb1cd7ddc0dbeb6002aab907e1e61d46055bf11a6a05ffee46bf7fa2ed53c42414f45b8bcf84abceb3e45588ea4a5095df54ea32a8b2cd0330a94a88d38993fb323b625a1dbe702bab0dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b55d00f577dade1c8311530010cfeb7a3049166d6d3d13f5176393de037107afc5e4ba8b4a06ed823af29b4a948d312fe60048003ef32be8dc5caeac9136f5452d933da8b02b58f1825de064c0a898c4f2b496cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27bc2e8f66b0bdb3c8e3fb774440a0d98ce8c64a7dc3279960d7894dc933f216c423d5ac704cd384a0839749dc729e4accf2eaa15c09d9c405aa2afc8213bdca79749b5810b7717259e60577d5cec5e4a9c48e015;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cc3f3e3cb62524ec396e4015b402686a7508c2f88757106fc133423cf7c4b005f10a7115567425b6c969011e925aa4e2e2ebc4173bdc5bea980eacc05cffeeb0de75252e7f0bef5ff70776f020f4dcfc834efbaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb983803d3488f6fabc9c816393ec431a2f8a56d6c57f4ab20f187a52bd8555cac13b2564511aede43dfb77d8413c13f971d709c6d06b4a7049508134fa248f8717898ba49ceb123c2f5ce4f068b1f74214260ee12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e5611f6852c774ab1dcaa45473d07ba19089d3850982efbb5d417bb9f6111b94c57cc365504b30ab2f3fce7b1e7411c25ac0fb82e64f6dd809c86da9f176f2bb9e479696ea83f5e042a6d87c99f08838f6f28d8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4470119dbdd7c57d5c5577a030b0eeaaf4c04163acb992919943591eef6f5d1e93c4e2310673b099bb2760e1324cff42082ac57e5cc9509e1f6d4149e5fd6daab94c2a2b9164176fed52c09b05f869c9104beed69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f54647d38f954eed0d80955cc9b439346255fcebcbaf6a47e9b4330e7f522c5e7e63dd2982b5cf119adcc573e39eb2ba7f44d2361a8091273353a149cc91e6ab0aef90c5f9408e08ece4968a495cd0af0e888e69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44c77f847a12b5bb342fdb471d93ffae03bff74350d1ec7499e7b60316d14cb971ba02ececda2b70c364f836a20f985479a42d3ab9509147e0b862e6cc722a78d92f09c9e349d269407955c813179b2707176aec2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c0b12e7c7e319cf40ec72611a1bea13dbf7221cfb50c63e5f666237be2fc11dafecf31af1d0c3117f7d5fbff8d4340a79dc5e263f144065eb78cf515597fff85c243bec572b4bc0588394cf1441924640a3cb19f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb429da163bb33fa28b6ba50e093a1404984d7d2db8e9068d52d87449f2e4b2928819d5d772c3b16ea29074f804936d436f0caf7aa639d28dbcd016eb6b06b55983759ae1ca1a6d3741ecc62c5b60c17651c4914f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d741c72cf02a468944c3837d5ff3eea4b235e483a63347ddb70ccc2a2d0a5234d235ea83898fddd1559d92d23e9c4a6b252648c8f68afd17804ea930196c71dc8a4669820cc8f48979cd8bd48e12f7d1a5a86ba7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9aa39c5c71a94b7ec164e33b246a6fe1f4d99fdb0357c80cf472e089b44787cda51364ad48898c94615c0228b4378c31c63e7c5fe9a6af5d2310da632f4d2b9d24d754f7f3a2eb22ff824065748946726bca6f0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h643571d0faf89d0fab07a4c79c4ca632db018e9316772b95d68b153f8a8ee173ffdc89da9be28e64066ccab7a600e33f2506b2866cabd50142265de719bd1dbb339fb6536ed7cd926101c04631cc05255ae174f54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c8be4282a35c86e64e20dc2aab951c0c8ce9cd0e43b8ab053d847fd5a0f405a9a0a9eb51a6d97235e818125fff35ae9def7af95ad190833fe8bbdb2ea0c9b75bb9bf18d0738f1a26798024627c694461fbe9e0fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e2560cc3eeda627b684fa9c8daa07ffc3bec41d91f986cc73bc36d03c7445c5a7d59e322eb2a6e006c054f489fee4761332ed981ee7fbcfba2ad877ddb3d145d32763cb72f49a3b6ffd7b86927567a8fb69ca22f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55a8880bc0e08f2d15e66df3e497a50ba606369706b2e6c7d462efcce10dea4dfe8e506c8e01b263bd794763801e64e2bd0fe163285dcb921c3528f2d4b5f97f53723e223635853e64ec504a600bf3cd2c44379a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d175a73a92a69aca0468cb1d9bfd1ec3e379ce21fd6e47b5d2bf1be9362255520661842b1b96b11fe3cf39b49c5346c834fd54dbc9ed72f500d149190ade986bfd1ef2d66b8c7a0646fb27b2ba3bb8d6ab70c970;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d92d722424511796bbe3809b0b760549d9201f07a9d090b21245de6b0b42509f38e993733616009743b23a28b48f9b7e0174f464b95c9f1cec3adc381ece5a8590f51688df1873362f00d8556462bb948ec44e2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha91e0b0f0ecc0d95f872bca149c49923f7d19bf2c6c6b2d0fc8cade7d51b91a61912a1edb3e1d87865996811742e22ec08c983fe73a0c5a09c98b9b4eebd5b40c0d19321c511fb0013039f2eeb0aaaddcd4f874f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb101ab554a06c84a7523ec1080ce62becd7c0d42ce6d8dc17c1f15928bf4414e69772f401d71fe5b42cde24f140f9c4007403db858c1d11871f1bf840f58f0a60eeb14b59bd94c2225636cde4f125dfd6ed45ca94;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3448fc88e79df1ad7484696f2a9f36943bd961159510f097d3add9ce2f47c11680a4e2cb61026ea14f44bef47d0f139323a156f0407d28a2d361446310380947bda0c7f8b643b5afeb003dd2b0325f4ffbcac417c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf70c816b491b36f74f147e83b2d8e8c26e5c59fbee1245a6ff5309e98102e6ca9f70fce3c9611f5b262859d3fd422567d8ded82a80edbe8047e30d20b405e4e81ce4fe10d1f83895942be23a72fab40748d52d0b4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67cb862a09272fd45e86fad48a3c53ffcabe4f76a0dc3c5b706822c48e02d2ee2aed1ef3f234ab9cbaef3ca6d3264203ee58e643f2b18c72d98c894a03c8c5fd2af008e95866aa9bff46dd301beb7b7ada9b7d72d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b19b0ba2c616ff2f80ee4611acbf3489eb5c82880562ba01b877ebd55d2cbe3c9894a11152d4231cc876cf27565032241ac9e6bea2e3dea0f87357e247a1e57ad5f9096ffe5adeccca3819dbb1b8960f79c16327;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46258902acf6d6bbe15cd039e5da1e0b377e96175d3ceceeb71248f69f0dc4c8059ce4cfb5c1ff36ebc98565ca7521fe8665bbc59887b465f92d62e9259d79503fb78df1a5a5b9cc6d1211f39f318c362b4bbca86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8d7c7ed2e025645c25e2be2b3171d9b73be076af45b48c5f295f947a87de7e384b48d05e9a5c93ca8eba0233335d87c6cf76f7dc138f02c2f8a938a818fd36ab9096d2eba4c4e8082274807cfca9981806c63403;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a15ac126b7e03d83b678598b87fdae5542cae80d6cee56b2f9cecf9bde412b0623880a67eab3bce632bf9dd5370ee4eb7f218f467ac61e85926595a24f44707f4fe3c1668744d7ce7a8b5da5f434d3034037b32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4b86862d24aea50019a5e65e7146f8c8183232702d1c19861eb465fa6195022a6066d9a65a0578aa3deee19648ff9ce2876117df1696767a865f56d8bfae7d5daa879f30be455f7ec20da29cefbc0e4560d0713d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h908f7d742b348f0ec3fbf282b5fb660d352cafd73bb995bb07710636873df020b1f16505b76bb6e5576ff8bc854129c7e26de66da1281f33c3bb8281c574e821fabe3b3e4e4954716eb55bc8acf6efb670be21115;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h704d1d24fd6d9946dd7dd55062d4c4860dd27929c8ced3615548bcdf0f741e20dca76add238b49153f14a5978e22a7d4c774e3c23eb86d6bba8f003704015a9f5d9020751d5b75a58ac8294811912eb19cd5476fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b1d0da8119ab11baa7820a2c818741366a66a1d8a6734aae4dc958f7b54197da57b5bb556f96c2508ec88f940f3731aad3d9dd65ed76e0221578fa21988971956277e38ccbfdb78deae706858db951b3264e7cc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37006ca35886930a6fe0136e8c88a6b3431eca6ef8367c554bf58b1b31c33bdab4d1ef28c7f42688b3c35177f183ce5b61bf5fd6d083c0b24cf4b236d815920b691738633981249dd8d1f302e3ba26ca5c0c40e21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd79d6d8501c58980e69af712f1c1600727ec01b3910836d6211c3bfe9a9c08a8657cbd386d6a150cdb52b8bac1b360aab09717cd2ae9b2a039898f1808bebb857e6ae9ee11970dd91c4373ff3ea2893dbacf04d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf351b58fbd46c2f0b8e39a5b426dc9c0e5d5dde6cc11c3509fb2d1f639a096a2d0e2412ebf722469dbac61048719f7e1c702c109c4395cfcd3754beff9e09bbe8a6acbac884fcf87857d429565b4932be30ca3c87;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5fce62a1c69f17211b6f163cacd320c7f7794b4e7825caf5203c87c995432f57fbd6708aa589c84ed144e67bf375c2f7e860f28efcb64c871cc545173387e8f83d95c7797fbe7860b21548dc50b772a6534aed37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4a91fa6de2f8d36a64e8c8bac4e1b4d6ce693d2369cc6f9f761f1e1becea17bf929d2a3042b9e3c573e3730a7f6b56dac152d466600dddeb54e710c86f8e89d0e8df5ae5627b54aa71821be05d7d350c2633ba3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc575623a6e37bf6633f2cf9d4dfb886c6cd96698414e02cb82cd6c125c4a62afaa6ff1919aba9c4c54a9521cae05599b41d6e9e135d32e7cd7bebc171169ba4d6833c6a21e60fd07819c17cd65eafe0cd327c6d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3d29c87090a7d0cb7be616c70520400084475ff0fdd048d8c750f5eb20101f536ba5c002e0c248724e80b7a4db17a5ee26b294b78f8ee0cb59798b1fa42b2be267868155308bbfe8a3c9d6a763ea81048166cd3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dbc2f0bffdb4a652df11eb38d31fe8b6ea9db7b21e717670d10d577f9b7f12771cefcbdef20ff47da1c2f84762e756a7790d4e945bc1a970442e007579744a16e07b1ff8ee54de22b11571187f01126664e3e475;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84efa107de70263eca23ef0dd624fb983e764feecb497b4b9034c21d18a0436df5776c4051407db493e063e2aff5fbf7367d15cfe140397f938495d3d7df7018af8e707e5f1fd6422f070f4a5928ac3aa9f6944ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca2177918e8973cda30dbd44a48d95ceb6093b43ff68380f72e7741d3dca24fbe2cca9cdff78f0f7cc461ebef77fa686f829402bd6b12f69afa7a891be1a8274e85906acc28d56436142d83294f25fefb8f015ccb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea49c228ce96aba0f3fad3876ad8764100e2e57ea0f3233fde51a34e8b4b37f882b46eb65aacfe9d554dc73b0864000419e022a9e3a51b94ab1fed5e961b14ffa5634e1077e0070cf9daadcd3b3ee86a77be49b7f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed2f80b0d4d9aabfa8bc2cb2585d52f09f5c44509045bd490b8d07709e2e5276f89663ddd48652bd7f341a6cbf83f910678218c73e004aee6030e7c378d323f7ef6a2b9040fbe226656ee546de2309acecbb0d7db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1715e66fd4441f22c9d1b70136cd4989059d94d82a1d4a32f5c62aa273433f1c35bd30895503a48dc60695be3069017044dc07424434fd039a49da66bc4b554e3d009c5598562c905de2ecd8f5aad3ee9cccaf40d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haef4a399ac290f7783d9175115aa4cf62236625fc1472f1c6c575afdea32f5b125e590b4ec7219e583857a83c73ad8c584d17a008655ea60f5b111512d8db7414dd8851a37dd6aaa8a93548e144295e357506f625;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1593c48576b1ea9a30abd3b8c7c68b2f889ce895eaf3b80191ab1c28bb4dc9a872de1413424db3fbad605a5539a077a993032df3c79ac25db1ba8278c893d2c91b77640e2cdbed27a88f4973690ded753069497d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8827038d659fabc6f81946a266d913d3229985d96df5442ef85b945b2ee59e6a3a1645593e79dafec5320e16d49b0e9e18ae6a77b458bb2ccecbe72ccbaad8472e19a11efae4a6537b9cf24dfab41733a07cfa7e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0c976e25aadf8737f0a3e601008f8dbedde167c1459bb006c8cd17c19033ee766fe95b8e5e9f9daed8d568de5b03fd9c4e593d0036598f929a09f3943508c66e5e5b81ea90f1d5ac62909f6bb12309dd6770e769;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha209016eb0cdf476540aa610b7d3eceaa1b644420def5db65fa59c1d9e64341ad3450bec8718797f916b01ac1105a557246c2062b85e8942d81878c96ae23d232d20a069271fbf8d1ddb230ef1de550d69e69934f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30c8e244b7246f0faa658eb98b1f39f2ee3980c03441996705569f3e445a3c37288ae988466c5d22be644353dad879252964f30a4cb4690ff5b94728b25304744f7febe21059d66b65e5d8dd7c9ed728ce9258b6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3496d97b433b494f236c27b290ba858100a2c9494ba68ce3cf484d0ee669124b23387ca4655bc4b51def26edf6dbc3a42ccdac0691731ad74d6c7080e7cefd7b73b1290afc6b6918f90457a15dd1043c58d84decf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf28fa06e95d86976f012af3984a630e3ec55096ec6a5d8924008b15c529fe0d55788c02ee9d40198a1ad4236b0ee5a79396685cee41257d74a8cf8138057dbefa1316f9c858f2549c51dfa7ed1aea33c82b80096a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37e1d3156e65b051124f4d354c9db1b6ba4a5c57bc17b3b0af5d492e4c74822c8cc5c4fe14b1a03500000153b577104d967b6e083521c3d86ce3dab8b988ae7d9940d4de65d4e48e61d92f8d360384542827c642c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97e9e95cb51520f7630e250f43359bef4b32be66cd49cec96fce680928db85881f8f0d858abb96ab4f583266ab4f4fe9586dff04c196c9acbc0960afbf2edc64e18d7c498784f615575988ce522a29dfbfa6e3409;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45068bf69e84ba8e25940e9a95aad1ce65a89bc54b46037dc0175a45bca849d204a4c3b4595e69dc6fb7764612c56277582e943808fb846edaaea6121f3375dee2616fcf65502a07ab3beb05d1cb3224100a97ec6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b9bbd5da4c56c734a819e52e0514d317e14d919ffb7a60a508e358fad1d544bef281edd0ed39afadb2a34cddb9f4c470f6af30385589474eb24e16e50bf515c0636f0453c5d722d64549e3461788bf295ecd4f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd05eab7327348addd63b3fea0859b04d080d22104e90ee91af5e08954d99517d70f732c1b7e1f723975ea5bce05ee3cc5c55f54e65ef7c020ab56a61d96870cf9dcd2f3ac9f37ba799ee90ce7040681425ae93578;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0b444e065a0a11f0d03ffe2a03dc92e60f060d6c6087df1ecdf5e52cd2c02a42942551bc652c01de2618e2025ae841b776019b62c96a8f7ba1aa971f405450cc08f4ab7092557a40b08f505310ba61a72ca8aa46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de2ec2c8105553120ef8df2a4f24ddb5d5a0c22e117bf9386a08db5e3fe9ce150d61f4c9a6adc3cc615444a6f9920deac3edcef33c9371c0531f51884d3d1910cc3803faa1ff8fe70b77e11f156557a958eb69cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a24761191aa06c2c45396c4770f60198bb7ca6d5663e197e0cec811244fa5a580684a52d1d7afd98e7815be46e8f3bb4d9cc0086558fe7eaa7a45cdda6463388b07c8b4ce35a581f8b35c255f0282631e9f3f4ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had31e9c143c698d0a85eb7dcacc69fcec088c744a341cdf10976017975b2c41e712627e95905d37d5db71946a904fbe09ddfe097659d2e9b950f4fc8590e19726af11ca8756018c9394d4d6bb386b4a3700d63a86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b850a96d2cc45cbe4a9e1d1ff3df357ca4cba0babc56bf21488d96b7470119d40b954507743562e720ca2b80bd56c2c69e159a9e7ae27ae656d8a8f52a2afb77f9b851bd13295fe814629e3b962f38934a20b6cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h938fb496da1b49a3149096e6c71397ac8907d11dae869c6e7e31485fd5c573e0744f747a3a195e51b977e1311e8f2458cb621b0f4b49a93df00b3cd22797be2c19e0c923c144eddd9a381c5aaa5f824688b85e4a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb114e67cd20bb6f8f831de2eedfa3cbd1573b78ace75258f3065330a7da2be77ad575627c717f8349d293216e32ffb6fba78c30b0213b60ab71eba7defac89e385d3f4f577466229119ebd8dfb08313385c23e536;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46add22e5d3727b7604264889898b999e37917647c974500c8eeea213689e93106f9201222902b46b357c51f4881c28a6a10b1b3420639a76264c8b2cb8828d16507f6bf45a4dd9b4fee66ffade252dd6c4927486;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ecb0594dbac31dd2d8b91f33b740e740fb6017aa0ab273c7d7a175c1dc03226ef5329ce1f69f7ac9b83145b85f214c38429fe14f6c6f16bb91cd2509b3404cadf1707b5986d463cd27eab25c13fb30a3a248a934;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7721ff00cbea97393741e63a457fab5dddeaa042ea0207e7f5eac99d43b40b7a1e499fe15e9e03f83f26fe73bb941c860af25ef03d521c6b6ab980f51143e7af18ca9029222352f72bc463a03917880d1faf32cae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87b4dddde5a0c84a14df2e60d6396cf13727056494a46601632313288e1efd1774be17cfb212de71e6b787ee288c885484e90ce927aed7feff975ae12a2167c75e18ed4ae9d34d9ef3f97f56a1ac99a6ea9881c74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec882dc8451f8f542cd9b715d3453c4adcfcc3926732d7f20133ceca6ed9795084b199cfa046266961fdbbc7d46656daebd1f89187ce135ab2978a62158291373a5d1e56335cb8f70a7e4dbcecb9aeaf556ded561;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3619c94dac814ea943c9ad5e49d39e3685567db4a6f54828278be8b6b19acdd43b6fa8cb10c4f25cabab428b71acc26db7f10f6d2e1abc6468a4e10656937b293ab846e5020deff472f1a6ca61e873fbf68e6e147;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c013508a51a3fc32fdf714c6f00f3185588dadb366a0618f5504c2a5405f835c97a16558f9525b13ec92ea8f5367c27db7b1f9d49b7d2061749e5c54843bf1b1dfcc392bace10cd9be0312286ba5dd545f579edd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4885e577e6e631e7881d0e4b5e6d253b644e19d55c4d1bd8417da7892b6e3c0e8a60325f4200344acaad78462275143e0c1eb95fdaf938cd541af175a1a08f7274133372177138e673efabf3230177f15e991829;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0d013de1d46c36b44b15c88ca9e2b446384cc0b3a82162852e3cc1777e9bef865e447cdc6e74813535a4bd0ce2f0a8ca805e349c2a796674a29b1150e2877f0f6016a060da631dfaa7504f634d9a1b160d96b923;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h879e06093e396799fa440b07fdae606887372740715f846f687b7dcfbc8fa49316414f76aa38b8add59c4ef22e1b3c5476658ce59e1e17b6f47c39e2cc9241e7cfb6e2ad1e0afebcfef692298fcf0854933353ddc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h617f0ce0ef22fe9b24ca505441a16966764accbe7ad28a636d57a062618db12b2adba821b60afef90f848448dc95d7be814f74689bbf5b94b792a426810ca605bfdd1433a6f3d4d16cf07a9581828fbee35afd09d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e2e6e1b30c2d7d67623ae22b80f25df5272dacb8989cc880fc71ad116c9eaa099261610385246bb70c5d7f22c25dd7aed82cfdc4a91a8d9216dd06544cc9cb2e48dcb710da99d938f77e9ae7f099eaf2239e0714;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h264c053d6eba48c21e7e9849ae174c2b2267075bddb425ffb7caee85cb8d5bddc598a4d7d99592f498bf3eaab46e6a7b45b4b483e35fef1d8f0218a1b0b627b562f934b308879446420d25ce03fedadbb1e71747e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79bedfa7495b6f6629892a5ceb7cea94b4257a735f2c3103a75e5b8f74d43b14c9ef1d18c1106b27b9a13f425b74d27b3acafe18796d1609d8bc78894d29bd27de29d24bb528be62ac2b5459fae9a6fe530f61cce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c6cb71753d8fa82ebfdf1f3902d90770e92041fe7283e5597bce7ba39dab8060e44a78c5dee4fd976b647c58ca5b58170a26e0a8aa5840c8ff315de7ba3ec584531145ff0d84cd1f390a71411ba3b80e6204c28b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79cf24580d0090f5879726c4843677eb678991549328ca40caea9827f2ab447957dbf96060d3f712e790c0b6a8e78dac3b363c58673e184077c68387befa9dc209b2dda9c14fc16ec1ee057177124772487786b4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha23f2948cb3e46f61f2f0140872047b91163dadf727ab689edc828f7d42c8503953784eef0411d9303ae6b4298f7b7be634b35fb658609616313abb1d01ce51d029e9ee0ac4838f45b4a0f01f6f089ee9bb22c507;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb430ec5b6983dbb95d6746588f31bd15454410dfe6d3671c47923cac104911af41aebd337b64a4d7094a6c808039539af3a1d2ca0c2ca264e1e5ac01d06b19edc59f378d8b54502668c64c5947b6b83fe6a0c1249;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h286e73335726f1fc4be5d67532f528702c3cc800660860c5208a4589419fa9db2da061ebb5ad2f5e0cf54aa7a1785532c224798507c8ddba2925233411f3f3d9a126ba1a648b7abab0b2c7f9217019ced5b60e8a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cd132a9a2f40e26bb65364ceb730ab0b3f0a087c9c74ca3d0a6c132e3f8253c88f73fc6787b35d19e8ce534a5c84171d18efedb3ec9373e099ca4c30dd44f75093e1c224bf8a19d4e240fc648f27685572ce0880;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7abcf97169d3b9f60b12b0c4e66120b20e9811e4049031f5c6318a366fcb23cb688ed241e8bdbf0b99bb0c7cefdf50462093f25e490fc4e93308e31485e8426384a2ba0909d6795a63343e58a49538efc3ad81976;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc90df69606237c6f49406b82fddfd063084c8113b606a076637776ac607771aa67196e8beec0ee8414541d85f41199732b2f9207d498291e0a56caa34a0becd8c282d27b9a217cb31714a62c7029fb881a76dece2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb15a4443fc9ab3a8799f693c33bb9d315929d1defa9e2d8265115ea1ec28c58d77b3da497aa4a92bcc03722553de04490dd568e04b54ac17278da474f7611321296c5e8815848dcda7a1b078d44368f1a29d7c7c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8233db854e7cef26d4ca67b005b9a184d5ef1cf768ee3aeeee3a9e35891807248acf365811d5986549e7854cac5e2079d38d4466f41956240d3fa2e896b192c9892e74c6e60c577756597f29551381acd4d288a1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfafae868ed62a899666425bc41a790f92eb16ff2b42fa54bd66f441d5994844be343f30cb5f3e90ce011c9e0c12f6544971aeb643d5d9b93a85e6a6f72eb1c28f2a78adfb3c55d0b20cdc4d699a206a393e2650f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4436899bc1a2b5572f4c231144ac9c97fda8aa178ac5e941edaef02a007d61eaddbde726c84fa90e6e764aef7ed265a2b679cfa3ee453fdafa79b7b02a77c84c4e83de4d56f1d8f08d2003da9ae9d008c54e8990e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5622cf2fcf707dc4274759bd6c3f4ea0c56c2eae6024f2c2ee2c2634792e73cc82a0c20be20bb4ee00e7484fd6ceff3bc9156595ee64d724b0db50da7871d2f40536d7fae78e9cb11538df05e6c3ccf28e325f95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc792726da8ac42cbfc98b598f413a196c73a442957f20a36ff1f25bebb9c2219fa1ff3d9a1395b9ad2bfeb745620e57aa268d1f6fd278fe6386fc4f02232d010eff5aac31c4431d332c45a6f5270566f3235b40b0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecaa57fb14db3cb30ddf258f6d60653eb43f24b4886b37202534072fbdb6d4c8b6d112480ff2662800821518eaa414014fceed1ae32d86861adf156270c1a645bc8559818422a42ec7b02c3dfdc65d2d7e4f9ebb7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc48793e97653feb58ec2eb723b0be3ad5442a20a410c7fe5f716e87e836217e7133d4ab6df136b15e61b7a851b6df2bd6727796e3d2873860723f6786106c18a88ce5a067798c2538bafa87b7d7bc5f61ebb016eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff68b8caa24343617eb4763a85f5389ceffa6648703455897f966fa1f007ccdd76aad9578237c7d0ddae922b787299dd6dbdf2e3d9fea75200185587abb9071f861630ec841a8947f86e9414dd2425f8ac1efdea1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c1198f3496d523e71c174c76c60a709b56ab8845cf87bec0b8c77a1725e579d7002a512e8c9ec66e431014a0262d955571f58705aaf5aef6dfad9ec3a6f3e3fcf2ab3c9015c75f99cfe66b962989a94de969c92a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92ed540b3a36bc1f9e2a19196c915853cfe94599107205c76eafa844b0b5b7821bd087b73d9cb9aba6d10576f7887d1b20ef171b56b62b2b4d620d99f71a84fe24215bb519e033b2628149f1931b6c8e1cbe29c82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21e8e7f0f34217bf0bd17f4f5507c688e787b70f6495d18cc39d7b5b7ec762a5b7cf31d05d3a791d365d0fb605fa1b8481d60415a4515714590b6fbf401b930de5eb908b4aa72e6e5a9c9c8d4fe1c512a5425faf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf97eeaa673f3ce41ad48e5c39e35bc751ad62e1c099c49060311efc5e6d0f9c38459ac363a002b97ca1d89c62123ddacb700606d3a32c0b2ca78b2e10c8837bc9d173daee6669516b04d48d4715551c99bfba3cfa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h109578844b5aff43cfefbba5c554ebbbfeec024bdd8bfd1cbfe57052a30558150c68d6be1c120f80da1e63c305e4e19d59daaca7601cc1891ad4852ce00f21f1ce26da50b532a9753941834e4755d5b9627f3b7e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b6db8a3187ec4c94c781c52019fea21c38c08ccd7ea757c69241712f78cac2f844e7d4794b455be649e16669c0407ec67245d18273f07c6b4fd99a2db98d289ee8a113637682309c5eeaf4c3e77a107de4b4f90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he012cac1b17232f99c43a305e25731396654825ff8730f215f55b4cd70b2bd013d520c7703b1914dbe058340e03964d8571d5256f8256e0851c8ba0634fa3055c9f66ffb22aa2f6338d2165c8340d96c73e20cd49;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32b002adcf246f86193137d29463321066863eaeb35142099cc8b1e6e84e4dbbee94cfe887cd2314ca1934958a0abf5e04539c7a9e08acdfcaf13bd5022fba7e328c2edfb58c50c53b2eef4ad1d096ba786b3a7ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he52d7d41f514def2540922d8ab4b8115b1b17b71d4d8a530f81376d19e438f65375958ba9985afba1e72672d7f4b9c56cf725adfb9c35af9d8a2a9491e087307634fa4a914a978d4714343484cbe765c488ad7850;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5bce8cdf2479bf54fa0bab55ba154ee88d9eb8a5a0598f817bc60eb065091f897e84a3028d1dcddad6d3cdaf5aabe8846bca68928c80ebb617d5625644b96fa09a9c8323e86833f4cad3a74223075e6dc1e7685c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74d294719fdfb3fa98181689146c711be83bc1aff822c7c5cab05070f2ab8b6e81ea80a9769bcd91c8302adb131f04e99581da4ff5b3f99cf1dc8c5ae1834551c038b3e312d577e1be4e31c63a2c7eb85e5521c6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcae09e5eedacd26654ff7ee67d3c1c421358a8b4c22d8d8d75ef18cca882be855c29542b6fa335fc5b2ae085585d26ceb61b7659cd3049f4d9cfece6495cd06c4381b1325f99a423e5593d681e2ec15f9c8f59674;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7e89be89aec81caddd3335d89cdf915525e8bc8192e3d7f37de8d1708ce8f095b2a464f0979a19c0f70afc077dfcabbda71db877fbe0f3f4d34b9a7456e63ecb44570c9cee77197ff2533cc69f654e80b7bdc464;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeef598df0b7ee450ae44692c4dec2273a156182a1d987bf237042dca6d85777f275731fe47cfd205896f93b21583cbd93d2826e52b682c8f7dd6d2f4428261d070ebc440253f509e605ec775518ef701865dd116;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d1d97af0798dfa2030c0b797b085b4c1fc47a6b66dcf070e1239974c2e180fa48a82dee49ffc5fea5b4ecec93540f13277b08a400eb37f7ff192b27b9c42e5e537774407d55e0820be14b12e0399f59b8b76acaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee32bd8e302a31570664c590a6557b24cc44fbf0956372b24e20e1a8f1e235b871e1cc8d0b5e7fdf671824c5523327ca618df815a7b2a765e4f056ad65fc4db26bc30a19f25334408fd80f4e2bf2bb4a4cdd5d201;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf691b29efb07bc490f12a4a4695bfc8090497a7508e4c4537f0de1aa40b15bf497059068f42b750ff2e693bd4a995479c8881dd0567a061bd764369d0052fc7cc0f79570ed458ee6156d67d010e88c96d573eb27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffbbfd056093fb6ed28c46f6f57d1e016e538e568dca63716a6766e91537e228ee2ca7818fdcaff7e2685a7b32a07e5ff65738253de4005261a00b09542d6e8da6f06fb2e49c7f24cb05370ecbe3c44cd98e84003;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h158b26538c6b3aae4437a1fd517c0cae0d9f6f4ff2f65032d5cf297066334e5a0f58d8a9c134ab9b1f08db912867c2e43fda0c03e42aab29cd8dea04e63c540828212e48fa54ee05beb51a842709ce39dd08b346f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4d1e7b0917c7abc7748ba20bdaf60e351600d63c9096fab86ca8eb1d399b9ba3d1a868549fedfdfa5df1ceb6d3e960054cc7e2b9ef03766fcc8e68fe0db84646680864057a935066e4f6fdea83b7ab0c3714bdd1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd88fc4c29027161d3e05855bdef18699f1ef2d0b5d7459b946e442f71a2348ca2e826d101fc97786f3d548a1a6410dd165c97caf73226ce74502ac81272de054f8657a589f240e20d7baf309fde23b1bc13acd51a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h689cefabf8d6a37a561afa9ebbd937583226f6a434b4fb67f8d67ad071354cadaf3a479ce69aa2518e8cd21a86eb4273a62c0da50590f09f4dd73cee2452ea84abc933e845dce0990f8f318dfc2ef3d19fc195c33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc90007fc56027159ac46588dfb265763606d53be04de5523f6dc6786eef23fc9f07ac0e1bd955d7d96d165dceed38bbe5c0cba790c73cc180e5b424990c510b4aaca61becd52f04438bd357bcc8b63ef8b33d29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3377af132167529c994296d208023c768c63dbd1526f7b99763a3ee2b9b3465c665238ce1ca6342dbfed378bcfab7bfd35dbf9ba53db20c83019a47284140769c5e625e0b4763f140c9ad5be26b8ac2d5975da5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdde238ea8586a50601e5581966147a3ad89872c659976d164044a52e644e5b84b49b5276e4e72f335ed3f02bdadb35fe4025d4046fd1ae2fd738eabd9cd17efa420c0c6c18867e2740d155545b40889ecec8e119;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc37721a8ea055908056c469ce3ccd6afd5289d9ebb78aeb253e9a94affe41c1de6618ff00d5fe6e9cc5b6cf43123e7b590b7667b03b3345c9a00a416a1b1c28b0f5015575144205bdba544b9031c083c13a6265dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9411bd5496161143a86fd7070212eeeedc2bfc3b15c213b111919ac45d1447b551065a067bed2858d2515f0defd7fe0ed2698ec6ffb86e706f0e92087d31fcf69cfdfbcae8f4e5a67e01cdb311fa2004ffa6cf4ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h539f45a985eef3942d88fc16104fa205d12e2d554e445cbc42cad46550a92af7482af012b902f6b4b13232445f95efed988ae565a09e3ea194d576132446a94fb7606b14ae9d26d8cd8c83f5071cf776c260f8f39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2d7273c5212bd973481fcc9342574de7c1d1a07f8720a3b5976f4d151e31a4282b7e52056b110d75d47e683a5c05a6a22cfd44300ba7ee049df34f05c1d80a9ad63b6bde73e2e776ddda6a5dbf78c975e400dbe2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a5691b90af9b3b57abce28d87bd180d4e39313aee4bae091c63b1ed83f8c7ff514b7bd0745b99efc0a25e6e011a4c0252466fe25f2615bbdcac4d7b7b03b76496d517356187f34253caa4b487b2115068ad47691;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6ab9145896b4656bc48c9e5ca345655c7f6b69982dbb77fcd27a26ca7a68906e97c16724756df97fb6c01258564ff43abf8fa3517dd4fe3c9f73eb324e703121f4efd05094095df1a5064207da8bb09a5352d782;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9330a44c41cf6c2061b89dceb348a8230050164b934733e8e13e9cec1690ea7ff34fafd83d8ce2ff87861d02cf006ebbd1136c8b46913675da65b288d09fafdc8849edc2c24c240e5ec6388a38a15ffb3138470a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b2137ac2eec5f2bfaf0122310337d62f47cd1eb8a994f5562d3875e1492ae9f74e4185cd893ea85f6b802d2139fce8b5719e72d225990024816432a5cccb15fff2afd99fa93eff6ba23fb3163c29dcbbb3b5006c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dab58edccc328b424bed9bf7bdf3e92dce67166b5bd3653f591828947bb7feb6d817f5572e5bfde4c0af0d5fb02e77b02e2568a5004269514a4f91e240e382ad9a8618656a40e2604e36e55d71d025c81ac104e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44cf2001e43cc00839e55cd7b5ebaeafd507aa52b13b3527cbc952e02226fb6c5e7bc63ec6f8ff4afcdf510a629ace6a3a1a13b44f7467d213b494a2ccc1d5b649abf63f34812cbf421bf7a263f4fd572cac692f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee1dcc3d5354de4ec53fb5602f3e40adbfe1a1156b1d3fdf81cbf01effe12d30f92d7446dc0d1966290c37ff2e24af1a5bd62d5b336ee196c9e2db7763b237445388f0a7fd7df91eb629d5f90edd0554935750de4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dce1a4f575a8fa548e2452ae5b84ddc41bc8659048474b4cb9f276c6c797b17d1ca42067ac5eeacafc76b00da8d958291ca8d47e41bb4ccea2227444a6855c1925551bc2f2cc2fda7674392f39d2944dc8cf6033;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafabfcf1abd5029822c91b7e571a584479e568b283937867f35680efa554024efc2758303f6758ad153a047c3c650ee696f58ef25cf0cac801fb92ade61c4d01d615de87fabe1f5d7050c9260acf96cefdd5c5888;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4e6901a90bb2a1c9a320e8106f7c72083e9c2977043492874484f582aa928a43b0db77eaec53a0124bfc212544808c77bb3606b167c5e36a4baa11363d700e3c63235e08d94d2a880aa31895accdf65d83eb2c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18ecc98fbe666a98697500ac78ad4e2fcd101e0084654f10c6b8a002ca7f4b463d53929f129d246f208b1f6aef24907998226067be0db0495cd11cae516eeae7a6a06ac2a68aca146d0710d006c5890b1fc7dcf75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7b9383ec27a29746f48564759b0374b3459c354c421e0fa1a7b87fbc24b5ce22472d618fd97254ca442a977e3c869051726ba4dc7ec9f1575b7b079ee4c0c62dec1a12c4ab09623a3ce623907c6a569bc7a1d9d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he44299800ebe95093777be33922f906a54d08429dc4cdbd81095128392394ad94aa0c9bd56a3b58eaeceb001a6b180aea8bd5f964e17433432b1517b293c364813655a489c42879096e21ce97ffb07d6604739c8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bd3c0b97b7547201db3f6e685893541bab74e160b222d7b9dcc93bbc65e8c264327b98a8fb03c406164b7fde6adcd0bff5d4dab40b0be7a6c6e35cf2f7ec7a12430ca77301f21ef3ffff17ab60ce2bb874583e73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd04314befaf501d1ab78fbc71ef5d1bb028c6d784e305b9b9cf1041fa08e177289bbc0c3ae0115505b8c6cc8b04137c8b4855b50953902b5973ed3fa03f7afc5c36bc0ea6e1cf3963bc2f1ede499a5852addff19f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c49b97f9c7eee33e4374791b5a4b869134141a96a2f757afa1eb9aecb37e1e349c089c02ef035af2c537a53a9d0e31a44ef3523488a170cb03a3602b28db2360c7d53c41465421da153e8fe943a58a147c1a6e5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5437fd5f90211fe9a11515cfb8a7a8ff00a04248b95417eacb4f345db5d068ab762336e987abd24461232f572838b725a01ab95c83e630e3ccb08dbdc2d25983b6f54c765bfbca43477a5f33b85759d04111e7d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27a9b1cd01fa3889145c9d540142d7445c51c98698816a31b9c6e82a6120b40fb820ca52598ba57d5adde76ed6b32fe611ee345e050e0e79f3dd5dad7ff68651cd9090ede3163a4a2378221073274bfb72227b5c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7cc452b840da50d71b685004ed8d378091407337cf37ae0208e68e7b2cd062e5c3fcdca78f6e98cbba79ae7cc3876028d55fb73e1c6eff9c4833d3d214b190004ee4bb40e3b750f370b1d4ae1f7ab2b038621e8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fbb348b499693c391b4bc28a9da31e9f2022df70ba6b499706e199a30f7ed20cefb479511280ff903ee6714b07f1fdb0c3924ac7b9394f9740f80bf2feef1edae312d4768d084356ac002e164b9ed9f545f35b4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2832875368f1cbd11c87c88b0dca4d89570946d4561c1dd34270ecedd9ce0f26223b5fbadfdf7e6823349f9926ea0b2aa1fbda3026fc572e01cfab8d34d34e2f6b9a49599e967d6a604d67cb248a6ecfd28e789b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a59d3a9d0e691937ec920893b5326826c436a230d9666c4c64d303b5a24d0ea8d1d0ebbe1367fd715cb209422f02a7a0c09261f56a779e39f1b632e2a63f61b1530f539423161d95a51f38cecd2816ab238a9a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fde284a1b2475126bc360e2911a43cfe57d180d38a624972bc61a9937dbdc027eb2f565c1f3e35918c9edb6c9345b3b22b387118c7c0f39a784d934a774e6189640457ac604e30505892a1e535c5ab3111c4abb7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha15ecc814fcb62fad6af69a720ab7e6b7de04a40ca46d7df1847abfa6602024e4188c73d8a123d9dcffdbf3d281176da607346815cdb215667e3b243dc7a6f77af5006149bc0ed29fbc4f5532b24c6c10170d8fd7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7386f4075375358752711442b534cd14ae0bf6dec5e60b96ffb5e255ead5f08de29ed609de2468790dd506f7f369e3a18f88acbe7f773199cf1ffc3a6e8c465c86831a1539dd880a4e1b5ad80f17c1c864ca03515;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23212908d867b41b43956c3e295aaa8b280d60f10ed9ee19517deb50d90850147a8ab8e675ef970b25f6b2173ac7dbd3cca5a1184a8ae57879c83d5f9e8d3262b9a7e51f05c224c70a5411f74f65e5f32cbd6927c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87ca21da07cc3a20148f463a9661e8de99a4fde5cdc47916368bb56f7174c5bb4f1e5fc853078c83b98cd31c5b545ad66bb1a904d2c4f73c0ad5913fed9a497ae44379e40e84d7c2859a497cc8abf7006d438cc13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde9320362a4b2926cc1c9bfbdc90f4efe3b51aa5224d09d74562233fa3c17315ce331d5a1a4934ca6c6f18d018df607ddf08e3f6e678d53714c22793ca6963809805e2ab9d95effac078fd6a64ca39118d0a0f352;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcba689a6a0a03ffda72d1e1e03dbc629e1b63ba628e0c6700ea6cf454e6bc86454fa07c68a9c83a2c4ad3ed019b711407199e214a131154bc05bc4c1a90b1d0487490a58cfaa68d60a314189566f06a3163e6c87d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbce4f8f79ca8772dc767104abdf06f849dffec393a409de0bc96a2eeb0e81281e79750b67ee5a252dfc4abe4b247604f07d89b54d264dce71ac0e195797907edebe263b3dbf1db5bbc2f6102d6baddb760ecc0a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb89bb218d15950d57006201fe5e165c178d8d3d849af67d9d6a62464a337d12f93715186d16b0187f920f87de66464d86c87637ede4aeac23cf5aac273166b94fd35d0753df4e84925db1b48ad9dd6bba3baadcf3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63f5a1a84bb25102fddd1976c03538826cf45c8f00560dfb646f18c3546f3ab4501e46814f6840ba28ab55922eb196199917ab2ab5c1fb4f54df8df610eaddbe9add6c313c7cc5eecac7570842ad53b0d5b542110;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9194158a1c3f1bfbd998a5a68179d41aba28db4270299fa9f35693a4bf961144ac9efa041662a5b188dcd8e4e3e951c218e6877d4882cc83b85c01ad48f2abdf99fa4212452f35ef8d8594b5fab3d1a5ebaa98dd7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ab49e2c459faac4826b8dff57fe4a126a701c70497bc235d92a82f477905acbcfc5fba83e4da127dc259310f525dc4a6fd4b1733c83af6454505d722226a5730a6f87f87171894e6d93401085bb8e01bc61fefa9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7056cde5ed8ee542fe9bc71799cf096fdcb6fca4ee1459a9b9ee99077f3e17d5e5e9e0fb5cf005e6bd330554593c37c912a15800b228f3babeb0f5b0c3b98a2d482bdf63d6b2f4af6f8be46d8d6f8848d5029784d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6065302dd6e20929237d0fca5f664dc8688b035bff205264252596fe6dc1307476d142a6ce4a8e59d80897a05da831855d5042c7a23a027395440da6a206c68947ebc847fd2f91fb82d4cfde23c0f68ffb035d949;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0cd88e5b630d86bb3a5defdb89fdadb8ed76013936265c4ff71abd7d4c80beaaeb154561ed7923abd9c6f13e75ddb03669b42211fc6cd55a08cb5905048686be79f587d85b5064d521a75e2506ba511f579a9506;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77805ae029626a724920d0b6c31d87b10a34644ec96569db0d67aae0c267aa186b792cad689c0eb08307bf91a00a42de5b4348dbba61f0e064bbf9e5415df6c5090f834cc0f6a9b377e7af4e0430f2e104432e7c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14a06664ab0e25f529be2378405aaeed2569cf2c1be85623af6a9045ef0d5c461891fbdfc5cf3dfe7872c63220778a998ac806084ad840a52bcde1d22968aa4b14d0079e92eb5d453abd5f405f655a2d8742162a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b04846cf1bab2b643bd722522c3aaaf89430bad50369318de48bd5d74ecb7f83aed2382b7c18b2a0b54dff3aed1377c75cf9a20b3aaa5ad32ab25599d148c828d9c4bdbf853bdd4515b5f7abd76a8ead7e752653;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5592683c2106de7b222516b5cbc0fc18886bbdae759f77ef0a323ff06fd69fd69826d18b84a724ae1a698a348b3065b9d2b7109e13721c6a571a2bc17f43ba86d40a6a9470ec5b6398fe5217e2a9a932b7a8e7cae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1da8b022c17166d5695ae135510fc8f84bd2157a24dd021ed720e643b1b29621cef3028ffeadb09097841127f61977d62fa0a881b21e7162a3827ddfd64f4230d72b1906eb64bd0b6faec39f336c756bb54b88dd4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h313115c0022e67fc3a2d51ce88ae23f3c71a82ef61c299652c84b05038c908a424529b45652e33bf6d74e61e642885e881dd0d26321d58e27acc84d22d763d6f1937fd77bd221fedfbfb692c6ad11babb8c2f2334;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2552b2cd00a4e3289bf9478e195b44523ea387ad28ca19411ac80dee3e30310c1401f597d72924080f79035e8c54f123409fb502968368347813f7813a9d39353f15ba9cbb784d5cb82fbda2a77c43fb935b0574d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ab4879ea0aa412e498c5e9e22a5b9b610a33909a04c9ef391e24a77339c7d137cbef0777f243afa7fdccd8b06f248a9210a8567fe10578d607dd5bfe6d7a93a0a6ba1946aef123cbcd5c89d383a2b4ca87fcc206;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f96ddb1dc89f5dc43f4c9f48fc6e076f81450fe975b0b1cee1bd473e0973f9d9ac525d4522fcc5850516bd691f6309779844125398fc0d706c1df4bf899532e0b17ba4644dad5674128b91bce1799fa780ca376d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b793943b04327022b1fae16514799810a3ee72a50a08cccaf929579f75ae197ce875382e732d6227f9b37324c40a39d0f89727be9785606402d66c574406e2f21b059a0cbe0ee7e1ba787fe4fb43e20d1d814d6c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36c2c14e40222cfc85d3136377829ee8b72f6ee72424ad06ca89c7fbf453c69dddff5826fb27f35b73060d2d2d204616083c94aeaa6bd16a109380e6f9c0431d9c2cf09cc3b1b6c6830b8d07ee207b0307b7c4533;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24aa92faef1c56eb5db2e04f7581eb713e78e294d3c52326ca04ca00dee0e6a08bf80fd136fdc0d66be419b5489b779133368307feff54e97fe8331d8a91ecaecba55435f91540a22dc5116130c0a00a4e548ebfb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b3590e04c5fc0dbeb68413296191d799d1276989590717b009dbd89aa4bfe17bd4ddb18303bbddc1f9a96fa67a62ea6a34c949dabe99607c97c21688b8f6262b592e2f936e3937fd0d7744d220dfa131a586d0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdacf98c9295848a8b6dc22e4e80c30f429b5f815db3c23a317b4ef1bd12204d878d869dbc88be53f30d2b50cfa04b45a7a382d489ee7eb79494879b6a825aaa329d79b2538fdfc75233b605b72daf6bd4fb4c698;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef7499f1c3dcc2a4205639caa2235e073f032fe01d37aa5e2405f7b2365a8f6ae94fd8f80e9c8d4086453d630b0d9bf6bb2eadbbda620b8fb3082bc2ddcf13715ff6a6225d6e70f4b2d5677e71930764768eeeba6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha191722e10e2c16a420e8683e46ffdf7b56fe90e1e65085181896c637af4e40d841301149b3c801a542b70fe00d6f35f4bf171fb95f20e1ef16c24a15cb05b6f69604ef1af2d86f05cce6514e699e1cf8c6df2a5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h140eda4b8e30a4aa3361610181a9d6b863209de635f51a824794c4728cdc6bcf06481bf0e6ad0659da7003ab1768629039be023ede533e9d2dbeb35dcf2159508df3e18f6b3f9ef8c6da016dd23058f40af31c333;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed925b06e921660de1224b40d837edb7d143b344b01cde3311d5bd50b00755299e7fb6867d1900d18427d39ca6d3eddda5eb408382c52107457f43384e597713e68dcc8582445065917c359be278284994b268b0e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68c0bf07684714c2cc733b1fa7d0f981b2430da5245294ffaa84253fa9b588d92bbdc992a92f404f249b58a4988edb2ed733ce627377908e1e99482f6d11edce4f7b50be12d72662bf9210faac3e0e5d100cb9c68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c172fc551336450b8bfa004576f9316a1010ac6af25a86e6a5bbacc476ab36d8a91a3b05178c01946a0ab57a4d3efc7214c8c4e8fb7f66b6404405c44aa4449ecc2cb8315e0f7252768736f141b4d73b8cc754c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd3b8650999b37715661c53a6577a2c92d5a04f11de2c09af11df308f4cf9fb3e1e04ab1e4110b88666574fd5397cdbe6dc01059a2793008c67d7ffc42a87d47ba098973f571747dae1fbe92e6523ab7ef9f4beed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc889298b1ed99da03c8432a5ab88c6dda9406f1bd1bfca224a7667a3ab7e2c3adb6a98ae4f9a1935000ee4dd64303305159255a03c36491f2a0d52d1f96e2c408c18ea18b357020e2142a0dc35ce03f5e5e3aac8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36df8ad07d1ec5999ff1161b2edb276913c6e7a2ddb764d0060ec9be26385bb32cd14c5dfc809b290433621b7e1463bf6e02fb745c374cf726607faeba8827e7f2847f81f27e41c7bc89486f20b34a835fbcc2c2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h914cac36b6b4c447cd7a72f4ccfa57e0f891936c1eb64266aed34564c4f80eb00e00c8d5dcb330610008aa9419c863f8cd02e588fbdecdf6777c01880d9d64ec6a5a27ffdfa2c6c4594eec559d0c513caf83cb70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26885506ce15dd787ff2dc2237e98bc5f6d04af64974e8b4a6cd80b18d2723cb58d36813306fbe7e70ebe41792e36f8a2fc90af0cf72c25b36a6825ced5a6de1767199fde584a24293eb225971f68868fd9f2b79e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f385f51e4e9943488a1c40ff402f3731a2da972f7d8a13bc35a41c245fd23c8c74d017ac29ea61cd1cf31dcc0b575b45b6dc878da23a8b6e749788522cc70668d42293bae37fb16fb7722e7e45069deafb258074;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5260b0aaa416396b9b90c7922c9f2f838a21e6744e3685c1c3dc7304cc2d676eb47aabbf475f8bf397454feee5507545d5ace988178c34374138fd54e0430d6e14b1fdedf6429fdcd86e4db1b8f24fb3e435e8cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h425544a223c866bdb99d9f840b33b6854c8a5f862c65fe75f52427b85091c59e7d6fb1b1c5efb8fa8f865a47ae0f6e22ecdd7493953ecd75ff30d0cac0d0721114a63bbfb9d6ebabf50315c274a95cf5b3b51be6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he39b514185e190de3d14eb62a73ed870b53e80affd70a496681c986f5740c975134314ce4f35d0575eb24b69fc245878bc7434f3f7d407a94152ddc66ccfcb7ab47aee6c2c1f54c3c8055e6fa66d25937c9cd52d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80bdb129a750df42ade6fbf978b8768637fcfebd5331cb0fc74f8711ed28f3a2b1804c986eecca78fbb7be856ae5cb833941892656807f71b227cfff045de94bbc9d57ce64bea513bc26d9212df648ea5c1c03f04;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1560c721c51a8c21409d2017be3c25e35384c99501261759cb5c921e1f870b2dd41a05c3c3f2dfaf41eea52791c7439088162e22d9454a5fe033aaeaafafd2cdbf9776e4f7c1023021d8050ee8de6425e55eb7fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h943be6b89e4a200d9a51d9bd3ea4348373b8ca81c93d90d6ba4804faa7ef044d1995cd6ae23f0910e1a8dd6aa3af68ed8248e18b625c17644bf4e28394d041103c1587c4713bbc0b654d9fffea03c72aabe1570ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4265b8cc887b57141984609665433a4f5d7eaac02a9eaec94281061bf4243d399c69a81f1f87efd8cf611bfbd6d45568108b46a014c5fea4a7fd2f09350e88ba7b189ee4f6cca095f125ed6eab85c1d05c596efc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d56e0ac10c7f9da2c8017a1d4efa80304cabee9afd83653acd2a0b69e09711aa8fb22bfb6b7c906f153e8347390b730897b956114a5368cc3011da5cc37725bfb25fc23584d4ee9ca9ab29def1f3419081aa2365;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bdbbd15a0cb951babb410168e3322f0b192c57531bf320f6442cdc6b26a00572455d03bc03d17a5c99b771ed7a7d17a8e055d1b01b1ffb4aba3ce2b79d8cb9e622fcebc5dff5510d89003f6b6098b464afe5c602;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9cfc6022df9e6a3659f4653d9916ddb0a3c6b24a17ae0013ed6305514cd69e3c0184d1b13ebf9fea990804b2b383d2c9bf9b43687455708822b624b0677ff88792f8659ca2a48ef3b2306f9bf895fa05151d2c81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44924d1ab45b9b1ea7af8a79afb08555ce20e860707ab4352b5c6099a6efd8d535ec145d61962fb37ea1dd4ce62cee48516778d2624c5de66c44ee9ccd98a7c6bfcb83473dbaee92004e02d9a67a3cc9daa68f61;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha822cf87ad4834f681c72ccc2c549b0a68a18bc9ad32995177fae362cb0b859a5c5bef6230b13cbc17b983f31b9b5c0c2190ce12bc751a3fe65e22641c2a837022ee1b6171b5e7ff59e959f1768c2f51f618d3ff2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37110e569de1ff43d9d560800ff4cd652c3b1952f2feb096c5cc229d065ce552f94b55da20db844404735b936e2a2d052d80ce8d89e706607e73b9df8c711b71e250c4a07476ef6c228fc1b96008fe2440dc6f775;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce12072a9e577b5efb6dd930d25c513673544d367ba4664cc997b6370d8411d6ce0ffb4cc9121fe5bcfe2c067a44ab425bf8727ed4c60b34ac1de1e4c7f6c4c379ac5fcb21f1b62e740215c9bb748cbee5fb97e5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26e7ad3475d9cac2f8225794747df13bff9815cc99ee3e7106caa7e65a3fe705ca2704cec3ea437b3b81f6ae6c862fdda32985bf9c7e9ece1853f6475123b9abb6a53ac4ca68a84628e2f2c08682b9d00bf4a958e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d2d30f1dcdec7b35bcc1b5ea080a6fcaa523f785a5e3ea1902af840951812992f4b453eea8a1c7683651b08f61fdd5d4058aad1b3dbc7fe5abc67835631303a27ba6988c146794c2fbf0968ddafe79e1a809f49e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf07dbf47a0b199bb41b9a04c5434d753c1e714f048ca024b3b80e1a30eb3260007ff2402fe64f4194382646b4190868a07c89e5a220ae354886412b00c5761beeb78fac4bb31f17f1d6ed339724e44a05e5483569;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb63f55032f04dd664ae50f5a6ccc3e5eea2866affc276f77bb8a12d635ab4a22e4474bd26d30ea0fc70c916ed9de237dcb6d117d4946b8c5e077240c5720479dfbd637a51c44344a091afb3e972bc40a75654842a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87055a15115dee9804d4c9a7c7be6a42b3f8e1dd0344664df0ae58057493c501908328ebf0829c26f90e16f3f0cfdff728be2374831ad145f3988d55188b3d9b7da172fc6c1d9a7cf728a636ebac7be38db85ad32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9daacdf75fa61a31ab008080dcc75d43c29ebc447961d8ff98ed5d6e098157f2e5231f3605956694efe25e71a21368ac1e704938db0b94b435c968e34f08835c20f53dce2c810d1d7f661fcf709850e4c75f7819;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd53b8b5534e84ca6d1a6073ad3d1d0876396551743132c6c4501a8a11097173dc3164d889f78cebf428653bbcaf73397c08316004190b777d6c08970f409d0961c647bac41ecdc467b1bc9d25758a352453f5776c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b9fe5020bdf80895338bd245833c9a023057061491786396c526faa6200933b6f367296a19bdbdb45dbc5fa894c23b28ea8602f3f237a38d49b66f05d6f202fb16b6c22c06420c84f3e6aa6f258ab8241a43f4c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14593c1d85e48a67817b25babfbb6f424580a54ca8030f194fdce2ff49fb8966a790f8430ccd8f763aea36678f6edbf660d6970bd797efbfc949a2a1fd9c182314e733240338b18d1e1ae6a7c8a8744a05b0d55c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4638aebd271f4c516f3902c052bc22c8638bd972e4e5595945b754109d72784606a9d9db8086d04bc52dd8dc3cbb256d8c7a7b1accafa95bda321199bc413da62ac5ab1ebe7da242e0af211ffa674482c2741c2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d57dbc8617c8f7ff21e379548ac8980983bd9b88e09fe36276c80b7c0b76962459c5e44b56f2ab665a9fc3f092663b65065499a18dee2964c93cfaff7e1bef00ea2c6e0fe9688f7ef09aec532279ecd84c5860bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9594a82fe993ed78ff4cd9de3735841af8ca30aded6236bc38aa2e6d9620bebfc5ebb6ccbca9a11a21e9eee74655eef3c9e66db1b8f5897a79e3ade9ec2943ab65d5fe4281567056f4a730fa6846dbcc89b57be07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96a89e63e0fba17f5776ae7568fe83973148a104e3d57efbe15b18e2d8d0f6e1570c0ab5e20f29b52c619de56cae33b7f58f66cbd1d9fa1a6b1bac6875bd6faf83d349d2a24658ad33890154530a5a9f19199ca55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h611ed5af821a951f995c72d437736edd249933969ea39f188136c186b4cb07e42e0004b5c9807c7720682cba0c2af4eaace68d24eec91cc95d02bfff3fced93dd609b847f9639647788a87ca429e22eaee5da15fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96c1b2551dd5de0e2d26080d39da8b3d178168c289934d5e4a32371e3e1068cef6bb89a506fdc9173bfe46c1f566e3ab56b706807e82284131aec7216cad4f16b333494692d69bc79e46c9d2993e2a098329e4064;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54186c62dc2a24a317ea00feb2b195fc48fac1025667e7eb34c360f3e6429943267d3dbabc7f9e9264d1b23ea636a8277f374611049f7c2e6c50d6a9cc29b9a43d44b28902992a4c993082625721b5f3737edc950;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h752b1bb833477489b7f07ff465fd097200f4fa401188516ddb5be46227ff8ed757d03f237f1c1012c3805c4af6ec1bde0340ddaf4c79a159bf9cfefbaf064eaf672844fa087f0ddb2e8ad157a30433eee92256c7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d714dbea2a6b25b0f831061e4befc1b218260875a11adfad91bc1fd67ed92fd74583b5910a0d50e331e46d8267f4c3c701317f618166bccc448158396b89dfa773dc0014224dfc391c7ec97e6e12658c5f0d9bc8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64eef255620165c2ebd1578e81168246aaddf2e157994faee98adf886609ac4669f88072e9ede195b40062a0ccc2097cfef2888fe8133b94bc68a6fd7ebbe321ef7ad19f62c60ca34b90277754fc34813d4204f59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9f89cb414b4a8d18d97a9ba8c8f115557c1ea36b9d4b63a5c7b125006e0a4ae397370ae300ab9d5e9c79cd77c26e935f794b1fc5d5ba29efcdfe430e4ab4512e584e7d719c86faebd2aa154e33a610292652d289;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7de7760a484cd1b86ede5c258d63568282973e24367064021eff652e956ea51ae35f81b92d862c3b799d59deb2dc06d9ca68ae0b30ac71552b42bb0837ffb45800a78eb31dba7dc6de838c46fd7679c7ecbb86f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h345603b13f8bd8d30a7f58f237b81d09539c00970690d7cb00c4d2778c9f084f382f6fe38158733c3f59b55c294130270b7dacfe2ba7c46aade990826781df9486e26debe99081dd6850813d5f750ce40b861f6cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h503914fc63670abb37454a0b583dc84b697a72f34aa086a63de99be70372c89b072e25fd348d41009eb65af7bd56907fc043b362e724c5d682c15b06c0068b2ab7836466d9c3a90535cd5ad70cc618755c09e659f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b383f00ab5f27874604c1d19c91b8155ea10e1d90f6b498d3a9e7d6a285a28d3d5511a71f758c4db41cb9748c5f3269f08463a1085d34c7e4f619c3c922d8a2567048fc839f5945e4bbbbdd63d6f0ea20eb26cdc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd304bb23faa5b4aa7afd854369d3b00cef60af403490aa861788b8ff216739e24d8cf19181c3781547407597dcc436d9779eaf47c9014234dfa88c08d4ccfed0ba21727dae82b1cfb81315368051ccb167a9930c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3b949c9d62121af8a172f5ff6e0b02a6f4e4d1a83edd41942e087ed1c44c5cedbd96873742e806bca7b267c1d2a53ab284f4bd0a097c31da8507e73599846283520dedd800d5e580810ef0657ab4f82dcb4c23f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9841e9c2a33c7db0a1d45b56b352a68fe2c3a801a4a0ac527b1563fa036bafd3eeba0b1b5fa391739b333f1f2910700ba5ac2634832d03d7be02c6fcad77ccd67c80b9d6ef0fd687cf8beab3a085b94760f1cde2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2af4b18f6d332c07e4d6f443a0ab1bdcad3c90e5d03866a2b49881bae314d7edcab1dba2a79dd8736ba7d41a7af8e9860528525e8452938553393c9c9aeb838241b2391b3314bf0ddc8304793fc41ec6b6322592e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2eac826277df9d8918512d60b611f4f3e60895615794480788c4c373fe2b353afd6f89c99fd7391304ad03e4d76b4bb015134f1bad348808537c63c26893dd8043fb9f99b7a399ee59244fb66451d105e3b3d2268;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9b3d36de1ae060abdae5b1109100149786e758daa9813090c693225cf341e50f633aebee27a7a98c31c484b496c59cf6de964b48d1430f6cd7696f9fa16beea8c579cfb5f4f3f2379082d97ccacdd8f4ca802a74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdc64b37193d7b2310cd40b846ef32c0f931e6c513a3aa2b195ca2652b4b256692a7d60d9449216a05bbbcb7300fd1218dc304902f1d7c88e63acce0df4babd8e1d91c7a899b5ea56a419a1eebfed9de44d874406;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54b63d88212771bd6d22353697afb745c50e4b67477f416b32e708c53ebc7c406ea54503f94191b15ec2aa2f37abd0fdbeae6e9fa2086d032e494e63f3e7b17d90d39a531bd728ec0d540ceef6662b8d0cf28a180;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc25821a56eb0a0960da37b9124091e85995f225cff26e784417c9de84248d8688b5f0b8e2b0d5d320c3ef76b3ffe54ecd0887323e629c9152c381dbecdc401b33464985b0f45f885f5aef685c468cabf667d91e01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9aee91991059a7ddb418d0b4020112236219b426b467df20e43c41ab0f261d78ad3d5696ce345fa82740073ead0e3fcad210503593e7521614c3ebbdee042686eca1987283ee68007fc645a68846a210d3e47a38b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha52ac1912cfc7333083ec4147f5b1f36d14760ef2aa1bb3c72556ed0fba8d8d3509f851ec2ed3d7f0fafaed9639080d2e95783a81a2a434bedcc4c5bcd645f280fb4b53942ecb92601529009deee523d5d52d9e16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95a356f22117f3947b9b93f3be7d508442249d048a20582ba157f7569c72fab42d019b45fb2f5c4e7bf95323b6c886c4799c92678a674d78cb4595a4f5ba75452dbde5a4d434e66051fe38baa988d57f57979bc6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bc34c70f27206554ba4087d8783e0900553bca7679b01537d51c451945e348ce45cc982c399f8d6f8b6c0cb56ca454b7bebd407092f518c67dd552b875a8783ebfc684d07b36e778cc36d06ef02b797ff6e7acad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4608bc9e69fd39cf411e746ba90f255b13f0ca2bd1e7ac7d57f1102fcb2756452f6482feeab3a5161431fdb72eb6d293fa9e7286cecdff84c8d8f0464fd2888064981779c2dbe08055aa1839343aec58e7d44edc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf75507aac4b35ae75a0fff39eea3ed99ef8f2c85517f96e22e83c4009cd1a80baec5c2355a7adc92c037251b7764e87e09d6f72ae45d829d46c19a0b969d5f6df463f62b447aab8098d70c4079b686facfb6ceab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73c1e17e25fe27b7f3a91e5794756e93db3b59644dc193d4e4905be2fe0b9e43ba339568b1f4ea53b69ae2f6c7ddf181bf8dda7ca2343a026d98ee056e1b52f298afe3836c39e78a612f5e59c8e75acf2f43c0a41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97bab2a920e435bf9c7dcdb56fd44eaa306a35737cb7060ae5c36da39ed2a28182d13d21ca334e1d8bb4828e0855bbd3ae16fe853930839ec266bbecdccb54480681fd1c5bf571e6d513fcc706f9745103d203258;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd00ee9a6bdddb81c443796c8a9d77aae23190f8199ad6685883f7c2eb0bb79461c1f281e21a031a836b47de2ac6ddb834d5fd7acbccc91cc4d633f32653b5e9836cc67e9c5da974111af8392b913ef03bca66bc4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68a50b200ef7d9a0843d8580998330172bdf0a5e55cbde60384f2254cfb3d3839ef308e73c3160d028d332694b8656829e6ec9fd1eada3bd894274c4b5b36229f307aadfe834645a72a0afcf7b7e51390d0379172;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb44ec0e8bc821b438a05a7a4891a2a7c4910b9fa9392fe7bd7b7040a3cf4785e262af92d108744d68f98f77937f68d9faba93f06ff400c64fb58bb468e81590f0471d35b9132d567254316a3971a6fff47cf0aae1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfdb78c9b7fa88d7f4319142c666d3aa78aa65bdb51459bab689ab4eeab71860ec4d375f6195a935b3158d5a2ecbfc42d4e1fbbd9f1fed894a68ea9474473af53334b8d3cd04cff76c0032f326045096afb5e83f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50e9f3d91f2113f8ce4b426c8785504f6488a068fc4c5d0ab80cfe48e4ec70d6b17fe9fc390a18905c049759a43e974776f5ea68b0b7b2d1552ce3f5c97e1260411a1333478c06f5cdd0c4f18f6c32768ccb1b1de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d24f47d2e82e872f3815c2b9d7a41ebe735390d57e63bae04fd15e0060a5917bc2bd464460768c8168bceaabfebf4e5cbe7510a4c9cf08c31405585d7f799474f456b08918930acf097a98bfa9c9b95275caff0e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd21e35cd415dd3f2300993f7b5cf3d303338b22b3bb107c25b601d426e1bdb2c7118a73dede291bce8677bb69c82d81d80899cfd76f947b99d51056fd1c01232148c1698275423cfd8aae8999e308895924b75d33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f662c251eb0f5140f8b98c4cb97243260bcf1e3b78ae6e8b58375a4d6907b7c7117e49850435cb37e1f17ef45a9285d92ae8f7eaa519a55c64d60faa3d5da328be97c72d447a973b4f7bd1a9aadddc967c03103a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9d870d878183c92715ef244547423cd44622dd25b84c74d64770ab672c624a28a79835698afd390deb346bd0e65d33cb70b8e975235029c0705fb175d51941db4799321e0090c41714fa44897185412109bde73e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf73b70256709f88bd1912db2e6b8ee45402b7d12643d7e3534b519dbb690fbced7619844978e4704df50456dcbe1d0b5be6591fddb6bf7588ecd04dd13127a87874e67bdeabe7bc6e115cc50cb9eea52f37c8a887;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5cf6b17ef3393e18a26711624b29fcf776c4f8ddd490312d3571d2bbb2b51759fb0b579d6ce2770c609517e85c7f053aaaea426435bdf510230f736e70aeace198445d4a0f8e63bffa621837c805b53c84c929c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafa29943a2b8b7114551aa23489f30185c22ac9a87fe90867541b779e628f4faf186298c04358f4d8f6ccc124dfe5781c7141e13f7f3e9a43b191022da5029a135200c1c53e05354dab34c756f39c336a8e000bfd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3ec677f1b31a78c74c69c3e6ab441b995b5dbb2a4a1ae123f375d88dcb49df56cf2c0cc45a31ef88122ae7ac34ade8879e00d276c3110cd918cb7a27097b94721e7ea8bdc0c5fa678d63a49e9a3fb6c142b6b284;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba695a5156c3d418801a406ecec48cd4fea8cf0534c18e64c431b30a90bdd638dd2ef9712fd008c07c18edc6fb156f298070d9f71ea66fe216d1cd6131031b76e9b44d0d29325f243702dddbe09b9c0d0787b3e5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc12d0c52bdc1f33fcbf68ee5067a03bffcdea1bee45a94180ec654a0e3c7985edd37a0a13d4588cd89ab9bc63cca46af64005442575833fda74d26517af946cc54e61e1e3d92c886cca41eeff210b031f5091a3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d8dcf3216747c728bcd770937c66136a4acbd6ed3213be1e3111ea032c05cd01bd7de96a4a8c0cba99beefb7291b7b806c2c340546d59a09559d824da889d13df1a55c0dcc83e301f18a9df169608a3b3828193f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cfe9145b6853d9267c1e7b8e9ac42adddcae419ea7eebad2115be1f47426e56a0a48643cad0d8432981221142cd2184a809c1f4997a71e941e7dcb752c434adadf5b062dcb5ebfde1ffcef44cea66aa5695da8f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e8321cc24fbba283110e943331b341404854f8464b617690adf02bd31f3ee8c912a048265aa3b48ebb88f0d46f3904d8d8e9cd4a5ce9ff34aac9fb2b6c43c41617bf4e7517d32adb9691144cde241c98af44251b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb6ff5380ced442ca9851343e4446e004d5e8b0a031c5fc9c7f597e17d25e6402004f4e30cc9353a002d5e3c6cbbd72c4908c576e3bee380481a084ba84f59906c51052c6c9a1977363f2b8892512a4e4908397e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98f8dd430251888a30c2d67c4807712f5ba10bf6bdb56920b50db3cd7047b0cba93a3a1fc0ad82d84dbad9c6493532af7a14486ddc4ec3021ba477615b34dc380b8f815f57495a2a1707322768a5d8c04d8151527;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc42a572e84ce008ab85a23f83c61f3ebd0b441c3e642371119f73b7661c35efb94072b570625780796991966942aa4ec033514f5e02527e5e714b92d5377516a15687c65125e5617179a7f623ed26a67aefb0d343;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1da8a38386fcc8065cb366e33ad8ddf873eec3ad9ac7a04172420654afd08a07c0e08922b230c8de1029599ef7694d580e05712a0e6b94248e2a34aa805cbc473c523e3308140b3c6c75ba33ca4277ddcad37c8a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b98419059198d5eebef32d45bca77a6f9d9c9b2090465efdb3b1c82a3fd7e3120634d19f125b8d1b0304ef29dbbd872a456912e54ebe8a394a92cd2a3a8c910c4593bf37a3721b7459c2905f27ab7629c7f63c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89d2d6ac5cfe2de553f3dcc3a7d9b37df25f275e80d70bbbe508dd4c4b22b980e53fe84e7a744a527e1c319425a4b2ebe97616c19454a23b86b87fa76f9fab4f659fd05286a914f5a87adde55f80ef0f6da0a12f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9c57e8d630c1f87f141981b1c32ef368d8e84f0cd8eb1db2051785c46a347a5c221672e16f279345b5c469c3e2a4c64284d88c472e51aea83d486f4392c5ff82d56eb893becb4c62e61b6da1c3f0927da482fb9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b79290251fb8ca5a9e1b156971eeda3bdce7fa3b81493cee5c310ccdc614e8cbbe72f8be24816eb2623e314bb2d44090ebd28b59560509c6d3ce0004e495d60b2f9878504803492e7c36324a5ad0cfee3b633165;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ce2eb7840fd23b63c070ad272f5b998f71c07f0ab2e052aabbf9d8b1ff9cc22717b95d97f61e67c1ff23edd7c63b045a235d9bcd10bf63706b1e0a5a4626c9fec4f290913619a8f8f81066d1c8d2c8f69236454a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f3fd62fda9ce144ef30616f904f25b85cb8af47c753d06b0b2dbe8d3b3556b26f1184eee744bc0ee22a0f13047fe09058c747e279d1d2a4c44b07bbc20133c938667db23993aee5ce4798214da153fbe58c38693;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7430035e5ef12d59b37bdeb9f36e8057456d66d43fe5dbaf24c0e1006da3763807bb039b33b0a2dec0d75fae44b4f50cad51e687578dad81ddee221e1c1aed38843533b92ef286a03de1b69c85249e61a137f1fc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf77685e105047104241c22be603c6c977e6116a70a8565dd48e1291ef1e1c3d6ca59c1dee7be4e8c7d2a32cb27ecc2360766adb4500d9b5d6bd9274629996eebbd3adec3e76ed3ac011951a9ec72066c707b96045;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dcc3bcb18cec60bb06aa3afaf915401b72b7de4db5e6b93e888f6aed462e6d934061c95abcb61ec6c326d53279e7356d6272d129f26b4264dfab39af38722c1e49ebb44e5dfe51900027d9b4450168674a26e467;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bb4b5eb445b4b52f9abc896dec9ff0479d339f4f72f57ee16e6d2eda6effec9e28913002b12d9b8c49e553c873a6ab868d39dc82eaf19a048bf95d071eba9b0ddd2c7682c4ceda0dae30031163500fdb193ee0d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cba7f3b0d870766fa84f134c37673a2de5c5c1df489d223340b404a422b83fc0684bd310c67b81fa92b3714069fccfa6e52565ab305a2b597064020c79d3a699876bdde43e7c821991a75a4e03f769a9fe1472cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7de3a9ac0c5ca4cb5ab7d4dfaad7b5f9e04461e9497cee56e9f573208b2f989472635cffaf72492879e1315497f572ce17f5ad38e1631623bdcc05607117bd1aa9228541606b8b5d150f55243b6b709790d350b63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4470511b18ee890b901c6ad561aa91f7e5a2850c1d54c5083e8741eb98c85202c1ec9994cabb3bf1c76bc84163d669617ca40b61604fbb9841588c85eef2f5978aa3d81af944a97be3d661a5d917e6ac4c8398314;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd36448683d7c548f3dce04c38791729409f8485fb94fe6ed8e8cb102fd4cf69b8dd9442951631e0b820522a2f65c76964c1594351b26572e624008d2fd6be828e5cde8ce3ae3f38f7b26baaafa8f25c3c8b88f106;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6101f4990676329f7f19f91291db7504216a1fc8719ad0eecf760e58c0e5db052e6d5871f5316e54ba8fdaf1ece35129077a101117a23c4387684084a0cfcd79d355cdda157ac345cbfd30f036219f5d733fae1d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h312ddc3d256553ad9ec6bcda42362db43996f4a1d5928a9a4089a79a707a456b1255aed11b5040f8b0ec8fc7c54e2fa9051c0307bfa8def5e8ddb9e1a8ce6559e29197c5b3399eb7420abda834ecfaa372dcabdf8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d368048ef85a575ad27303b25b35f9eadd51f309fc888bb12437cb3a2c82b116e7815e3b3b1cfe436e05cb8281ab1643bd494f5a7916c2119229cbb269484120d3d475ab255fb736354f79125ec39e13e7d90743;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f5f1cc4a0c4b3924104eca488ff4a1c8d0ff92a610133b42868126f43d944ec0b9023a312212a43c91205bfaee7bdbc83a4e249c8535f6d2345afd1f4f2eb23296bea00a18f5a9de157a786f4f9af96592859ccf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e39c320118695f9b1d7a81111d7c16387f2d84da063096ccf19f284c28731668dede38205eec7fdd2bac5470d64437e1df79896e6cfbc25d6cf54a21c6b8e0d6f8e95acbc14053a1e604815078172ed0d87408b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3aba68aebd771dd6f36baf6bb1d22f68cd0376b7b8a33f8ed21edf29b6e04ffb7b6a634f61ab0434daebcaaf2e80caa35ef2f12422be74c6b3ba772a15497777067724ef3738b90b109d652f9155d042a22fb690b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec20c2ac88b8c28257ae026a0b6c93af419dc4109861af3dbcae6af5ca1cc837a6667941a3cd222c28c90633a2cddd16d32a4454fa93114338becc3b1ec404dbbdab272d81eddd297ef9052191e97b65a06d50faf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d7b523c72d12fa4fcbdb480a966e2512bdcf4f4c26fee719b6fcb0ed87de1d06c90dc085e69670e061ff92790eee1cd86fefc56e9769af4fe5f231dfd30eba7cd578e28df55b52fc4ca2c774450023290eb5072b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f3ad69b4d44c95651c03c7e27f6d150fb3250c81380d19cfab6095d33422ce76e6509c311520ab70d508394e8422a2e90a16bbc1622a8c8e1e528abda783dfb2f473862df7014797a7d665cd35e4da1eb5846521;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bab8736a1042e25bbf7410cb87e31216963a87916629c86dc89d39e99d3169b2889ecd29de77393b0806aef9b89810d1045896b2870d951e660fec77a205338e1eda92ce800fa3271527fddce48e7b63476b8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h894b9b50571919dda9d3ee8e48975b56e1b33670f7b4e79c55d94d41438b603f834a581f973dadd0f4f200e75c112d2970e5e42fc1cc1eb17ec7957d3b21a214eef8cb9fcdb477768cce5643ee67fbf04317f845b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he30a00b412a9aaa049cf711f864d3ae4138a368e2b6055c9a65b340ea7534f8f08994cea49b80c51d4259d44e672fb39d63f1020ef469b38d1f96b5ec901aa1caabf1526b2f4ae2e8bb9ec42b51944e3dd5e37b59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55ec07e3d1b3a13678878fd657e3109b2a62aad6810c7ef9cc12a3bf879e2e8d8dd62bd90a2a82b34815a02c5d65a3d3ddc44f38a636335d05570a0dc4e4ef234f305c88bebddfdc465240e77c1096faa65705e37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5433177c8fdedc60fc6f0ab97fd5f3d77345713a59cfc8b867404698f67df4c0f273610886dde04a3cdedee67d2128b2eb7796d9471fb4026948f54d14a553a7221e8afa91e245f7d948bfd396caf341f4a645d42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2474aa3e607cdc2b46db381178eab1c6da2aa2c25c3f5f32632f940885b1bdb339a0968b64b4f4acf5e9a775aa853b2936273e06f355750242f00db3ae09ad666de3641ff4cb9e483e4d49f1d38e718e1857b4c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he611139a8d5d4b2b269b2dbef2c2a9f341d1ba51c306177c08895ec76f607170e7575d29e116670b2f35f18ae3e134281aa3780706543c8f17ddcf5446cbec58e8312b99846438888cae2c0f3b12b9460ade82661;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65e6bb98f3c14804088f815b1a7a20a0295a241c106a87f0cc56c48ff30a04f2319a501aa23a7cced6faf6c23619aec20bf1bd43c293de5a7007cfa6ae67485a770fe087ba77eff14a39bffd78b003f4190779dd2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15df94c6e23e77285031b2dc3dd29345972d8d490fa428f3c6b81127bfa2390f2a6d89080a6291971c30815801b5632333eeb9daf4bae41e48aaed780d9e430196f2a4569dd957c200d569babb9051d06c4813c08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aeeab00adcabce3a9ad2a8b85c7455a81e52938b42ab5f96d96ae0f369b6f787a3852dd6028a7916ef864d741e99f748349f7a81a27f5b4b9c9a406e699ea94a0ba0d3af3bbd33ae513d07df8d8706ac06711774;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf6f27c8e791023d1403d6da68ab6de6658a864f68101d3b0f649ed993ad072cdb6b5ceca603dba84e97164af118bcaf6c8db6ff7b2a6e8716586d1d349edaf123ce6fb66c8a0ffa9d63f3ffd28cee2bcb9faa5e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d1972b021d965043921b6c1807d904b7f76c3f122064bb2a6b350adcb5821284eb59d4770d33dd029fe065cc2529fd90b469c2771d85471b194a4d21c7239e389472cc4202861bc279257e7b1abf866c37e2cd5f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1536aa1025c9219cbf7ed73fa9aa139bcfc918ea411cdff77fe86038f069b8fc3144a3c97a3227b6b8c9851395c55d5abd801b5b57238ac9b5eabb8bcb651b9eea871f7371d8eb72001d340151c0d7498caf274d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cd5319cdb527c9bbee3085d4cc5917872cc5cf9587703ba80bf2431b97f187cdb3679c5f4a280d5c4d4e4aa93e375f2d1980bb2962c9b1839127dcebe43fc0808b62c0b9c7ddf72affdb359b3c9e7a1390610149;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc053ba55079782cedf81ced79fa2d6e555fe4e0faebead32fb2b9e44a0171aac5ae5e1fb3ea7b2db4e6b4fc9a9caf78eb6eb7f0d25fdf3676c8ef4d47479d35967fe062177aeacc0b56d62eb0bc6641d13fd6133;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13d62a31afd809bfc6de17e61a51cc886186c90c51b8b7efd411d83427fb5e65759338ffa4155a496614d590ab2b2cb7c600adf78a83551af580f8a19a2fd5e62e15073c7c9db761d9616d3ea806dbc718d2b68dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd44d49a4e56baf7abe26958117632f897c0f3a41b84e9ec7e8e8c284adac1377c8feae9daa2d7be2cf59c5521dc95c191f74801badb11a7230f02283826b22afa44d8a382a55d4f7a5b53b82fc10200db2b0043c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2611cfeec94ff71a08193f03b6fe5f4fdd8b167b773ac50c02cc113be48116bff962c76d14cc41e37185f5b19accb07316fa7e6d3b111ad241fb566d7e285a26012cb544a6aa418151e6c9933a6a0e291abf1460e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h709fb0f9d5b2d3f6ab85c9a35ce322366d9362f31949d05250965aebe30387619d3a34a06b6a60884f782c90cee9230cea7f6e61a7bcd46bc04bd404ee4e367f827490cf46074cd98f0a481b1fa66de56dafb14bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f154a1a508a6bbae7c09ff1f565db02a52fbd78800ed10c7300d84f87830d8eee09834c3073b943e99f08cb4891431cce9be64263c598e171fbacd27d12e57ef3eb9a18b084cd376f6ef21cdc7f17308ecc078fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef1d345a60e1e280448f1b4a9646241e033439079617782ec911f6080fee79d964c31a360f3f453313dda599887247ac3d4f82bebea85a535435d5e85dd0311e9314112ee14a4a447b8f2062ba93ce9320c22ff61;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd091ef4e55b7518ea932b65685bea44ea53e49a0c63b68868755f889628a724e556c603d603d073472dfc25f2c5e48db93e1d37598b18a45b0c3079be9637a501857575f2a2f908284934ceab36ecc346acfb6c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d3d62016b961d96ba26f22c46e2fd7b7fe31680964efecc97af897c886f03ba8dcb18913f5d7654f94fc6259defffea61e9c1a3629d66e4c3695e54e3375ca6365c678882218e44b0ab9d574a87b7233d1a0375b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a870045391df68b2c395abbce38fd22a1ca32a5a7e14bc8e0ab201b9f38732f018fcf064eb0a76687bee908845b9dcd8e5daacbdca05ef61606f6ffd927c145f3c2eeeab61b3651a635b59159af710960fe4fa70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd34294c0cc26c0fc21ceb66d6c8248bba65b21bb69361fbb2ac7370d024e466a4721d99412778b9725ddad6397218527d566a70cdf77c8c9c7bb6beb05e52e808e0eaf3e979fa611534c8f8bf6e456cb4d527335;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48e8a7a7e451247ad5eb4fd35e21306f33a131412bbf3d3bd22a638fdabbbe6cd32751a1e49693fc4feee711ef1b58ff9a4f8e79fc7b456374e2ba4e6354c66d0b3bcf77bb5e34caa6ba94db75dfa10252bab2f4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4a5399946c2cdb5cf2fd33f586982960cc023cae6f8b77a130169130189a11bfb8b5eb398359ee09c9a03bb918becf64ff396d956a77da48bcca1fc0389e4441f47f624c60931a5b9529e32ae45d92aa9e8c6e91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19ec2d73501655ac931b6487eb725ce418e8ae8291c3a4f4801b4ec3601bfa8e8f02969ffc3053b71e1941d500ad6fb3a4d522a32f5c534ef5d45094dd4da01fc22cd839cf2c0a7b460c818817c503929273dba33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19239134b9faf6c35a310eb4762afbef9e9df1b97bc6520d2b1c26d65ac2a470386916b217a10d81e1546999bc8cb3271d2cf21df411a8b12dc0268ca5ccd708600bacb863c08af877a1a44b77125f740c45b69e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf346499f23723aff8cd67aaea4807a8f100da153e07c310daf894cc851d0546965cd6caf7a6024f98ab0a672dcd3e8c23eea5ae77751b7454ab5d9f7adcc3be3e26be9724b14ddae798c74b19bcbc41b21e25ce03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a419b5ec807fd35ef01eadcf5af7273a0ba00d7033da3ec52da8d66aa68dbff8d0bcb5a0f9c4458d8206403f0a0259531fedf7fedf0edfc6e0981f1532cf38c3ac845ee55a01a3e996e978d5cde7914d5d129031;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a589c4e112e0a2cc8ac9d634cef66e2625b8286e9c62317eb133500c3671a8ffca195242c20f55df6f9121109f1a14395b155a95bf245bc6de9afbf36d74386d84b4bdd5d67b4ee0d8659b0aada65fd59f07abd7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89eb3f3ed31ea7de8101df6b3ccd40eb80781fc1622b3f3b37e50c1fcc9581be2a3ef0df57582c2804559e6d68e7cfded9d0e4b1e714392070f4dce0f0b744a1a2719357ef7f7f2e206669e7197c5e5c9e2d21afb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf62a7ac43f339ba30aaff37641f6b3832aabc0aa06c4108f81c6c6feb893d78585ab2d851587ed3e02c140366ac1588c45794957f9d08173269878576b044cc4a91223b8370552ab9d3d101a4d7f80e962a275c09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h201e8c2232f343e849773eccecbbc24f47ccc2e0d2bfe6215c1992583dff2f0b4bf78808386b8828a5524e8d7cad701731353dcace77e07091e4fa6e9142c1c6383ad3f346073b4551fdf8c5eb34773cfe068f4fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h914ca3267efa38013216d5ef832b5deaff7e78a6bd2562465414f1b9aa7137291bd75b46f2a6e379a94d7bfa93785fd9bf4e42af8caf068ff25bf8252826159e603e9647fcf593396252279e9a82c8ac15bc8abee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40a8652b035993acc815af21de2948ea78f0bfe410e568028a280aba2743b9b2f0e2cf323216e2247126b66349f211bf577eb0a37ef4fcfe224b1944ccc32485740702b17e9a0aba7614363003abf7865bb91a9a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7df2f1675c3c8e723ccb74c50dce16fc23a3a85795ef1e4202d2c9b4029c2fe50c68bb7ba1bd983bb9e7f5aef96e9f0767fe48fde50c18e6f6a0663b04f249e3637cb11372021634a1306a6c377d61542357222f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf73843b3ffb2553d395c609b96b53968c4d88e61b9962eff696d3ca6efef5f7edc9a0ccbbd0b358cfb0b25ba84be82d554a3f49bb4901cd1ef93c27fa1ecc285c73cc7d4c3a9c9674d601a776088861a01f54ebb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c59ba0e775aa02876061ca412587607f2c91fef8091c9eec98a501336438b3e5f8f5021e6cb945038d9f01578a44ec8134c397ccda5544f15563abf0bb1c1f30f960bc331b87761f437e36a9adcc053d021b8c60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7e4c72b84e568e19863a2d1d4452b7ccad802c03c5347369911f49df7ef8aad2feafbecdb61f1839be3358d51ef9415e627de059a2eca1600f333ff0658080e9b2eaefd65c1d4ad9f0cd47fa83801cb735ea0b29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b40465f1eee995da973a29d47da753d5a4797ca0b48d55fe1466630c640d06d5ecee35617ba92d2b01bd55c9150d75b4299e0bc0d2ed6864f5a23ca827d8905446c27efe33524e16a7c6946f45817b2841415503;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9c3dc03b3b0e8854e0b5892421901b69c241919505a32a991c86150aa65f41e837ba6be839575eb8a119a0900525cd54815606618e069cf201cd7892e76430265aa01236650e9a44904a30eb43f565b50e92dbb0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cf1cc6dd55d4f1b9d42801f3a0943320f7c4f488b6ec282a06d92664ee05501fafba12b25dbc88ba682181989e7cfd95f99d174db81422d4bdc842ddcba496d7d22c63f88a838af8c4de5c2eeec0de10bef65ac0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9751829fad07e457eba41619f225b3b498136b34291d0ac4f307a0a7b7c01fa71a38600e7114d032f6113e0d4528d09ef5ef092f27e1fa7c9e20de2615cd1f6927c093a57588ff9dfea00e9a4783981dae8599e5f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4386e98397614e7a54638f4c49e0317c591be5951577c9332254cdc77dcaa93052b21c07b4069e6279c0060bd668fcb52fd76b9e54598cae0d11df7fbd7d5c7c503e1ea684169f718175f8b8be0bf2fb770e0bb35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc53b80bf36315cd88e785ebf19accf190a0912afbaf7eb47899a0613d3dd16022d4a924726fa6aaf997f7981cd8162acca161d618821130159bb9b5d0ab4b106c249922842425464673ce3c64379ed71dae60501a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5109a707394706452cea2f0bdf11f9a21e4504dff29e3e6e8f2c58b6f19c7b003a11a2850970df4e95d930b2b3f873dd70c84f2fe1f15dc8db048d407d4d113069941c9a5f1fc09796d7e960915c73b4a953af8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57b3977e937b8e24b899ce16a6b0dacc1e733da12e49e7466db6ffa84b04742162ef014a18b73d54366d5a40953dab56d99dafc95d8f87ad9967040d89b62610108f8f017a8a6272034ee1e0144fec7fa1933e6de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68dced5776393ffcabdab477fd906346d24a21e162d045fed1a6ea6ffa11d967ce54be8cd0a0058dd916d0f895057d71dee2d0fd4e595dd990b6b8566baf72d0e0c7bd7fc7d17b8d900dc550716eceb42d1979a8d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1db6d0b32c116db730ad65e98f637216e7e61a92ef44c722a749e18eee35a99e4082b77880cac567e2272294940069f02b446df761e6476df8503d2bd6d2ca18107e6bac6648195b89745eb9482b30bcd92ee959;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1752e5ea9cf84c33bfad411f3e78f8e24585d5a41e43355eaf7163ced481de79190fc6563bd2972984cac60ad6bca8fb6e5045ec9908fc89fb0ee60cbec4816628e019aa599a273681937b639dc0a52ad3b5aa0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h310594a05fe5250eb9f3c066a99028219dfc0a2efc13231c003fd8b65794d0d3c10fa49baf57741e904882b5ecf164747c25f5a665906d79f8000f9a948717f6a8a64869becee76720cb14409ed71b7efe8b6b85b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7b1ca116046fe95d79cc3820bc3cc5f855065e87727d4ae91e697de4f2e1e25923697baea6939336603c46bee09a3b58aaa217549bf48cc3a11be395b8e66b1b9bc8e698086599217609cd824dd5d7fee9e1b6ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b48939ce97daea75ca202d8381a928db04689ba5fd9b1749195e21d8165fb18c4b761aa122096dc01cad78ccbdbbfcedd9697692816eab1fd60a12895c4d19c6e0682e8e4f6e60d03fb8d13527b475f32458a1ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h868ddecd9afc44f7015ec53e72254e1e2a31b1769946ec29acd4c877790dced25bd57098b1a5cffcf68b4da722b479a87946bf754a6aaafa41bc22ef94442a40bf5b3178c7b636f4147fbf02f52e9b7ec1c6e9f60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc69d8a7deb0a3119cbd34d8ec08d032fd034629965d7196f3f04a4960ca989ea6b17349ba8246f621a68b1bf64c372e6dbaf3d503f286a6861b22622cf14d6091d63ea9b35cc1a932eade0c15a5e9a4295acfc252;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae5680ce764829f3eaa212367b57d2354fd2c174f0b97bcc9f4a9e7153cf0de607444f0a85e2a3b2ae697ea05a2d62a61d178abf08c6b9e8ed504416a72fa15d2e00779ac4f26f29ef5a9afd018f3030dc95c2447;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41154e170428c64e4996a79befb07b3dc92114fc1e170c41d8f0beaa0eec4a3d203e35a73b33f4d2a2dcf14f74fbe06eb998eac9b20768da99888d24ba16d23f0153f5846e6abced9d837da38c7ddef2f70a38892;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba662d83cef7b00498de400935a1b8300eceb606070499194772012e6133eb91db2ab822050314af0ffb45d4ffabb991146dbc0ca689eca95418c8449e80e9ce2fff3f6c19a8972689d49c622a37a789cf71a585;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2766ebad86ddfe1ba44528fd088587f00491648685b3ef0b20e2b6779ad1ca34fba28aca57e604f3413d1e2752c65ed44fa5af769ea79dd58487186b4d2940e4fc16e275b133e9af123f2acd7c03c193c1bd6e9d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha396216a1741dd9a536c6546f044e9b3c1661fd83eb33ddf3bb1c2fa93433d39f85e5396c762cafbdf52ec008b9e7a7386413ea29f97b4bfbe6e24c035ff2d7ffba8f921df5ddf48e46bc0a9ccab21e857a968e2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7efb993fdf831cec4982709713562e58e27073867c2bb3d93215c23fd6b15a57093bfb2de939b979b34f0382538879ac828989fc50174d79545452384cf1d43a72b95f7927df6664a3aeedbcaa9e131b660a1f4dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbab26330d7dd3dbfc906d8a184474e69ddc275a31005eb1cb34fb504216ea6c669957f08e7bee693b044852e6c2010369dafc349a5bef925207d24fac824b81d433f47772b13709b79c96ac90cd07f549242c658;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf986d982b831dd96d4612cd189ca9651ab1854d3ba1f76efe26f251455a89a978ecb47a86fcb42beed8dfce7458a8b08b8f88769904455801103de74221c11fc323ef3fc33907d3f3619a7c5a78b5d7fa55cc2eaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bf9f2f1b3a35b3293aeaf15c19fc92b5e6e244bda75a8cd6df3b00eb4a8d8375caf08b2d3adbb2e718771e8216e78b9d09ba9e033f9fae19c093e724798903f8ccb215bec10488177d363b9e28a7f7b3bf67d89c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha40de119a8c2c261488c5a676c18284e228b95d27eb1dcdf53c3fa3005164dad960403777edd4c9faef7998f0a6687824ed656952ab3ea12c6f571a78da5bc4c89d3973179f81d73fc89dabd30d611f2168e51640;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6e5b36574a9334dd0ff798d05fbcfc90c4cc3a58d59e2d701bfacd9ca24e0dd58a194e0f930c394e75187ba5ef21f462a762ea130a9d7941d8aa064993df25cfd22bd11d21f6b11db22b5e0f93bced329bd108f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h347af0c5a3e36e7fabcf5e184d1f2d2dba7356667f2aae731e2e8dc6b441cb79846693db97082cca44d97b83b75263713e71eaab92787a2e010fa1bc34d4b98bebfa13dc1fe71495f80c01a71e7cd65a9a94235c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb71db36f4f5b3bedbe279edd14f7b4c79bcb0c1cf7702daf50ad43bf7c3b0d45978ca46a64963113ac446c19a45df038055fe1c3523139e45b2a5316c624b2671263b2e92b771282c042713d431a451cdc9d8aa34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h939ace9b7101dc8de01cadc9c53f144545e979279cae90e807995291c63d69403119521cb14b194d99a673fa03043e20d009559f2a8927d876728e1e792f550bc6ed2117d319a613a856a75ff4e474ac7751b4cc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffece7ecb6b8395efb0c77d6de24a3ef1868a1c4a1f0c02447b60ddb27b0f8a1ae91cd80d5994c55876813dd2d1f34fe9ddf3c274c64c70f3583cdb52efc206bcd13da4c0e8cfa3198504b6d709e3087997a2c7fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60d7e8dcbb5c3eef20da6f4b9e4e410a01af9056224f4c0f1b50abf8f8f99ee0e93f990a7ee5cc15fd18967f8943f2055eb5e17d5fb1c79bb42b67df206b33bb9d7abe91e0c1bf22dd3a6afa3c8a2b33ea7bba8d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfda7c240064a06bcaec7cc016cdb7a7d8eee9a667ee1417f7c627f4a4753c147427da5fc41895b6e070067bd687a136ea39ba94d4b307fcfd06381f4c4ab337ea8f5dfd88cfb2a958cb1009e1a7234352300b1447;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcad6284a81241fbd5c45a95f997749fd6071dcd3f1ba7c6e1fa88f0568790aff533079559a09564ae350263ac7421f25e588ac7bd006edb8e7a3623b6cf559cc3bb374e3b9e1bb4d52ccf92c0cec6f89167610290;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedf8fe628cf42f32884de1ce7a4c62670570b74565a882acb8b84dd3c789ea3db60adb2b58c3852c6633a6bb68194e9fa02733948bd6d1819216583d1d81628d508ab997d718300661f18a0f38a8ce3acba689f3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa119de2b71894dedf3914da095832ae2e12bf8c501b0e78316a0d09ae76889ccd5fcdae1666b1beeded3ddac5ca9f5bb6256ba586c117a4e5e8c9302442da24d2688da16ccae5ce5ef7b2cc5459cab30e56086fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he11444649cc9789494f15ef7f914056ed09aec6b545307709f03c50b61d77af5ef0ef9f9b9d439af1889856ec2723213606c6f2cabfbf9e34338d73708bfc6d7dd251e6254d354f1145c859d571db5f5e22fed67c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83fe95d76e142f40939dacb9014cb4c51a64a03f61397b5a6054a85ec622d24cb92cc6a3eda5e12a547336bc50b6b9bd821966b365457715716ad037774bf12ea25f738194d7605f15a625674248a693e0946a6c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a24ce5b86563d8bf4bc98a9d2d3b2242b45036a71dd746c5e27088ae1a3b803e26faaefaafe5672455761c4896e4eae664eaced772d52005faaf96cd068ac38dcd3bead444ae7a65351abb7f019dae675cd1ee4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha81db662a6b68664a91eeff91d79bfa7d91f6467c5fad0c1fbd6e6dd2cb69f85b4414a07b231fe2d4acfd0b855fe3fbb833e3ef9c39186a5186530579a49c35f34e32606df21ab119a33c0397d90f229378270e40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h701f1f5b16c23a46209ffd933191608c7077b24cda13a5c77a268f750212419e1f14c637948d2f9f1e427f682615d809f3e5b9cc8934bcf7ad3bf4dd03e51c2cd84c1611c29b818299961c2ae4e1d468108d19736;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3eb9205b994137f49a14fa83d3700afaa7c5a5317681adb16aa7e5934af085eb8851052227acd9997b16ef6cc349261de8b59c17a993f4f18801a56ce170312d87f75d028515db806d954cc638ecab5eb61aab4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3f1929ba205584c6245191af6027d9a00d7b6e9af2a87a0b0b3ca7f60a9673bcc5d19be767407d6f2cf760437ed7b0acdbc26840358b24c2f45da48a25d64461539e661999cde8406440b9d94cc06c2956729eec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5633ce643741ed53f1d1c26ed732b3d6620e9f4209da4c02d80ce2428d75718f83b5528e8b20e8a2fdaea140eec2d8b85496bebdf6d377a8cb84f6e7331963ca82fcb2048bf4e2f08893a25b3008868916da0d54c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac25bf2d4f2764d6ef4a1f6204b1771113bf43647247afd9179c7fef14d3f7f86e5427fb128fede31381ee59311b7d38cdfe22a5f5808fd504b2abcad32693e9eeb567a97a18776e0408dbf53c1dfa0ebe2245259;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d72e108779f0c19f02d98e10fa76efc46d560941c40aa07f21faf7358e2229c2ece6ba9635130158fc473f1c067e86523aec169c0c47ee554a1b095c177d91c17c3c0e650aab22d41a9fe764b303769304e23742;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d7dca8ccf642c05159326f27b5a357af7c882696fed9a9a8ad859d0c3977ac13e9233ac903c1c6b08adaa3c8e6e0564179093470b5e457d6ffa7ff681e1730566dce46a820e068a05164b241f1075d3508306957;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he97a96b8f57489b239da1f20802c82c705fddd01b02f3d4361f974eae6a8a289fac5389d20d227040242061f337939a2041595575e4122a848e600305d252e931ed59ec8607295ddfa25639c87d912a094f80586b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d5e99578b2e1f5fe9676c29bc07d03abe1d194fccdb1286bc3ed3deb06c619db7206c2bbcc9f1baab37f4973f0a891175ff773d7b8b66a008edff1a8ea8c3a9e20829bb3046fbe4f19748f7d28692c7c80c72771;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43a605b5ceef61b4dca3867f87b15dd542a0baf860879353b4ee2b78511e03f1231d2a791a04ca39f4e565b6ef51b810b6e143e591027109e4320fcca4ee9466f1c550b532c8b37498db08460c43538074e219165;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha61b8e806aea86bbd0d77a80ed6bddf3b72265bd9801a22b4ca122be3283e777d19db80a164e2195a09b9d6628394a3ab89d77956f5839bb073686825279b37d728e33a0d3b1d370359ee8be6fe4f71a7aec3b601;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd15ce9e465bf90e1ad43d8a68083e38614fff489fddfa51423a013ebca03700b25a5d8874ffebbd9bebe00d50e8065bde5b65084960d0ca85741b999cf3bf73b1ea2e166e7d0a4053ee56e91caca76ac628f3c0fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb499a47fc611052ff35e1ad6be0c92064be30ee19460806d0ecde005acc738de787a670395ef5de0b50eb44f8b6aa46853cc8ffc8f0433df5eaa1094f24f24a8f69de17efd5bac9d86768cc133d6a19997f519fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9731201d1506c96f81784cfa07f12b3e801cd99e637a085cb2a1970069f2cb1f58dd9e941aeeb6e0049bb49efd5e941fe38074ce0b96fc5d0b1773da1fcb48a7b549f93aa7ec2f1f8500b3ed68403f51afe56ea70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5d6495d101c046d926344ce29990d765243e7bca35d9803e4f1f1ea634555cdfd00a283fb5eaed83cb1f54de9ef6293353b226546197cc07089a06f0639b65e13075bd3153972a0b07046d2eb7a34f977dea2832;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73f00074e5cf562abf1437460916a76a00b366ff2a9782793e590197e4c8a24cb953b8fa5c5081e63ed6dfd876f0c98aa6481a76baa2b7a908c18c82e67f574836f3df77131f6a7cb98a1bdb84e0da89172df5d82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h861cbf57eedcdef0343a1b570a6210f5a9542600a2426391cdfbaf4affcd093ef3a4f606f30b773e8671942e3f92386014788a280d1a64a8a6ff9c24604728b358832807d6636c0019809752c867452b7e6dbe8ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30221a8dd4f23d2ad244138131ca06c3d83bb1b84c439ac7292a6f061da56bddf4b850a06409b351400c4d712c3b1f929ed4cc4bb7ad398751ea6ca0d40449e4b154058c352cb16b070c1d1b49608a53f41c2b2d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc06f79608920d1993c77ab4971abbb9c0bb30a2d8b457efdbd310fcf6ac5ca1c101013de6eca9e4e31b34589e62ae020f548c34540ff3c4af1ce2beeed3ce6cf2fe20ffcec8bc6ee8bd250b9ff8c0368636d1536;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf636ac76ce8c9bab71ea6c6a257915e0b9c682ce30992f615364387130b9fb5acfbd8f9940ade452eced89073e4fe34e0e006a66511efd449d54a59c04b3bba2496f76da5f2c2a56cb2cf11a2a250c09a51e8df8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3353107199eccd5a464a5e1bd8d225945f93261487856dd38f0c99c488d6e8f4de258912ea21a466af221563db0adde272c8329d2760ac7c41475e333bf6304ed445b63f79669f555656ce3a2f95e1ae613a30664;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6c9b8582ebbca208b7dc2eac40d30f6180f782446419aa3efd5a8d0024ed249fbaab6fd9185121aa5997002b78c051f19b164bc2739cff2300b39c5cb8b3e9e435baec52fdb8ebe4343d8fd6aa84a9d316747b3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc15aad2963686d617dec854c60825591de5b23e616b53cec646d9ad2e8fe9ee2ed95f1d73130c0f2be6c13708a6ad0dd08ef1756d35901b70726b9b2fc61c84761d708d420d7455cdd5e7c69daa4b3915d8b3183c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13725ffb780b2ebfc077cb7c9b405b6795ec8f50bdba61a2a88197dbf173fca9568ed9832c09eef9ca25d17be9d3e08d85b97efa72df118bc02b14dc00e644f2aff2b7138e0227b16f8a06d044dd638b90eceb3dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4b727b1f65f6a1a0a1a754dbd3d2330453b9a868b22596a7db259c6c0f53f93a6eda610a5379c4849ae11e0f11e03887c4e93beee1b2242ff20ab04ec073b448da0e9a7ec3e786c9c90fdc24a3c4b08a77bf1b4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcea994ca2dfe7db0cde717525cef6bc02a2bd9c45c259ae6aa38c0f949d81dbc8d1b5205d1d41eec148429428d8dafc0bc2b3fcdc05d058aa2ebe37d8bfc428537cbf5353e9b0f57f7de14433e58abff8e4a1f83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ef1bad59eeafa4d46e71ffc2a37f8c2ae65f1cc3301575ddb0c25ad836866eeb45b5f0983581540c1d194b842d823d3195946968f5fb66771f4493ba92d4cd5038fa7f982e5acb34ba26bded9f9ad45f27bb8c8f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41bc99c1586f72d6c2ef2672ddb1ccc78e416dd468781dcfe2a54cb98cf10bb5be7510ae84f0fbafe7f162eddc1ac20eada5d20abe9201ee791f2cf5d404c7c1fcff28e73f86fa635f0778d4a612b3fc52ba6e07a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1098c0ba43f68118023b10308bb549e4a938c9b81f86bb768003a355d440fdce6b01dd94980949328abc7ba24dffa6e6ddbfa3dc83714072c40a6205910ca6c50e10066d5c9a2a7993e31136f804c8d5cad5f7811;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1f83befa445f05422f74a9611558e2ceb19d2b9d3f1612d058aa1bbc77f4837f5ab7eb25a61123c3881c3d1c001d9b0287a564674baaf55626439861892a7a2125b26934d257d19a1962e54c78948f86a3a7ec38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ecd60bf42018046620275f1397a10479a9e5e42ee9be0ed2e99ac885a19893d3ca65f6ef72f8196186a0cde4d986c439120e3c6b0544f13fee8cecbb8acec34ab0b42bf8cad9fc9cd919f9d6b153580327b3c6db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he987b1c66a04b49fc6e7cbbcd85370c771d86691d06a7434e51fdfc4289c92177488b35e4282d536037d039a775b3827edc3e3dda12fe9525e36d55df7a9c3852eeacf81fd024091dff65876ad7c2ab6f2e977aab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc87c9bf2e9a649bb20b8434104d7c9f30ba9259f1d1f7936f214ee1f377fd52c2239aecfce860d7010e87e09cee443ee3ee3f08b2f35ea42dcc9284efb0a19a6f6946df830c1762bd693dc5b17eb3ccd7fddcf2f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1305efb8dff562e00af40da27aa174a97fb8ddb8c248f6f6bc52b72c330bb464696277723d4bb799b4397ba71a7469191852c81fb3bfdefc5553c4d24f19a9449c27fd1dd735903028e18a37f50abb53bfca6bec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97c5af3bf885601c36f81bbbba4713c5a1287f8a3d82cd4e974caa54fbd573ee56add55842c6ae05dbe89ecd058a0473f5d5bc28528030aeeee9197aa4fc8cec9732341b371492c37d40dad634512e97dd1f028b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe8418a6babee78df1d1ca0871389fc8e4d9f110d219740c74b92d197d43d9d941629d00f0b037bd35811980dc4278f121bf7de232bd74a287c7fe6adfa83f20f5c54f26b1fe0709421fb156025094fa60508fc36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34cf91a747d7f4e0398f9c4b972ee63a0404943a632307a59c912927be4a90b4267dff53879f7795ed6e7370d730e40ebce016e7d3bbedbb408d53fed1702f0e7cd4bae51fa108bcf40fbc41abbdc87e957b5db15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88a8550f07f13441b69955d94c1908bb6d8f813d94b23758826615d4f44db576c367c722ae5e6d402259ec7d8e0635f3b34b137a21bbd4567d9a522ef33452927815dc735442e2cf2d60c45f18785f154fb6c3053;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5da41fb1cb2e2aadfc26437c23d8fa8437ae4a041e290d9188aad7bcf622a0b129d43ff74a2b24df81f0cac00edd9d17adf13a9af4cb07fc1bb847b89c5849f8532c80677671d0b36256e5fd03084a1c1c410edfa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdad9f3a8c47a51271e7b83c31bbbd807a1a2825b8987fc322960b4e2782cf3d204e6c5cb1cb657d70187a456c52cbc96c13687e0a705a3b74181bddf9b1cb80c2b988c336f5e268724ad28df994fa21018c1fbbfd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha23968005a10e5a4823acdb2b35b76494973bd524d3257f3acf712d10cfef4fd2895dc3854c0eaa2cbbd208f8986013ffb2d685ba8df21bac9070edd4d122067cfc712cbb0b5c08abed9e5c5ce434fb4019f429c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc55d573d526b8b46c903d2d2ebd2c70086024e59889e6b580867cbec6c8a2ac95f84fb89a2d75d5159116f287c7106257416054299739a325aa2a9fc29541615ec4c5df078756bf0cc14e58841c6c7e9b09241f56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb6268b115a5f5e08ceb20aa22a22eade45cb2811b896d1c8341e62c20208e386dd2e1c876b912415feac8c9167f0b917eca3a11212f6f332cc225aca17cc0119c93439a401c07749842335c816b497aaebe9e4a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13ddf3b735d5912ff7f9236baa878198ee48eb5fa9a533a8af753a4ae06960f673daa60160be77a46ac638beb1ab307b23979dbe3480f04f1f12b7a2d6fb7364af4968f6a685961da7e02ef425626f1c7aac191c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b8a8ad9abdccfe364288b1c58f28b21ee8297f7679873b342051cc47765e29fa80993653f04c96c1b4655a0ce583150db6c7bc2bcfefbd82dee2f136917b585bd5f7533de807b03562382c65dd953ee664922d8d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeb246ada022adbe9235c7e476d93c26e4b8c0e320de0bea56ff30e5992e6e67ef3f3a180ef1bb5af3a00c43f588766d2422f6b76f2a2c5f7790a1c8590feae0ecaf2c96b7a0d6dfbb718b4a702b1b4cad022c784;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h568cb45d94744884e43b37f14e66cb9b8a293873985dfe2facebfa9961aaecd8bcef8a913b4b98ffe18fb41d63ae549ef24c03f79b057a00ad7ed78a2ad447cb11e2826e4453906776bed00fc0723f9bb6421702b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha31bd760a11f89ce7a63c26ed302667f2e592f2f5ab8e05f2625ef2c2eb9e8d612854990f43922caf6de324d35bfd7f51a04b01ceefb638570643d1c27426ca3e6e147001c9f86de68528aff3c6aca19c4faf1447;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1eff0d7fa088bf4e1fc4f412ca65161383fafac8f26b974770aa529b7dfc6e052750e3efe5a6f6a991ad3cf35e3bf5e311c45eb75b8081a707b2c7addc2b9b2e56c65e70c7aedfb69502faed457c47ab29c9dd143;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91e448f8bcff860f2c8544947804503a8b05f39d6755943af216426a0aa0cc4012f1af35354468bf38f6037cf4914b2619db739437b5a1b2f88442ba8945ecfd144730a0c5c1c5c34bd1144b46394341c9377e857;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb80a1cfa36cb2f7f9f72153781231bf4be882216f0a64672af96168c7e496a9468b307a8ab3674ee25c8da9e1897b0923d591c9d4cb11ecfb374fe8fb312a8f2a897d9a10bee51a145b546639b85feea94c5b6c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b2048dbcfb4935de80330cdd419a3edd14c338ab861de63f66e870397a2411ab47b3672a5721d84370b4b190d7129a21e352c07d3668552455188f8abd64f47ca69c6d57d9c0ba68659542a0f21711a23dda6475;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c51eac9c73912fb0e5015061c7111cac426ef98c4a1ebedad02cce9711fa927b66c633eed66069b8bc122a0b6a5be57c76390842da8aa4350e0ac2f90781c98941217c53b523ff141e8f620b28af5fcca88bc42e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3208eed3ac8b20eb72b6bdaa9c1c7a43db6bed6495e528ca1a6dd0cd07c9d9040674f365c68a38bd81c3280675ed6bde530e4541b100d4f86a759b14eceb04b9e51f8f10fa69a70bd5346e5dfecfa9a10efc72c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e19d00a4116ecd6ac9254e5d1cdeb37a798e7489346c8765b504174f4fdbc6800ac3d3cf24b1f072a350bd63a2c3eeddc9fd7cffe55a2767d5022ad0dc46ca9c037929c251c38ab9fe2ce12b7ca3ef3e29acf6bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha14f1be9c719bd485d5b1db84c7780e4fc02bb1709bc1e2d3f2ea64556fd07a1ec7dcfdd3ae032ff8514ea42eb8e23cb047ddf3076977f721e9b299258bf5cd8b8a5a3647e7aa815d7f9a4c95c1958a9bdbf37acb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3bc73d1e6198a1872957a9015bd2ae2d81e47b2a080e2238573c8e376c66cac163d76c8dd58771517c3928eeaa317bd4ed9ead33558436e27bc8fbec3e9d30bec00ec7d5d4d576eef8e523ecbecbfa116a61a723;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73f811dbb61dd6b353d6cf9cc94cf4c382ff039faa9aeb1a8a2064e185768c43f7bf77f9d5e46cd17d876a20206d8e452e7a0fc4b7712938ec685c3749f5f638c4d66357cab8b5c8bbdbd7b4b871107b26ce1bccb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b5481aaed8a51c9565993e9c9fd0f897dfe74942dd0352654cb853829b3f8ea69b82ca71be36cd18d224339dbb39eb8b62733e1ce30d7626087150593eb486e72e06caccebb14498c253135eecdc45b0f6de0d1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca487d517f93bfe71354b4539fd8ae386773bc7e6277a1675ca5f4adc1183e6b50f5d5e6ce7e011c0fa4d28e3579231ed5ba57eb921c3453edec5fd03b8d54816a2796b5bb37d07a0df66d6e9b4a302576cb46556;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42b7f29f10ee98e5bc15c7788dfab06dd2d669e92c5ec90c9791a06ce35c1256bccf5ea1cc7fb16e119f11edc7b63dd9e899c405934d313d1778938329a2b4640e95b68eb6101cc3b4ec6e7504833dd63669d8a8f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8f40ea825291db23586d7718a916e9b8210e5a52eaa90802dbc3f735dcfcbef6b7580b9fb607613eff6b78f839e669ce44a2228545d5aae01495561f1f1e488715f327ec845a1a94e742d582c3f0d2a4fb998b7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23a8af10db815a0a79b17fb92719b988f9156172a2efbc27110bf811dacd47100c63b3a4e8c3348a27e37c180a93e946c5db9fddd3359ea57ea99e4b862e2566e79850e2da65bec5e5c935086ed241d04b9803517;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a66076139ef8362fb700b1e94923785747fa0fd4d49f4ed7ef69bc0f86d376a79df9af9048f4da0e337f8cea189c15a2a9943621bfb3c4326ec582c24ca7f147478637ccc9aa1001eae1a36dc38b693e40338222;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5517912bc380e69eec5d7a00291c92de0ac64b8dcffc6bd6e4d947085054777e73cd2205269541d24a5285a57cf48143d32bdb31b842428f7dcbe3a466e9fffa4376bfe96cb1eafc66f48432d9a4cbd67fe14ca09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb444559c94f2272d16bd5edb418fc8c4f507c2b3369611e19007bdd96852acc0b8db998e448c99d70dbb6a1df908f699a77bf9f26704e7b26fa096b51ae5541e01591dc0d74f89933cb56b79a576a2ebfcbb2ee6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dcb861e786eb8cfa3150f314a0d10671596537dbef9801bf65c6507757cd94767a43354672963428f0227799fa9fd7f721545d4d8f6e4bed5091b9b02b271e68f69c391ed86b291039361c7d51bc144ab8ef6b05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbad9c46eeabf0db9ab0db494c78ae1399188367827a92bde844abc44762d62c9fcd641d42512abb823e12ff008ffe3bb845cdf5b4e02905236b23038f7fb0c39d27951400c37560f8845d491fed8b7680314fdb69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef1706bd4d3cae62711df92ce33b00a6a1b9d61c4537bd177a79ae2e44c46f4c7e69fefd0e42e6c7cff182fee6883dcd8716f63c81e0842555edf588107efe83ffb055591fbd9dbdfe7d4552815673b59f74ae1f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1c874ba96bdb2b623236703f275d1eda5f1b9f504a773920cbacc79eb82d96ea0a0a74e0ce9df9f383513a3b3fb73f10dd5da700073b4afab002bf83934ae7281245b971bce4deabd5f84426399acddee99a8292;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4ce04dbf130d4a7f4fa1190927194e703266d5e1ab495d6961dfaeaac53cba9c3d7d9e88766036763c614258bc80d443ff300341a03d820c23fdcf50e29aadb046921fa886280ad169a7bfee8321f3647a64794a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59d7da46acd7b1d0b14d7b49ba272f40540555efe027a1ff49eccb823c0e207ccf76a593019d93de68a527889b890a81830e9ac9159cca307dab0a91cef8e11800700c32f32d7edef69bdeed8ec52241f135a36b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca059590202de82878f69a1ffadb13bc4a2e97caf391c304d619ce23c5750a74208d2c26988be8d3c8ef5df7a0d9f8d9cc8cd5fdd9ce524ef5395ba567c580aadf708b285ad49d2ba82fa5f6e992c7d7d1c37ffbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e37c3bf2026beb14e759f52b03d67f12dbeefbf120e75dbb57fcd2c43c80ac3cc0844f080627508bc30b83d6ea13f54bd6aa8511dbe1b0a9bba7bfb94241e8ef72b5656fa2f780d1207694d901070f27a75e6a3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c91155e341bd26f9a6ee765fb27e2755e1a285a046b19e61e31ff9bfe9cc65beaa357ef753afde489e707bb46d7e5fbda93cc7600bbb55697c04b154d0209579aaba441cc5cba930f50a33b69afbacba171fccfb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28eb6a0bc7392205c26c233e7467903e36e765df35d415df2c36f09c36a0985e1aee746b749a4cc6264b55b96ce784951540461598307141cf7e4179d157d0cacf3611cb101b5745e99bc8d550692bbb9be00439e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63a134319c216ad7b63e9a9f4ed149ec59f391e9cfdd98f3ae0abbb0c845b591e61fd9bf340397ac681e7bd466b0ecbab5471577eb547f7a77287d65ace34ea753829b27dbe7078683d5694666124c588a29a96da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7799079dfc58cfa6a48020bd830bf61720fb215e904cc802393c36f26bcabec491e43bea9166587ccb2145c8b4e858d13242b1454abcaa4103acf95f610177f6f6589d3105e2686fcf3213403d4bbb0541331e829;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8887a016664f34b59ee7f514c0b977f0863431af1f151a7b4d21eba8b17b86b370e5df31d287e78978c859edae682e07808f77584ee0d85b26c168aceaac31a53998ed4b6a0b3a47d8b439d10d27152e18d7a4c42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf56726393dc23bdc16add97e2afb356beb47e950109bf9e0462cab8aae6039716d6400a4dc476d1f90a5a381e9240a64cc91bca0f50c127a7abc7773a34cefada18d6a55a9cf4bd5efa2cacc66666cca7642d1efc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cddc82bf41889e04c34fa4ffd91b927dce22c845c06fcbb6c2e4347e61a5f009e9d9ededef263a6bb131ed8b70fd821f23d97bf16401d4562e934edc6e75fbee88332653d235631b269bac75a5988013c941d2f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7482d436079f1baeda1183dfc97ee7f0552cced748754de8b4de03cf7fc9cf538618877fee2128d544fea7bd9ad119ff41557fe27c8b18915dbc463e60f5e1a5317d0ddf9d1bed9e3d917b15f066404bad7ef2df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ab8d72eb6798a11ad781b054ba5a2c3b9f2fc7e45dff1e648ce6bfa40f5597df810fa5670db42851ad40f23582704d6ccbd4b6c856e8abd283cc6093c16086e516f7c91b906445c4ed56fd0115bf8aa9ebbcc50a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16945df59ce7e8914632818ad4e9063becddfa7f0226aeecd08b3fbe573776d831ffc2c3e108afab14ee2181957fc3e1ac08a2a5811a17b940cbba1ab0019798dbac70eb3bca0c31d68b7dfd2ccfeacd0c4e943af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5424c7a65d92441f663a24132f970f274fd62b8f5d23f06890eadc5fdf4f71fa86766e13bc18340403fbef4e1733e1d81bc60afb9d4f480aa5f2f5ac4c79b94daffab90457d82676ae828ad219d19c4ac7dcd5c0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbd0d99186845b61d736c23077bcf7576c3bc41baeef659d69bd7f3b547f2637517e0d19139a4775e5c13acb8041282ee0e02c5de89852e1fe9ee87d2fd3db2bd046b7c278cd4b8be777542ab72f2ff8c7ed53804;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd006637d760de5e0d07e3ab1460048e463c9efd0122fc8916e30b2613a6694c40fce557be4c2e18cc85de8aafc032059dd20dcd3e3b00ba2f5ef9a6a88901478c4a227fe2b8ab2a2648d1ad97aa744eb4f78a3522;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h710ff2775e656d439b6a5a7a68db9c552c13f18462fb288ddbcc85a783b4a68caf663caa58b2ee91212c9172bd3103b22944d6d0f8af321ba840b1ba054117023f6663199520ddb39f0fe8860958d25d2fa406b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h575aad45b4d2f333dd3caa66d9828c9c831d14e3986cf560a3a4b9ea1376b8fa758a76b2d99ff79987cf6c4faabf17b848159a14ea5a449dbc7cb1d8afdad9b5655be26724321e62ec32fc6255c996ba8abc1b423;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc61a545682b45cb860490e80c1c2a75bf0b974a5f61373636665910d78cc201eddc95a4f65fff51c7a703f9f48807df49c29b39f6fef3198380ee88d253aab910c57de2ed197d5e06283ff5735adb5622567be3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18edd047d8bf9bd451f633a23770f512b51e7ba3b8f55a117504d7021b5ce56e7423aea6708819a544971fbacfca313f3dfe73799e9a41204b299bdf66ceab6e4cb17c9408e93d8fd3f8819cb47d2a37641f93c68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f922627b2c28455516194d7e309cd13d1c691ca5d595aa93b5d072e0271a26a3752041c56110ac32c28d94080d1aae1747cf361b3b6a31732aef967f3369bd74e76f968012dba41b9a6cd008b82f9ece5bfed9d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf59f4f94dc4f91dacd7127bae04c105bde35668e72d30eac665eaa561e2356352704431a853f6579b2756c1d3f381acae127d200f5181decf3443338e0cb593c85c100b39f4e9e75b752a714ebf298683f3fb4d17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99ff5a51af521c2c15e6684d286e61460b35e86de4b277c7d2ec79a12e59f102a53f5f8eaa2d8dd241f7a087a47484949018d5ce266ed8b9e6e940a1cde16f0ca83a1548e3bca59bc5e2d35b2bbe33320a1a1f159;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2db149813f1d8f6af27d19f3b9b876bd12ffef74a642f1b35e44599e1c4c68ff9ab4478afa4ca7b0b87bce459801b600f629a6f245d711389bd43c70e2e247af8ab05ed4538764d09d5a8f1db1693d5efd3e875d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3079162261200bf9c182adb1ad22f42288b7b5505f12ca3733cbfc4281a2350d8082dc0bd8e979a1d0d845f7ac3f8eadc4caab5e075c17791ffffd2ccc233c2618c9127392fa0f1aeae95dc66ef24c11d4f10368;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fd7da02bcec0f018c46a2e0cff93c09122152099a97018f70beee352a17ee17874247647eb945581f34e963df9fa28d66d75778c372553e5521d10cd0e03abf16675eaa6a4fa1ae2186d2d5fd5f8260fcf985eaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d99a3deadee45688b9bd4e9c46c55ea060895aa9c4fb32ce9137baf611df043fb0b4cee415be423395176549cc7d09cf41f52948e294177830185e4ef929a32f471bc2f7be7a874e9c83d6bc368e39b0a286b714;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bc5c870d9952afbc37bee4324dec4407e31e805d6af51bb7778e1efbd1267bde3d81e65cb41da1b66ad00ae8db854f403a417076549f2c9dd2d6593f9863bb2e98f544dde294667bd6b7679f6bb7fd527cf1c57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedf0d8a31704465813ee70490d91b389e337a3a3bb1a75aa0f266ef98f498fa5b558f926e9fba22a1c78aa3d496ca6f77506ae746f1aa78c8038542f4c42ee5478f29331ba7d070b3f04aacb247a4f763baffa1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dd2a2abb8211a20e14ddc3b69d20efca7c1b6c5a68ed0fbfe0231fafd07d86fd3be8b42c30ff0fddf9057e8b651b5129f78a9127ef8ab43641accb1bf19b81f24e9b3cc5cfefd396d863aa2bd194e5883ed99bba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0774f8f5825a8ec97a74005d804ee10cab796340dc36dbcef44665494482fd674ceba66d0cec11edb7d20b553f049a8685a09e143c28338fee32a7a0dbb7ce590c7f392a86887993779d80eca94aab2c6bcf1ec1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3872e2e81d22dea460dffed71aea875e1a5476171d3f33cfabfec3260f99b726ed1358a930f214b8f7b2eae11954799048eca2a97ebe763d542b1b0381214241d4821d6bfe59c1b112a7e217724f306e26aa9ceac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf8c740a1e7f1763911cabfea8a92bf810646eb1a4b41ed3a391bf74b95a8f68ed9fd6c6672b3e24b347733fee28c5d6bbe9860fbd155ef923ba02a0f5bbfe3fc42e429c5fb9f18ce7e7f4f4027ab5165a691c6d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0dbaac66ba5159e2d6d0716e043af02632d115962433cc8d7cd4a450b5fc07e698dcfdce1c5c7e8dbe42525fa830c3f9b24e29b654f5837049532982ea327e061a4bfc158b0120d2baa75900b1d34ebf1faae5d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4952db990fd8f85fff799858d087340d17961cfe11dd748e3356567553e349c23ee7dc86270503a1331662a6cd9b07425dc9386709369b1d36bdf06762e00a9d56676feff326780c433596a7ba0327bb0efe0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98ac2570b2d818a3b8bb92cf9389248d4c0f1aca40e44cecb4d144d6c5c93bba0cc811ad78241df8b6a7146088b841fb88a660251ae1fa8f516e1210bc34d199a7a3287fbd822bdc6f0d4d350402b5fde21fdce2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1046ea8dc7b0092233e7d0872d76e4eae0cad258967ecdff25b42186f9971b11571aaaa00dcbe19b0b9058e6f0dab7253ec8245ad56e7c1f923537a33a1e99e6fd1ec24c6334165fe9ba9c68b3aea782757a0b571;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h893a7aa3ae6da04d2ec95546d48cd316e36d6009217d43b23643d36a0ec2efbf41f1b0294a67f4cff24658759814c1bd57ede817c498715bf120e901951e2420d674fdf6b531f86af74f30fcb0969d6c2983b469c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1775ec1b0112ac3e24adfa50761d1b5187000be2e9508c99b3918b8a73f9cd7830fedd53fdf57b8646fcf1bdb981be1271d24a855de7e5b6785d9e54ddd82ddd6f69ac5eb564c26bed63378456c2b6432b5e6102d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce459272473416dd84578d877c05074ef172e63ce7438dfa70c1485d54939509430b6bf64fdb97d467a7eaf51ca21a11d82de8eaf038ed771542b3103509f9762f0644d945b6365d80375e2ce5c7e7d617a24a52c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70dbbc0f7454408c70e1a907e52890d2068befb1cacaf1ced7429e94c07f021a767c68dfb0b1d3fde91160ac4f194ae063320c4612a88c005fa66586a155faa067e8a6bf2d85fa895cfd88f28048442e3a818700e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79666a89735d5fd88669f67cd26716d1972c5ae7f6b47cac5cf95ed46b8dc4afd38d6b6c35e0dd819ebcd17ca28a5771836b8cc21933c6093b39ca167cdd9d96324a46895b33fef3ef73e081345e2bdda9f15e4eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccb0e3e57da6b0b840be9f75570c96af706ae097900ffaee6acbe3ec90abcdf2cc7796d16ffb9e869cf9f9599e4382dcb1bfea20404b177ad2feeb9fe10910c6ff942c9042eb1010ce6f972f4475ee71676389f92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bfe587f812f14e1dfadcb9ab8c05407f4d9f904c6235cc58df554298f69b06e270174a080948a4fca0ed310de5a567b71c4975ca89860995e4643e5cee54b53d5e1b06f0f15aebc6f2949617be276a085f5dd9cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69df916e909735bfaa762fe13efaa3380aeaa861c8ebf352cd7e607fdd1f930743d3e6d0f9021ba1eeee04403cd6769f75a675bc19f0177e66d891d343d969782ff26cc256db911bb34ae8c4482ac3860203eaddd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25db2f28cf6a9f5a5cd003da38fc78ac15c6d12d5d46baf5dfc79499a35d760357dfbfb2f28f73fd3979fd578d08de01b29353141f4b01856327a35b4b29bb0f829db50118c741cb3cf4668cf8717ebd0880a6528;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800c2bc82333ddcf4412e0b669af96ed0a2388e0d0fdb573c7123516f2d2a0a3728ea1a5e7c58778b2a4e8ee744efa893c05b876c0cf923714ce95c58d3e9b962cf8fdcd712f67bc0767b23ce364f992507da640c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2972d216348f1b4da3d7e7f867ed174c15614df14706fa002321524f1ae097fc4545459f39ab0528dedf0e25181c0f646c3ba9336bc122b3fcf16008f123643d246b346a820310d2fc3da2f24b3f9af486c2503d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41209c3b34a488974e65005f6e6b8a6dff00865677dfede7cd0b99b8dcf1aa87fbb2259e490e6ceaad9adb8c43e8a2625d4a60971a88aff9e0fde32748edd29681b062d8adb1acefbb71ea9eb8426bc2f82adb397;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a93b53fb9a7792f49c1986e924f0a1a79b2dd56fa8c238cdffa04ce80cc5bee39be2a8651a053a310a96d944bea5ef341114d2c21e50e3c6b398b6f9db119be68ea4e2f0b754a536f9a2c8a56826f7ba53e38369;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42e7c6a22bf0fffcc6e0af2cb2572cca0d8191b928a4b3fc2f57f133bc76987473b30703decb5226809db5a5f69790a5d70b2fe64f062497590962388f07b0b694d950d71dea5d28f3fd9e372398d19cfbbbdc7ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h140de05f2e00eb27108e7fece0e941e878e8eff7290e43ec1edb1fa2c9fde287317d5422e15f51e9e91d1cffefd2328815e019a7e47f783be1447efe98c5eaa47e7588c06f184e4ef4939f413b7f71a09ae2e6b28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3c483c40a49872c27d2d1006730a091e16eb1ca9e912c8dbc5f71319adae36f9f3b12013858764ce54fd44c4d26ea42cedc51d1dd24c37b165222a1cd99231e3a1e7b3dbe338ef639b8acb9565065b9e2e1ad73c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54d67a721df13fd87e6fda3b7fdb448d1c325f21208bfc16065e15b3bff421ebda12f1a3f4d7d85dcaca673b7c86c6438ae3997bac64e70a52db60703ee88645ee111f6dfb6e9a17b0d0c6dfb7ca6d3d7de25b911;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f5972082a8d6d8fc306bcee0aadd474bb9133856f079e2d6e1ac3849246dfbb37c0180cdc5aba80bd4f19a1182a1b748ed720250ae39bf84a5d82d7354ac7391cd6fd323700087b554ecb68ca72aecb980ca0521;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e15e0c827ab1a8ee7190625d34644906c8de349fabc66f5ff683436dbb2d22d948f7bec84e0f39cf1cb954afbf4f07996d602dc23f99dee264e380b788b375b51ca100a118fa9905e224bc43df4917e7a1179a3f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98df72704a3a46b19cc7a0c66f0ccacd3add3212cf4c59631a23043546a095b345335a95766275710e911e2217a968a0bdba596b644ca2e05786e90921ed3e078690330769ad67dc55390149692d36046ee476161;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc806cbc68e3fd1f61db172510cd8424a345deeead8e3819125f1c458f42cc6532185e4c59c7d6c664cb8f74022307144bcfad6dcf7327dfcb1afaad5b427bc3c1709b87bde9d4979ec1cb5e4603159e939ed0c361;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h933668c3caaf954fbc0190d84a214da6dfd65df2add310f811c8686d8e9c356f112f56e2d487f348500a0268068ba66a8bbd536ff714d5051f123c3ab9c1a79b923e0e6661b2e979175275821e9de7f3ea3c04be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30d88ebaa85592ceeb4c49310889bbdde78a1314cb307fad2788bae7d134dbb4d8c5dfb1a86d2be2555162c2b565fd2905d9d426721f2ca578fb9ae15ac56e070b93a0efed061577519446c5e90a652b395a1c922;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85ef56e9b54985cbc6a4d518b8c216e63a35d160807e6c35ebd2de88b1da736c78d3f67834c6286a8c102dbcb9da3d35f8634ed3cf97d5e58100227586d1f1bab3bdbda02837d1ae0a4f05e108178168a779aef91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbc053950e4efe2690d46ad1db9e835cbb539ceafd69a84c82a6e21d725e0fc168a04ef4bf3f409779aaf086ff47c77085b044b01444508dcb70fa61eb88992eee6c293bcf4a5677ef5c279225e54db6920866a6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2364af2918291c118dd3955923c0dda0f7a6fb59fcf6c6a30a560ca26be1b300d6d25f0e944bf256062982a1575650970624c8af5fd1b284ed70c3fef3f4f94d887c658ec82f8d3fdb66b1decb86bb596dfad4723;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b7a42ae77725ddda10b6e857a76285ef43d71f55040b27979f4c222d5bddcd2426b5c57af7f078ab6d57925e5f7a112304ba8449b580e28dbdeafbef9bf7b02fa4d1738c56c04c8f114dba6f307f8103f63674b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaa25dfa0d884de03a5a8ef2329b593c2e23ee26de15d2ba2c8f610c81938601646201d66a5f499c7522ee39022f4037fc4fd07f98a338660a94256ab63eafd7caf5e12e9eadb014ea8b9cbac738cfd08e5253b2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35c7612efbc41ce3b6cec3e6460da68853052cd811d14f23dd98cab730ddca3cd5d1b442f35dd2b6bef1b79e992cf63fb4c9f79436055ab26d027be417f8315a920c1f939eb8309f22b8009250ed182b7493fd10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h190a71ac14c55a9682785715bcb13f55d2893c658d0661206bbd40493ad340e2c71f098a21957f513451d80b0012157ea903a7629732f5ea883c5bf8c6da4eca454eed051bce9879951beca5cd01ba5b8ba3d081d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9e32524e3005a157e08de77b8a05314667009d3bf838f3179feaacaa811866c0e367e1d189782b5b1475d4c88c41181dc4159e260c66310c02dd13e2976c45340b7a5b9afe87b42184d5fc13a077fe122a200e31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha01ded16371ef6f5f4c33a1d0099b095e4530b34a84466fb3c3e84fa4796c041977c7b6de94415820e33b076ee6f5e321cc90a5f39037a23feb03737ba4b54e4e3bf6bbb3ccb4a717c4a24e83b853b810f63018e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha84b283bad89eb36a8779248f6b80e14057823bb660ea4c9fd73005bb2ea779b5a8e62712db2a48204fc18a873d11c256272ee3f8f0857a72353cbecd4d787d7bc3a0ae97313f3fe71adbaf0a4f48a4420b7043a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf588128fe89b6ff712f0301d5a29835e2fca59b6806ca5fc7e89480fdeea7965df738b4a2a20d9df9cb00cba8515e1eccd9ccab0f99fcdcbcc0eaa2195c2fb8000bb78ce7dcba87f911a9fb306cde60ffe44c800;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0f6af70127d4b22f4368c0d8deb3b42331bc7940827cff15d9e4357db743bd1b9a50f2a815b510c7a15d72d59eca251fc9e5c2ade5ca7f7ed048c8a928e9d679408a0b366833be4e33f30bfde450cf5b47715c3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20f701b90676745057b0baaf44eb654a79e939a3a150f02d5da11325a2a80ef195e770725f772642fa06b8c9aaaea8abc9e7c70ffc51d1be5e9eb10a1eb961d09436d9c10f82df83ee0a77f16ac4885072d51c5b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52cee55aff7ab5eaf83425f90fdde3bd05b4c9b4011259bcc69438f573d685b0bad84c968cca327be9d7add666159d9c971f2548af93a7ec698b4d40be16969b02ba208dee1c7ae2f2511ee29e7fdde86ccf61d30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bf30dc7d49034935447131362042f2ae5c5b361a616e89158d5f24b1cbe6bdd70cf2c5da1c109ed35c7295500dadb6a2f5485b9fc74d478f4dcf55a16a76cee18bb236ab3dede004e9c23afc2d74c0ef9576a525;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f93062dc3de5392326cf072b9dadf2e774657668ce478acb0f59c28bdf14a75d6fb9c3ebb9b4f6b30f9551c6f126a96805d02cef1c4a7523120e974c073a3f1df506ce0c564694b4b0840428f620dc251ab8ad11;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46c286e7922c68656e2d5798d2f9d050abc39fe9ef2487799a5cd018a2dbaed68dfcdb9a9b530831ee618e29f8f23e2ca959f0fea45fa5acc2ec702f7fc311717745860f52768900931400010ee56f07c4e4edd5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9940eb5625e21092769a183213a037153945552eaca2c6310268186844731fd61c26dd3e8223605da41494814566f5acac5999419891589357822c4df4e3174198354f6bea944ae3e13c83b2906a319c930b1fb1e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7db84559daa306cf57ab44f21441dabda01d74e78ea3c869e241e928928b08b7d935859f52eac21d7447f2953efeb5df6660ccd6cb4a2a6d71a5446b2f01d0257cf63b6c166d9b4cd3cc63740fa8e776307ed9efe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5e0d7524c357645c45436a85146fb3fe8e92432ceac374ffdc393e8b769fa2234ddfb171c4505a41ddf1938b21ea32cb3c87d571d586be6b7da41b5864fdbd6c90143784afdc1c48c579f8079e941c5720196bc4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha720d4034ed1ef71f1fe791940214a5d2a679945826dbbad7ebd35dabbb47d30f8b41ebd0dc4c34790f65334206feeb622d0595771d8204c72039ce1ee7a63e81bce778e067063ed2c74e2511c34d373dd5b82988;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h995c7bb5cfc2e7f88c9a78c4ceef1629ab986a30ac55a5f923b4dae0db8db864c2caba9e0cb422fc77deb8fc005b6629423935035a07fefdee5c5aaddedb1c3f66ed01550d618324e74052b6d1c5848231211cdf0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd06a43fdc775d609583fe6396a7537e753ddcf74224a6883470c9f4b7830a05f24efe41bd5231280093602370cfa81816efbefc3c302776500c0314566895dc704597991e0209f37890582634ad291e62f2d9b8db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50f00993116b2b0568cd138ff36e755af8827caded9e674aa7520ecfa810567cb0b39fbdf56da0b501b0a86c820ba5ddc35368eca529f696c2551c7c214b2bbd54d759e48fee1bb494551df5cbbc1654e8ccce6f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h510ecbbf6bedff6c86ae340fd5ed2ddb89ae8c47cb8b55c3b8e5e15b9ae4fea1909f08393a5977ad9b7759bb546c732d64b02fc033498989bc76b9ca3cec4188d73b0fbf062151446a587b8a49806bcb9ab4c08b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he248fb8b09567ddaccd88945510f625a5d73485d8af8506decea2c3c502a79371a1e42e5d618be54928d262bdf029d41506f7e65f0891e893a6b79980eb0c2933d02003207d7a020b34e0f8ec73dfb16d9dec31f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4335ac89e1e22fbc2940f111ce392ebc06b65f664fb367c5035258b6b2c3e4355794185586b7c9bfb0206b4f51261ae8be3b9b843f4958e27bba5b3c3e952aa51e7db9a6b5d6a89857a8dc54c30b4bcce7e69b51e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2591251c2a42c52f4231542a156b3b01288c28e8f58bdc4c20b66cc0bf796495ef04839757fed296baf74786c38ed084797a805366b4aa0135ba19a82eceeaed6e56308840b87c1c949ff68a91c5d2ccb9200e21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfd0767a2b592a3da1c832b3aafb1612160893c8b1e67fbc0db99099d443fa06877c7091119ebae5d5541d81e75c5e51ef875639044ff7d9737e7644e856fd51c80035b0952daaac21ea8b4ef2a81a1eb1e422e5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd68c317e2e9714ad763d493f18f6296f235092b430c29f938bb00407f556161adbcfd101110fe6017e5631b565b43c3e2d1852b59a79271196d041a1a85e350b497bbd119046e83bceeac4ba7731ea1b705f785c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4076d8c5eff4e4318810736f8d9e76eb9f36c153e7bfb72fc98f61a677be23cd4b9a225453591c4151ab8339256f306edad830ec9cc07ca71a263e87779d9d30abe0d0b639f5b85e08af8742d35ff11bf3b3e29fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58878448afd7ceec16d6599d62cb24fde826bf04ddd20e9307ac6e6c43ecf6dd2d41ad01fe93ee44985f8c37dda13efbb98312a5f10fc8902b402b6577bfabe0143843130aa0ddb35ad836494a5aa62478eacc45f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5439c824eace12fc758cc62799150054c0b69c25097b3d43154a17d1ecd97eef0b78ec632b1d9f38f94bca0e82317a1d94104e5e2ed11f21e8081297c66537d5aa40ef54f059c69cfaa2006d32bc783bcaaa3e30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40190e6b71a977bccdc9ef3c596b70f607db4ca86edd75ea8e0a6d31191018f58d311a9a1848c72214495a4dc92a76d272872c0d53ad9a94a4fb1028a8af06e739f2e29982b0a4ca1a63b507cc01ce5bb7ca7620f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3edaa6376f8228dc588c2d39ec9c52a3d6e3b8fdaefc50dfd7b2123409fe75d60e5050f8f5dcf76c43b1bffa7e97ce83c77faed16683f7b35340be297c1b981c17f3a055c317eb7ccb71de1523fa9193ede5a766;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89f35b1f61df1ede418f16d6fdfbe86204c475d53bd7d854d835c94996e1a3f669fa1895758a5d17d5c505cc3766c7496a2d5d9a257eeb310d464ccb2bae9008b243c20d40fc1dd9cb351943b2c79559d7fba4247;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55e57624203f71bc7a624748d54de50c3745f50baf71b531c57ec9d183c1cb53979a60256a24e7f218a99beb8681931decead16e8d402aa3d9d0db0525d37ef43af11beb6875275eb249f8713b8c364c55c246105;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2089313841d30285bc0d9d1d6cf9a2e59491b2056ad2beee4df32a5e6dd26d33bad21bfea51e7ac85d4bfb9a2ef569852ea6c9137d4abf3b5db81efe2e7df3c2c0b70c581e4269b13f48d42879750ff0d85fd88f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d5d79d3a0605b5a54f25ef1074838d61446c75e0ad243243b1729c7225459c4c8c3b5ba6c149b17024c29571baef0892b17f27a352a76e33ac237d5efefe34cce70b258dd0897afe8c4197f68ad8fdfac322449c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0dcea363283f9fa7a352d9597081369bdff51b293f545bd6d422bfc4c8c136c62783b11fa1981a2f680fce2ffb7f62087ce4446226ddf406cfcc6ce69359115e37a6dfefeaaaeaa20e5b1ede0edb26f010698425;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e172bbd112f46b12912025752ca79fc662c6371e6d21b90c1467ce2e54ee5af7b6ee61d0e31d28171d026e8945f218ad0e4294f6d42df7d6d0c7bca8d14f307d91c91dfbec16df2607faf282d095fe849f162ecc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1f4e89c83ad6431c835232bef30be22ddefde79dd139b0f71ea66286d691570ab819f5d5af95cea9db900bea751847fed441c71be1e13a11da70a88536a5a333ee1e0e3e6cdb8516279682424f166a0f2a9b7676;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56fc4cacd8c2bb63594c0b22eb724bf70d11827ac4dd2bc1dda76238e5ca97d6c75d952935194a48bff306827adfa538b061c5f4570035e2fec317e449f0719457d03df1d26368adc5591f8843993248a8c71c2d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5accda87b5dd5884fd8521aeb9b31dc703f026b443b9d7e03f11afd6c3aca7635cab4f2f6b47e192d8f5bb25532011661df7dd7891c3c863fa5ef5295ea7c90e4f0954c497387173a66a50cd851531acce84e992;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ac811015b650268e774212a7094cfa29710c4104b523b83d3033bd15fde28372d845f3a95c23db03494a0fe739c8f0150e85cb5fa6e7d97920af589583e9b0db9034b76f3bc834adfbfb65bda9290cde60edae05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1ba00eefb698e9a6c749c1abf85d124698f3d3343061e01127a70bb6cf735e0264ea5bef7b8c9837a4cf31a1f79d54f97245a579583b06ff599f438dbe7907a553bf713ce38c78f6bc87a7aea325154ca893e6e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6be05afa41cf8c28f0d543ec9fd39a45d3ff655e88361948123d20b77e1d8c7b7f78d420c46995d157b3665c751c049d1f5d0b4fc8393a952088c3a4326d4c94ad97dbcb0f67214a0796da20d4bcb06dd57a2e6de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14c09919188a40294c0fbb816fd5301031217f0bc2323453afe0f88afa4b88d49879c9e7725604fe8c3c1dd01aa6d23273c4fae9b6d454d41c0185da3faa58997626197fd27f7ab614e347a1f537f6d3b396a8e01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaaf5c848206538af51d375e9c2caf9b77bf008f7df6b095e030fcea2c008baa7491665c9cd35e9e6edb8c6f727e1c7504fa74c8f39cf524474ddd6bf0fa018765b59735964058cbc78692888684dba4cf56bdeb2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5882ee7e4eb9113e7cfc9c2f2105fd548a6e1f74622a41ca042d7fc78754499d8d1e828c5881746221903abde5f9a0bbde48fb01e8c40b40dc0d882cb26e2f61d4ce349fe52a3b1e5d0cda1e1d6ce82b4249ecb94;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23d3a159948e3727f9d347fc2396254aff77a62aa18d140cd4a403199c9092bc09c00302ccad2ee0bc3427e5ace598ef1fcf8f915bdf7a7c59208386a28ad5d1c09622bf8067814e7ad88163e69ca0820102704cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fcfa3fc69a85569815f6ff64aa6121b9ff6ae2f4cdd727b6923b33c45fe41b8c9e218966049a1ead3da1d062248e70c28c85988f305a4cfd505cea228a77f833d489e45b0687027cc392ab39655f103fc0a54ccf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26757d45c8bfd7e26ffbcd99e9cc7876a3f3b1da36f87a7a4a2300888cd522283e690dae79af0efc29328c264800cf8116463bb8b7bfb5e9d50b8a9914d74a1ecb291ed109cf50e8126279bbd550ff8f781b945be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb251190c0534e38fd114eab52e30c1c9ac75f5b74cf15498c3cd309a44b2bc87ea4122b81a6de4ebbd336374791407b71d5f7195143817ce497fe11cd4717beab14f1f529184caddd9fea0c3590b1f09e3512778;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he93fd0af650165cfba0f2d3e007caae123a6dd1f969c7aedd3b3a1e70d6eb383e5530224d4e4d52e11adba6643bd113f1dc4f36422397b20fb114db36f72583cc6e410432f01d5d44e546e1795b829f28f2ca36c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h499344a20de61b5b9e00ac5c3c46fbc52e98eb22cdac2c3f7d2ce7371eb7c2b3e8e6bd9973797ac4035669d95992775bccbcd83e8f1810e303174688f7b0d2bca341e3e866947e2ab33a82f4aaf455ebc45696f59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ca3f8cb795bb415eba87284e8dda606c999c2fb91551ee4d3f30b94002b437a5f8f2eb4de2360f8aae30c0bb2e8e78bf52623d1e9f0e3ad9a2f17e7aa175a945970a2e5eee16dcad4b3d4131aeb3b9a5bd625e5e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h834af82f1b20b49d014bf73856d0d75a4e9d9133f4dda6fa296519151fbb900d7c886b651b04f21eed1f3b839df4d5df9b5901c55aebc338d01a97a6e968703a1fc35d4357aafa546756f8f6e00bc678965061abf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd13ec58b26b5595f6390b649aee34576dfaaee7e501237b1e141bfc11932127720d7842227d3a8866f932d0e07db85400516eb58a575afa6e5303dbd5175dd0e0688c140d06e4433720f3d0aae5eaba433b6eda3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haebe369de919fb10db3b396b4626fd62f5d6ab0b6ab98452fa9a03f283d00211541666d752092d9265f2dde69d7933f7a03a99995167d5bea0768977e0d96acf0d542ad02eaadd3ff324a8e7e7231a770ce523317;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cfce1aff81e6cf65029ec74d449ec58d1b2bbe6a0d087f6399028b7272a5f529419caed303650b9f2798f76fc7e4b3f03696379fbf01f30e09453fb4590048c25431c4be0a229796cb092992421218439e5cc234;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hada0a1d2468b8235c1efc1b12816c64129b00601bcf1774c38094248739c5689a3f2e8971362eea4903e51e5e9e55c19278a1307c400da8a49c67c1d42dca0f99af90de2662b4b84c14c9c7eba27789217620d89d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6834b0bd3b9bcc723821cb2c738d417ac2e2937f96796c2277fe541e0a8fc3c65087abee666d1c1613948a1e7dbbeb8c600bff3609e773d1da4385951bc0d34168cfb8e69b8f0e221b2430c4a2c3022f8c8b3340;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb24b52c2c4c1b0ee45d6afb6c800ccd24e6bc27f92f918dba8bbad3aa3c3330c21efd8eacd7fae91be6774f3680a0b800467c876b993a5495c9280730fd3fd81206f60d7363a9cc00209b17eb917fc8926c4c046d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h739afa88ce9d5110769be60b5320e3dbabb12e458515601252826f7b72f15bd28c25915081ec3524f4098fbf6d2a8f4b457d8d7a20102a07dfd87706aa8e0f1522704be297b04baa7dd29ae843ccba34e93639ea2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75cd822b8eb162ceed6d5316f2bdf05a66f37161ce2a83ae377ae3654ed5e3f7ae3e74e096180f64b184c7a84d31ba67a37c21a872d48c491f15d724242ef5ae86e7c63d3e46883a47cec0e7e84e10b64f1ad9ac6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h444c052b81e35e397642e15f5dd08f97a0823852c8a1f4ebfdd263abd41555ce6163388b03a2d5d8192e8aae8b2c3f1b425aab86ebb96ec1a78c20d13093acc44571b01f123094fb158f60c167a99e05ac87ac71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fec169bb86f2fa9c18a64c2f718627824abe6fd96754ace8b05c49859f91e7ea079ec500ca08fae82178412b2a4bc4ba9188421a7928df4708dcf0772fdf73aed0bdec4962407f0d7caf92b5bbec3e03059edf07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d3d7f9431293d719e3a1c1401c5113d3c81973497093c8299b6ac31fab653c52ea73d64787be9e24e2501093d41abc9e241d5b81161680fba94b98833ccff49d3c0ff4cf6f98382f885a8eceb7e332262c2e3d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2c3381a6542fd1270198843b0839ce25b49db91ac3bd556e21ff8dcdcb51e26db6463a68fa0c62d81894d0389e957b9bf6c954ee1d5ca7eabae80a52ab598815267d81a23692f8c19bd4d8676b898f3d13054648;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7141cdadc7b656095fca515bb44221f7cec21a61f96d1cf8e678a6b957b6a784d758c315af0166bbde4737d50742d3fa1e5237ed0c7d9b921a4d3545a529201ae711e90b1d7da16a9cfc0d96b02f1307e34bcd78;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dfce097cbfeede4d3fcc63337eda7bf87e4f624d11b2c6f8303f34c3130b8d9f3bc955c9e4ded64c62de9046099f5fb3bccb1894890c8b98f625acaa957c3c2225ca558560a8781998b1f392fffa06bfbc0de6b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bf906a13329fc14f6a424b6835523d470d6539cb4a1ac8b345ec5d5e8702d56984d676e137128c227bb26cc527d428f20c4fd01d50f780d56f0ad121e83f4c3aa40f4ebdec2b1a6201306216d3c693b274d328a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66ba741bff51fb3db3526d3ea31d7ba99393c336fb7092b4f5550181ede66ae2f6b6f5749900f6616a9080b5a42a06f9ff4ddd0249308c545ca38685312354b6ac86a53849edad65c599b0072d1b43ece162d31e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81178b51728fff9f3bde3c39790ccf294718fe8c98f6fc59ca2b84fe0ec0328e97fbf81c9ea58bdbf37b36d182390c1d87abb0a3384b54fe282493bdf52c076206e6f9a56e1e2384d7c20681536a315d4f2b8c02e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76995ff7b420762f62dfaa2f36e79772f29b0ddb82f156483e30feac29bdc16fdce690bfb2cabdd50b176c792155b4425225c547d2956fbbe74f32d72ae366e6e440ea78ce965184c82bc3bd61ae54d914ea73304;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he27a5462bfdeb13829045636942a03fba115c64a5dce040e75aef57b173343969c726f54ae498eab550a54c8451f943ac10addb8c7e10384755d7818724e5f31220e268e9f6f5f78271fb00af1acbce81e1e41602;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2dc1fe20a4e700560bf8f7b39071bae2ac02a58857e6d4c122b533b875da0f577d35e88e1431760387b28be496087e13a4a3a88a29ea88373ed0f11d4d79b23c5992362ebc100e0d777df9f73c002648d768794ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34b4cb5e154d827e008ba7eb54da40bb2d44e07de7302a7510e4d80468d2716cd4cb663b2d28a958baa36025277bebc709f595bdac93db50f0bad02bbac205dbfad297ba0ec8271d0caea0eec9d7a974f872e1b10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbd4acafdae9fa6e26c6051f16ccfb4ecac338ca2037ae86f583ce2a63b4779f951ebdce110612fd71e154a9b925a41b08ae92d3da38c40bd2b9c80a61265ce9767331c9cdcfd6d3dc72ac1cc462de2c0cbbc3085;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8816df1d6807763cf6f426456b4524a6884cc8f54b98c5db51c7c227bcf32bfeb44c009f648bc845ad9e7b7ab4934aa7bcf2f4c9fa845a8c5e91f42f3058c5913922aa1d631e0d47f37dab64c6b481e9747355f7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h683ff257dcd817a6b359ed449ec4d273ace39e724c0d48d3399afc70436c7166e82ae0744aa114cbc0e8488cad2eca0860918e1c3bae8a6f54483361c6b920302268b57acb4828b61c166b7effcc43bf2eedb1903;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc443eb393298c3ecf650fe7f929cded6ce7beeaaaa681c58e58ad2433f3371066e71e4b3f6412c0812b59dfe2d0d6f5509c55a952092eac3eee41dcd1cadf1258983fb4cf4081a533afc24a1a6e6e4f95f969ec8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb669c7d214b3be2be8f95a7d8c45ccd31196b01c12d3ffaff80328bb23023364422b9c0bb2b6c5278990b1802ec9496d2f48b994b8defdf79a5d90f4ba0ce1f52f05f4e9b46053a254ab0c678c8b2ca6220457c85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h141cc6b49f512f009e99871cf401016145bb62b1714dc78e6a782d6c6d8bfe769834be579bd163f294272a83d98e60e2737605a809ec1a4dc9b51b82ce5d0512c1b87521e23db0bfa7fcafe65a986519d0d57dbee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h472639f945a1fb15b3f00e5ba09463e37a3ab70492ab82ef09b24307f7bc24d4dcd337eb1806e0bbc01fb98ab8fae817636f0ff7a91751cfad1ebe9937f48a03322ef6213916ef4704989177088aac895f10ee6c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha030fd092c83aafa0e6590507454bf85ebf95949ad9571deb6ff2ba3a8fd3f379f92ac8d8f1d11439308a36e54dafa35d56fac56e44ad66b239928793ae70ee677788b0d0c208282920550a97f11d731f6967f23d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d7c9fbe39cd06eff7e039aaeb42ed2f062aea338749fe39e007334b8f020f736a219866af74c88514d48e6ec28495e4a768854246031ef957afed9bebbfb23b6f04c8c6cacf1c222261575b491b9f5a34ffa9e5a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccddd80648bfb56db0e6a26a0dd5a47095dad42d02da741a0db8707f84823baaa8a9dd75789f5a8f95da35521f0aa4089f91ffa3720aa0e791376ce405ad629f56fc1e0d3647acff67349e86809480908cc573606;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48a938f85a89551306d27850c4762fd2db337aab40f8a4989188ea5d458872788668f5bde5589b4dfa8ad3089e3eeb0ef0570b647b36978ba4928470b46a52ba0e336fec3e029f793f34a6e02c91ad51358a6db54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6dd9336808a00989221828eb8b6137368973d19d7097df921eea64919371b7e05d545a5a356f43ad57bceb6f9fe8e176c4137ed99b0965c64552ffa62207669dff0394efbf7e6a86b0af1bf079d8bc4585c3aab5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha375f6b3626ab0650f5f963a74b3db07facae998afe6c306afa070b26dc17e6a6d4d405fe32cf33b2846cf7118a602167299d12a60c819c7b668f7a90b7b8812624e45b150109067a2767917ae5d00b9f09a2f0a7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1fa03b869ebf82f857929d70c6dc1d0bdbcc10bc9d6fea7e0a4ace5fe9cb76c1df0f6d5306577c93b06264b98425c00f271fd01a16f355e3106c68f6e28f944ff86df5e4c94048d943939e1554c266b1af9c3d6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39b7485a1907ef00b7ba1da849dce2f0b3385ddedd5c60faab9251c0ce2417e97b385404f4ea20132e182c51ad6ebb54fece27b6ddb07638e2b68eb3151091b914a08a4d4ac2db8abbc6b8f601d72c8d9272f247b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdabc6a456987d4757b69554f170b1982a3c49efa4b7157a3572d5307cc402661df0accd8e35f449d8c5cd20aa02213f6bea53a6d19ca831e91c3c928e192b08345d582c0f24c4633a2d3a5c4ac62cce3d4e2c5469;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2778b0e68571a573fe9630f333ae5e4d322517d86b66cbe2b7f2d81f51438401d8861e436a5ac0bd7f9402be71f3c8e9cbc4d9398e26956cdccc79f02957ce81892421d7cf4dc2a835a2bf0229a772afcfe86c878;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf69027a9c1919a9a7779eb744fea326d910d58ff8faa4e8af0acd4d96332be2d24e109f42b257e5578fe14e1c235185eda8e67c5031b8e8e1780c4151301e28b7160c4689763ecc16c12324e9739b0148cf41f687;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h772b7ecfd7929942a57d3ecbe48cfb28ac3db7f8365cd4ccbb60fbc39e659452116f755ecf2fdbc500af4aaf02f5ab9943ab31506ef352b3eed68b16826d7e602d5adba2a0277d1a72831d59752a0ab1d5c830ac1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa5dc5e0aa39b711a9abfa97ea48ce49928e868eb3aee0c3f4d979eaaa6a9937cd351e1bdde291ee6eafcd2fd047547149b2308f7b1ac12516b8f2c159df2c78292ed149eed1d93cdac3a00bfc71d2d3b355fa751;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb620333a75d9a952109a7aa5f0e47142ec8e298c103c52acc6b0d4a8618657ca81a22f698f49a78aa494a1786b451a5b529e13ce6c780834b1f7b5e9b064373239e68fee44346df703db03635413e45bea6acc071;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cc606b84d15569b8911b56372c765229e65987fa2ab6cd41d3941d079c48f918f4a073077ff5af8a124de5445ad1df25fb63f455c50431d9b00e3bde379557270ca035f50472ac364bfbeea15aaf7f4cf38cf9f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74c35d6c17feec7ecec0d9ad1fce18d84cf4353a83cf9ff068a2b3b97967b454c1c626854b92926a5e67f424b616e67f15e90c6bf84f694c8d12a8865ddd549bf633cbe26a20cbfdc9cf25b88e3d1943546245dde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc5d7532e79bb076e2777059e3f0dd2a5042ef0d716a4c4cec3682981cc4f2316a6683145e8f3ff0eae98a3bd71b2bb85eb3b1ab5456ec758ea16990b7ef7805d1c9c008f6bc8e49515acf7e5718329553eb0371;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h324f3fdf8b8d0c6ed89705cf3f632f111846efc46b57cd93726b8f26a9aa03c2fc9daf881600869f37e8348c19eab070b2a62ab2fc28a8b39f5fcaed825188a38a6b6d3abc91af0c5c657067c367fb3ef99e216cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11d928702cc2a30eacc8b82c60332ecace66268025988f3f00923f01b7744f7edfd3e9f58f5b8f2372fca89bc4cd91a702a4ae40a0d74f8f5378b8bb9b95f588a6f03c0046f7e3a6b3bf5e1f8a1d36ff933e2fcab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he76119fb75e6da3ea97554761bc43633b6db5a9928a92e25370138519551bdfe49cae8d9b1fa548d68bc9ee4586b30109452714c4ae03896fc01991636b2d57d2725d05a515b5777365afb43d0979ab36443b24db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he764277d2840cbd5d4be0a60aacd066a7a5252e4a64ef0849589f4f640d84ba3e31b251d6f3876e43c780efafcb330415a9a2e537a4ab98d2bf46036bcf9956f1f5f200072b53da4268f83c3356280d2ac43c6fb5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23eb35ba23f64046683e1cdf2ad36908c339fcb7301ac5f33f6de1cee6c9f802b5accb37d669c21e24298230f93a0dce13b51e94df8e93cf7e80069894b27db640bd683c3269f7814d2a292284350583061e9070b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbea4918eabbc5064569413714d74b9c10ccfe183ab2c77411d4dfe606a518b98216cf36bb3d7d2994fe96db45166756a2a905450c018dbf1d7bee863f38bdb59a964506fb48cf08cdb8f4b490429421cd2de9a0fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bdbb9f70e4fb7a810df08d8eb508563361c889d068e5d76940363679ecf987af41c47c7921df4a4ef388c365c48f08bb583104b51e0d3d36be433f5377f54ccea52429ea8134af3b4af2dc8ff972c2129223ae45;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62461450ba53e9cef947e2ed1bfb1c77f1a9a7780659df7f68ee2c021c1b82eb80877eb79c05de01a636fa8b5f32883d2eace7efc2e0349683920168251ff32456ced81c0352612aca4f40bb77fd9e04ca5f7878e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2434d618f5cdb9f34aec27f88c0cf394e138e0179b242b6d6d4122ddec33adc19fa647a4c6fcb109648b14a42d0c32e126ef4f021dd715f7a16b4421f90bca4f2a0c441ce56f3d1fd65c5372fb6a9d8d7ad544b7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa47a617f4a0727e6939f935c77692619d9dc1ea139d31e9347d6bd34de626b8140505b6d913c73d6ca24340e56e9a118f25bb37cad1ae44b241bf5d7497e08b16e2773c1bc8bf4f0735015e395ece292a1e106fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h523f12fc369c53d0179b4a4cc81deaa6628638254f9a298d04fc060a2c9d99119fc89341b4fbd666420cae0a6deb593f387d9884aa8f76e66cda579230f62c296956fcc97d0f0f71a49a06f7c4245469d437bff05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9572c9bc3cebc4f9b385582891f7b6528802372a726c49db2cc3392a56bcbd9115aaf58930c57eb8f224ca487527804a96a1dd74cf4daa0293621a772ed0ac78daac6a52de322f8db40a63884304fd18f52c9a918;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb974dbf07bf9f340cbaa92dbbfdc4da4d1b8e40ee44ca10ff49805b5286849f02ced189965c7276ba9cb784d73ec34393b64c368a5fe60a5fffa0a9dcb9f245ce204a20d9d28a5b97fd45eba483a170da6d54b18f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2be3a7b50e8076ac0bf5de0ec9b9322f4afa314ec36591c386fdf7ee1cfa566d3e4b93b3ac090619ac7e45aeae2d774517113dad4c8bbe287d2ae24234006d39a3ea31bc94622332a5cfa2fac0a1352c86c68662;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h718aa6955758aa4906ea52aad239c628f396cc1db98163060c36a86356e412caa20b9ce0b38050e1d0d6f84ccb0af669a317d2f5c6c25f45e5205c7a67aa0aa9a90acb4e62534b224ac3003997d2b7ea0dfb14a1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7697d60fac3bb436c1f8d16d05d9cf94a89401e1e84ba40c049e39a67ea85a5b1b683f0d1e258789076adbf0c34bc66c6cdd4a6413bf920f5e17f992afbcaa44a568ab97d7d812b9ac6a9c4e215b4e9e06cc5dde6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95c39244157f165045fa54f5913ea35f884e6d570cb2b876910c609386ef5e702c5230f0b60c6f30077b158bca6d6dd35c4b786bd58e670664bc0afea301c49d63bb5fb2257f856906c73de77b6c58309bb33729;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1da9cd78413cb97939a671c4c0b59e1ae64508a0bbd54b301d20947c253c87779fa09702a837b6e012975bf54940e62cb8e423023f2e5b712e38856eb5f27fda30ead80aa5a02219c2f447b44a02a553c7fefc682;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ac32989806e474ada3490974c233f52bafe426049b6fa5acaee0ed66d610616b081660f2a37f551f0be2199c8762967c9ef9d59f33efeb1cbc2599126bcbee0c6ebac21ba5be8127a10d937b0c276cb4bd724d46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h395c988c7210351197a396a9bf1d699a39e6c1a0440e4c3ad1e336c0dce425686407a5abb791691324f17534e28450d0aa62959d80e95aa5074b1ed77c7aab77ac5833148f670684db9e829ab2605b61105abe40a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9596fae0e74a753c0ea1b3389f1bf97b2cdcd1f6cdaf97f7d4f69eb653b0c11393eb42842bb51e903935a38f2e79df022b9667535018dd2a60c16050c4ee77bd6f2864a4dbc541e25cb2bea889160974ae89b462;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he44a8d0f7b08dfc67bc52d57dd08e8f3eb3c311e8f59665204603d1b3a10b041df27cd6117cdfcc2b385716fdb924f7fe2d59faec732582a2836abdaf409e581cbfa9db484fffd92cc27369cd3ac5d3b7cf10b666;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf94c7b730ed295e2520b9f775aba16056740885d23ed746533b812b6665636a12ba5ac60188b90c37dd810bb58cd1ba086592169c98ee81f7dc21e317c4db8397cac55ff2ebcb42c3216a350dff42be21afed5f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8d1df62ee691956f4d1581282fe9de0d69add8327ca0c91c570e23fb3729f9d3cf7c8c9babb0c0d2b9dbcb0a0ae1f082b4cc02b2ddc20354fd3142e0fa22de3cc2e7c42fdea9d30fbf278d197fd221a348f58f26;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76d5c40df2ab9936de9a5ffe660051f0d681437209ff9ab9230901a5fa73e30eefd7e34f28ba3cf24bca2515a0f25e4b4733e95c14476bd5cc8232c1f63b8c12aee446c71f405f481aa3ee54023f428e63f96cf12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c338bb24baafc0e949d50039ff912603e6467ce4f199a47b93c9c5d313218db2be103ac4f6a49571503d252e176d02f1405e915720e0fda394c66007b85ec951261f37c0776a66d43117437dbbe98313e3c245d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53b34f8aaa636928de326aa5faff1849a15583802c5dbed7135ebbb9670077139bff54449e19c74f13486827485aae70f34dc3087bcec143f92a512d11b10a308aca6764824ab33c9c3a229489852c3767169b89c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8875ca411fd7ff6f457ea441d92d50f2bbaa4b6a30bde4008eec68dd06ce30d18a8d7b38a68ff607b65a22edd7dd0d41da7065c6c6f2280b553f03d48d1945a1504ea3b569c56b9ad3862543dd74a3f16702982dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ebb654a8d97ebd2f43a8edf7abfba942be951fe5fd5100fbf25f4935f26e0027c731b6431073c242831d7b802f049309f71564b14829825f101b3cb6928b7732f55b0b4159f0da1249de2591f22ba105b18c1ee7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c6e742e41da592f9a2d94c1a3559398382b0b2d849cbb6f97bb687dd857acbd285d64f4a909233d38dda422983730a8ddfa5e87440ce111526f8c8acacd9430dc5c9da7b77e4e022b4ed8e01089c460d41bb84a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94c07bc33f5f2c057b040ef92070b2be9aba28b6555cd538386c42ae17674b4528a066ba1faf195cfeac480689d8004d3725e98ca505af922ea2cd69826993e29b683c0704daf6a27cee956382089f45746a42c73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73ab325e10e8c3a6fcf6b394079c11a0baa2aac03fcea4e6f9e908dfd5b65925c226b19a523ffc8a356101697982f2bb5cf7a76c8ad9bfad7324c8cbc337a15d6415ad63207e50975086170e78db00a448627ce4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97a80f1676eceeb25a0c204daf51866c6d75656d2998d0bcb57fc9bda4116a2f348ffa58df4ca14ee6877ca932a72d1ad2dcd42eec01d5b83c1bae54e6bc0fca06443a37d63d459a71cd646d52535d1ed980a5c66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heee47080078a03247944a3aa1af96f7ce824fa11c653305deffedae37afba5dd3a0707671b798253504f0d36ecdbfad4b2861dedf1ccaf34d2bb38c12ac9340179f9d27b20148674f5d7e0f20735362d61456f8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48710692548381949e11db6c943bdffc9fc234c9c085ea5699613dc7510fa80701670dff9c1f79cf78b7dcfd36a0eea026e14b30ea38995d61bb68e8e0944700a29c00b4d8d79ff177cc5915e1df20d9b856e6ae1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffaa1a505c15a7338afb005508b35c6f44b307c6699cebb47f9601ddd896d3eae2c96184cc45cdd329141bd4f2f890524e90fb9601ba5020634accdfe29d13ba04ed5d61607e7610ee1304d84ec4facbed6f5eb7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5da6dae6bba1f265c493966bf2997ebe6b13432286847d335d61928c63fdd200314756e71aba26876597484bdfddee0d2e17603805d4a6063987a58811c7204e88c445f8df43f5cdbd8657a736af9907095b26bde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19405bf798ff84665e573898616beebc4f2a82dcbf30a69cf82e3b2f6c6ddf72046b1e1dc9ed63eb62645e1b04dd6322235b2dece2d56d64bfbe4d1b89cdc64c5620b4ecaf24bda85c1df5184bb2574428261976c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1ab96755555764018d925fd1c407efe31c32f53524c2e20126c52bb09264229029608b0aa939ebfe194a21dd496840c1019a0a77eb63c52a91dd8446af58ee3684c30a36a258972619b1e532339cca9842e6e704;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac6c977dd214cc83ed6990ab3c58efedaa389e42d1bd1cd21d84a978ab2dd9c8215087acabcacfae296648f267423bf23ec75523688e4119207586963f0ec471f5ab140587f65f6333a47c9487fb4ccab5eb1658f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he81f2048d83e04536189ae96e58bbfe39c945cd20513a781311b5b5078ec18af957719e3bb0f28f6b57728f1a6ef567f6fe504af8fe290e3c481fc601d98812162449c19ec3ad53a4b780c14ce10e8a26a9c8f9c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde46bfc36e86839ea907b48c5971322ae09f0d74c7777fec53aa63286eb89ad9199d098cbe02151789434d4fa37a715ceb266045b69c2034e6883eab4d85ce95a278a12d5191d57897ca19cd927591796042aae34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc99b4ad8e33b9a63e769a64c9dfd4fa4d8cb71c2654a203633ee539e3aecd7ea0dd9d83ff31dff4dc61258259165d5ab1c6d3e58bda53f67352d76e6d77ac693ca2c902837ff480df565c22ffa7cb4db9ddb2eb2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8aa11fd63d46bfae3d087b3c9f4b313c049517823d12a4278ad67af2c8eb633df2ab1ad426c07a4feb5e3957d1459f4a4b1fa0a6b76f910fa6bfb6ff70dc3a47dbec278c3e50fc4f6ee8ad5b3e806749a4df9af3d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7790d591b2e955070a126c23c28b7612ccd22643de969d7ccdc99cb311297855eedd5baa39514b6bb4cd35aa3902a37883e90ecafce96976fce5ac3f3b64e7f0bda32ebcde209e04d1c8dfcc7789d75d205470396;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7f87e546ff39dad49b957983266519742d927dbb683046e7e84e82fb4a25a2d1b38e278f331ace9f4f12b293791705f6ceb538688faafceb980b9be7f6b77ed3d5cd6d728712f59ea68c916a54c599652ed94a2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf147c342560b3a8320a008172f54cd2839893f02ed82f20e763d5b7044ac78b4456592326a8e03c4135c9ceb5a4c2a6bdefaac239e2a591297e2eb99b223aace58be1d6155a46373ba8fd236098329f41815f8297;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2b04fe40d43e36ce9592696803d753229e5dac20250a3cf3547e013a40b24864bee7e90f7ecc04bd5bdd28b5e39f577ff1539c4f38bb231201c8dff85da136a29e1549930da71b3632afb53ccf65a5ed6f87b513;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2833b88d5c3b65950c9fa8085d8efb659bbe8286a97059c6c7b78b929e4c208fcab9e911b41897a05ba98e394553bbcbaba5bac76e7d92092ccd545ddfb3846479f13d0dfda9eb474847aa1664ed57cfde55ed1c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5a8130cc8bc206766ec3e66d67fbd342b5b68490049ca1896b34d2021987b7ab7ad4dfde2c71aa6c184d1e6128f8e1acbbd355d5e11254633e34f8e2df0c57f1c9f5341147c65101ec1e8ae63d4198018f6c06fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1db1ff020a3e77453e318acc982e14f4fbbbde0055413d506e21dfcb92736b4f00d2c9e993e42c205d7440d31f6fe4b87a13b4a372b10763be7e91609f09ac875e475904e3e1b8d17f45b00af9ab0384adb872d33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha096b8db11eafe0715fb104332ab0da8bb16b117b9fa16483898baabb4ac195dad0330b8834579b132237cc7401e40605d17599a765ee5338635385c68ac13437d976c0f66ec9cb998b9e42f3e6d071145129fa46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36dc3ae7d82c13afb5fa8e48609e950c3bfaa746ca4eb8c3d4cb881fe34b8cbb6743dcaf7cc8033e82f1c794f0a1cae2dcc83d3192d4661b256b5f7941a42004e5b9be314d9bbd787a4a2458f24dc96b10009eb16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6177b7875a82f7df6ed40b32774c1673c645a53291b747623ad2617ade938a402deb27215aeda0bd9ba8d9ccb1cb20b3b5ddbfd112076d3f45bda152b2f03a3db1e6896e0710e2fc97dab8375358a89896d5187d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca5afa39ec62c0b0cd589427b45508b372ad292fad9b3ea41a401254bc7afe8f2905b3ecbefcdfdf0118151399340eb87f8e04c172048af37bfd888fbe1cc45064e0be8a1d22e8290ed92b648d22b90497bfd5554;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ac8f0a4666903336abf250663bab4942c1374b91a0ef7c5a35cce88f875ba14b649f5165ad0808bd36c99cd490df2013e41d3da81665f4acd26f2734ee22f410fc8cd362010ce6899c2bf3707b2a09476b355daa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6744b4eed2ea3ea4b0534c7790b167ca98eb202a6744552597ebb11d5bcbc8ebbdea4f52d4b812da67177b9eff2e1abc1425266b3ada736db57139f70e71cc3c32ae3b00572017a57defcaa879cd2097f0c4d741;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86856bff3e31c4ec4ced0ef0ae879d1edb17fc4ba37f6d7b0ea13fa1772198af0fe5db0d17720d518d757ee26ad5440ee25d7c2b0edb32f046828040f567bb3b1a2d1d14102bdbbedc292dc63af2ffc2b2f2fcbea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3cf32092f9dc07314b1561c27bf3e7c6742c7e581b752998fb1db99ac949d785de32fba682b2da101738e8ca8d2604a292465460c9884e31037d873ebd4314abf9ee47d864070134bf53d6891f4341e213cbc9e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb2485dedcdb0e9286d8d14bc38c75bad42a7fc94d5061595093ce03580ec714fdca1af57f607e56affcbbe3c61523834c1e0e6cd5c8f2f9fcbd7e669d1afc52add890a5b811250c9fcda11352165ab09fd7a6d57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h627efe43c05225b09f80e3a7d72108fe6f65afab429ab713d57ba9ec3e1ebe7e8da476291c875709658a9d14f6b6c1d94a9e6226ee5f12b65cd25f7f542cebbe02f8012b1ac0cfa37244e53ac54fcb214c467c9e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f225e9903aa804b1aebb1c4e205ec5109c09eeb7b27b5bea6a31d05a7dc65280fa98f99dcbc30b76e4645fd9a043884e62cfd37d484b998ca42995bd108cb4b8ecd8505459a0b94080554db5ed947baf15722625;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha793c67cc47c6ef11eb2249016f4a0a10f71bc72291e31bae35433b55248eeb4825dc33fd40e870e0726436af86b7f785d8c2a011a4bf032865817e0808fd59ec08604a6d41a8ed91bef5c0dc612fa0de84ac01c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2be4ed2e92f6e3bb475d5614116cd1bcc66be2622c54a870f6ec8ba94c7c8e854d0477855417dd084493d9a8c60c89a811117f49232d6dca4ea7bd7b7aafb6cadfdcc2ad204b219717c6536c996bac0365336d8ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e576de38a8461e3f7bef1b26ef692eebd3ca0a4f029db0a6d9e9de7ab44e665ef4abd635a74a1dae24a7cf51aef6eaa20a99c6ed28b97d5c736e2395c909f34a572eee712b370fcd4b8f96fb2dd2e84956dc23f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5ef01aba499858fb07e1cad671982c9ed63946db6b20f2fdfe68fca50865d0b3a31af886a1ff3481a03a31320f055b727aff7c7780c23f78186d17d39959fcbf99c88e33369e35fc5a94835bd44f4c21aff39a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c0b388a9501fbdbb9f6389f973083548bb348a8b0061e50a60e93ab0ee89a3611e8ab94ec77075914404a88fcfb823f9dd398b07124a914833e5c595aec67941959f150fe092dd7b6c28a3f1bf37381bbb249830;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7c03a82b9d18e45833e3a9d1a7570216b7f5ff052b57192152a011196075a70226a4f502a8a73cbdae44171f9ee5a2fd8de5438d2822c3fa10d9d0d3cd0b53104ee532c30876246bfe7ad630f5cc1fe42fa3b54c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf240fbaf476343b5150d0f122fdc0340600c638466ff853d93c023ca06838784924c9a9a660072a3eae7e021718364078ae50de0a13bf49f4735b6f7e3314a2a9c3932d003dc11fa409bb51881ce29e82528f8ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0afb5e6b0eaf4cf489f7b4970c99cedb4ca80f1965a8a3c689d01dad474fb8f8296b2162e5c0f623a1e3dd59826f7420a75b42e72e3d8e2a03c950d6dba432dfc76550931942ef9a5a1814664cda4f09d0ef520e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab8f92b5222b0918333ab11534b8ccccba4e67dc95a19d00f7fb72c34b833e0bea1262668275326583cf5c3c738eea383e5ec575a3612d9e836b933ffd5b9a16acb9a4c3757ecf1069989422adb964ec9409ad877;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56220dd2f9613033b9c2219960d5e3cb923be9d4db9d60fafd64f8967a51dfb70df010b1f5dd35b3f741bf1adfeeddd8c71f9fb45948ef67b4040fca5d5dd4883f451cd7a99d51c086befb79c6c405475bc988174;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17a9923cfec300f528881de47d7f9fa735a774d9f13d893027eaca81fde31246331c8486303656d1b317b13e367e8eab8349d54a0807062db4afeac2b8faacf440412e3d72c9198b4af04d208e0719637e8601a1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4c4d90486af328dc1776e2d088f6c3f06fe7e72b9ed216367401d4beb812e11a367834b1814597e9068eabee6ab7d01ffe285f359d049d36bab98997bd215872f66191804ce8bb3450362aa67ed59f8f722b389c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7eaa54d93c6d631b2a2830e827b562c5a75bb133f7a4ba4aff5bcb1f20d3ab47c81784fb6a1be077ef2b9259c5967a68385c3da0498a19b480b6f4cbfd2e6b8673330a4b99227df9d75e77682e4eac3f3923e35f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h329cc01f4d804dcdebf8b3afb55c8477920aa33c9dbb4bb16c2d1fc004fd6ac1be6da114f0e227eb015e5dee851466d524fe4756718bd6ced98ff167cad2d710bf8d3dfe7cd22cb180d0c98853ce723630b7b29a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h127fb465d2769475cf2d86563875d03c4fdbf1dfdc578b0174440145c38241d08c4fe9dabca260593357701b5ababf7b9f5f85cbadf7c6e3350352e510b904f2a6dc32a43cf6d7b232440447c0c46e2ed42c63066;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b04f12f2c84845c41a2e7625433b62c07d1f76507be45b07cd1a7f37ddea98231b9247b311cae8a2b5c1d0b5b10d8cdd369529494cec48a40eb60d68bc768b9efb0570cb99aea62549442c607ea79fc2492c7385;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h296c2ba3a1dc6541d5cabbd78460142b24a963754fdd453b454d0ec0f6a06352f60782bf709145e7967bac789cb722ad3dc4d9609ea499f60015e257727e5149aaa7bf17538af84818efa2f8ab774f7a9ee10b865;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc2210a180803038398dae50bf4cc9fb960fb0f1d494cca6fc91b1452e0e32fb00acf9deea82d4e996d864afcb00f1f31bf37e547ef8b2e7a941d2dec9e7bfdb937e046724394c6c6c602203064344e3abfd15b3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92ad80c04d7e38c83226905cce2287512b7443ad7bd1f6a86148c0c1be48934efbf2901942393463c2f8d4531999f74ce161b00d538c3ff45f76668b4c32562e921aef5f4ba71f0d6fa2acaf969679f7be8c38c90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76cbd01c69d20edaa209f2c5bec2e0aa430b529fc5b5e99773d8d68e266f49e57075f5961e58c8864b656b74bf88de6bbd0b7fef3095865bd67deb9eb4087b5cee8d5dbb72a482b520637ffc1513b403e9805ba7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he29f64a8467e71daab83e465da32841d1ad43850ce5458a80f316f8c86d7935343283e9983e279675fd5623027cd409ced5e869b07bc1726fbeb476914952cac9e4970e67cbdec7169961dcbc81be19ed1ec71555;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7e6d2f4e210ff7beaf466ff017fad52bf4fcffb6b5d7186a7e715eb60bca34b40a92c46b7e4eb915954bfc43eaa5030d993ed156681122302861c4d0c6419284cfcd84d3a6f93d2e02b04d1b72235212983bb629;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc43857a15ed5e97bc7624890a6d1f1a4a3f583c04f7281ffc806cb2e4277d90c7fe161ef6e0af0627e553dffd2148356d0d0220b1ded2f10467ba3990e11ead734799d98b8e27de2f9c0b27535aa690eab482054;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbd56e941ed203a46e61654d2522655ef14e1b8045278dbd43e7b8dddaf24d5cca9d8b354794a1dacbd054b7c21fe5e2863a87d975520f380686f60241f6d4aa05a60369414f9a14975366f62df5107fd09cdf68f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdc115b53cd263685faeaa2d1c78beb4f460ce0382e5da02317a6ce5e0826e17798c09059af1a17809513ee11979a29bca7f6f6792bca8daefe2ae6c6f5323501a2c8b49e358517e22e4bf457ba932fdad3039205;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d72287e7114bf7a037d3fae5de46597295418b168f597147ccf8ca91ff8445b44a8723b898e2972114018e91c43ab7e097ae16dd0866392cf1612edf9fffa2704b0af56771939d89dff5865a53c2d53c441e7ce9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49b281fe64b574c190a1816543e8f7fc3043e2bfbe023e6fcf79d97d73e6b3f4af01510fc1adec1cf3398bebb2126df2c1a7f3d0f7aee37cb4ecb6dbda099f44034ef9ba83977994aa8887dc6c64af27456fcde85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he18d96c3c706b528beecad957b54a0ca06c41745352dfb684380b493a8a7c2c65123703a7b36c1aab24acbbd03a75405fe834acfa299b8aa152767d10b971c510ede9476eb85d830bccc49744a15139391b5dcb2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc070838b17c8a60a70666ebad9bd32ff394b3df3ab0b6d05d2824356fb790caea91695a61bc387136c0eda8191264174027595d7081d39325e37e022e6eb2ec55575b2d0fd53531d0e68daa66077e5b638c7d2ca4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef76df8a37b59d02579561f06eba74a70d253843820a9e9fc622da55ef1ce5a5a325ac7ebbfefe9bbaf418221b86d5fcf7b96d2d22b4952ca2f68ed0222f8bf5ad15511c567b7ea2eeafd9e6ade082ab6be40b956;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc3e245e06b96c2f1a3d59c18d1c37d27782f33b1180551dcb3e7842d55f1fa1ce7b287d8bc444bcefee52156c1fbc3cd0704685bf751e7b052f6aa4188e856ec74cd5728ad8054c43c5ed607add479841fd4fd9e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f576bc1fda7284a133cd73b0a7e7e82aa594487f284f1762a77ec393e31488f4ddf9f202a9d3d687f048386b7c2102221341054203c6d9b14949ea59223781336095b561c53931ac382b63d3be49e42f12f6a67a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5acf23ee7d553031f48e6b95efce85bcda9d606a9941284bffac3d1e31b4d1cf41c568890308fe2c333b347c86a60034c35a721abef6309335ce3e115506a081e8795f4312fce8cb23be0ba427c0da0b266628af9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb57c295da70c8c2775e85a34383fd36d8dc75d113f737dae5b1e838b32d191ea0ec8a50564ed4babf816523dcb07887c464fa065cd16471b8121e02dc694dac2df677c7ec38b68173bc76cdb004c20e3ebc2ce3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed9b2a63cf81fa04603210ea034e8de59932ebedbd3816a6d75c4b496c2319b3d35c231ec0343707a9b39f375454af203b094628ef2c2cb10ea1300f8840e692089a6746422f7eb4c4f1a983c01aee09521897cd3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h162787e47d24e79835e7ff2c50e35cfff63a08d5d5b5ea7bad02f008fd891ddb19d47def71c7a337aaeabf1836f4c9ebd263e363c18b78c36f1f7d0d25208b52b1c10ab802d8d5dafde03dea21aac56aa68c46407;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29eb31426af05763dfeb70583b2bcab0439d89599976cd5aa10e7a8560d54ea1c2d7fa0cf8b0e13891542d9b397d959ba5250b447dfcb7e958ad98cfd016d83063330768f45a5622e07f377969a035a462cb68b23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c59928ebe060124c9dce7079d095bd1f6aeb7596e1d40b740bd00990f2364d210a096d5dfe88cd07cbd09af384f966c0eef8098b28b4587d7564569aacef72ae2ad719cddda92a7c85f79d1a85e2f7203577ee68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h222658c9d41912eaadb640a462188c28d05a4b871ed7283495abf158a6addea4798b31dc1bf3c60873dadf8218541667b79c71f2455add8dbbee37172e6ccce76ac424a058d28bf8b0bfebe4b4a816624e152c59f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cd3c7218a65c83fdd64bf8c928e97eafab305536090a151fc1a5b1e47232f735a6ae97b39efd4211a9c19e3d661d7e7ddd5d3bc2227f5167fb7bd46e07dd2bed8c18df7d52de733fe9d0df284270eef55960613;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf98bc8d3198d0173c78ca93c63e4464a92883ae86dc6df27ce412fb55eb061adca85a30078cf06ed33d865cbd1c923a79d1068203acef35300bd911ef1ed9c2bf31176941f6d4339a08aad997e2f041165dd7740;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85189a69b13bde805812682459f46ccb3b918d067fd8300f649689f27233b1d0f512c55150a50b99ae98758f46592d472eb0b8c02e6c499fb8e226c5c5ab999fcaa7a27fba0e5192c7147d6e90d69b0e96157d9bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55d85b92746910cdcce7eb3f9984cd395c998804a265cf1272d241d4a47c1581e0b751a8b8c8e7682c8e981649f4f25e67a1d4b12810cf7ec6f0547afac63f1e7432afbdf8ce1ecf61b66d13ffdd666b43a55a605;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h839705e24909b5049adb369d42a58a120d90f7e4142f23736f0968829012fa64216a272043227845f68bddb8398ba2891c0c56f874d1a1f07bbf3ad00031d4129abef77584ded4e21bb620f81f81ae56743e2dcb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b5e3c614b1fc3e9ac79a864f88ed644a62a131261f8adf3993b6d756ca62f57d78cd0ad8bbd8c08cb918d2e43a50be07a58f4f24449d235186f57fe84d00add3032725a9de4767aab7de0f10d7f6e1729e3bfe4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6a1f154af61b13009487ce4cfaab226f83f45c3127f9ca80d9273510c4c79c7687a042c32358b7a1725fbef26111445e4731eb38ec43d9232c65e9b8359c5a99ead076bd80740b74894fa04531e1039ae33eec29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52bfba893177b41db9baa42905654f16067c80b2739824b972701e063c429593e829b117d7f62631c8672865c9273013d1aaa15fa670be646211b858564836f4e9d1a6b7926637ae76f33e54fc62807ba965833ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h237a65f530268d57be65e4a5f7a4725773054c3ca57390b8056be6a0c69bd016d5f0eefce84b43cf098ea40d5158ac0e7cd4afc40ef24e9ba87b9f7620d7005d9a4e397ffa00ed0ad4b0c108874718e66aa2bf684;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a434464c7934ff8bce723fa5e28d5541a9da5684e5b91986fcc152550a443f0adc43cbde9d94dfd5a342b0e35e2187afacd42a2ec16772b96a57c3b0f8af85fcf78fbf2c2cf647493e18b6cdeee85e466c5c095;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b9e1238f0a6c735a1941acefc7855375e723d2170fc496f1e8a62460c23342d8b48743db8e0118fdc21b0cd6c557a68ea4e9c203e86d1eaca2c9234ba34cae92e9830bd4908e9c75e3aaf98177ca51dd556a0df0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcb4574dc9e01c815a86357704da8ff034e68dbe0e75af94d04ee9a60b3a456e870fcda8abf147c7e05d637045f39a3e5b4d10f008f12ba1071cc710f1646c519eca013feef62ca3f7a7f6eca4153c4aa69c4da6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27aeb5dd9e2ed5ba402d9c4d56978114e3c5ad926787675ee46c39923a9482878228fd319318b63f9d902948d02677141439e62ec27931cd02ee11039538cd279d84f15c974ee5d43ed6c2665472c9c0e68bc4ad5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b62f399ada816270cd6ecadaa53a8a9b842110d11bbd0160d64c8246c1682a5432a767bd69ed36d1e2227c2286e4a37995f18bfc1616cf1cfc08f9fac14f7439eff484b0cc8a49ec25c4e9ea1cd744ef84adf100;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6c6069078fab4a5ff959cedc69d49a166daede454b3e1eb2b5a61fdd86720deddebc0f0cef4851303fa30edb23ef3852ddc89a7b69d4e6dc0c4c8ebacd4fb74320be420a810b301c7a39bc64f9467ca713a9dda6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52a3bc20dbbb5da60717b9d0c8da5eea14945b26a268dc740ea5fc01559f4b6e9d90cfb458fc4252692356c2a2de2ed851e3c04d9a926a18653e1b9346e29dd7931adf50e245a220c49ccb9c58f2d5852bb5600d4;
        #1
        $finish();
    end
endmodule
