module testbench();
    reg [25:0] src0;
    reg [25:0] src1;
    reg [25:0] src2;
    reg [25:0] src3;
    reg [25:0] src4;
    reg [25:0] src5;
    reg [25:0] src6;
    reg [25:0] src7;
    reg [25:0] src8;
    reg [25:0] src9;
    reg [25:0] src10;
    reg [25:0] src11;
    reg [25:0] src12;
    reg [25:0] src13;
    reg [25:0] src14;
    reg [25:0] src15;
    reg [25:0] src16;
    reg [25:0] src17;
    reg [25:0] src18;
    reg [25:0] src19;
    reg [25:0] src20;
    reg [25:0] src21;
    reg [25:0] src22;
    reg [25:0] src23;
    reg [25:0] src24;
    reg [25:0] src25;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [30:0] srcsum;
    wire [30:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92f06a335244412c4b1420b2af96db601fafe5f26ff63eac8b1f89d258e7f7a8c5de9d75b7fba84e17de95ae6b410f07aa3a5249625c67c2666d7d57bbe00e02b0c9e3937e5ff63443db83e65efbe5ebe6fae2093;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45588fa8ca0dbd0fd9a4ccb99d0aa8092101848acdbbb314eb355d53ffd96e55a9904c3c010dace528db88e0f38b5fdbf95e8aa4548dddc77071435c6c021f8c302f0bf881573ffe5aad46510608da4acc8fa5d75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4a5c18837b7a5ccf107c0914f08cc788da55eb179da5bae8454c26707aa767d61f6231fd4075230df44a3e44991629088375d1b8451764be52b7a1a21453be432aac6fd447458a14fc85cdce28cb2ca0fb818fdf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc31d83075aac8c639ae21f6c9ccea2b0fe2c965a43d63b6ca3b09f23b486c681d563f5ddb0cf15a60452291ab4be9968ddf7861f4a9a78de54b037914aedd7b3e113460a74298583f5c17075697bfa3c909c1ec92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa331e5d6895ca4d7da8ee3201db46f064aa624f2200948270026c10a1ffda9733c8521b349c106d2c8f81883a07f96e948aa71ba49077eddfdd3352e48a463c331ca077eb1cce71813a962ce3c6a0863b5aaa2e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8980713c5d18c1f6ead8616dfb6b21f7e37bc59b0500b97327b387481d1f497e4aedc3000693c14430c46a5f8dea3a3c59338b5b0f5e0db9749539f1de08fcee9b43649e089b0f8253cc9350210b7256e09b9fb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76a38b4e9e8cc8d491c58ad63066b851e07559fb4ae38a8004a2794c10699b6ab342563780957174731a17750129fbe9dea3ad72e1bb1276981eac2f37f2b31abab5f20aa4822ed0d7948dbef1d059daab46cebdd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55c1550e820fa8b2affd317ca3b92af7c12f1b96cb10b12e03840ed5af4cc7ff15e389874fc30eb2b51acc49e7c0b8271dbef261dfcb3b9236026b00200d1e8f96944bf0ef0e07a78f2afbbf288d6e7965fc6e7a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57890146fb53f8399127b3a4c3048990b2cc9f1afb92c6106ac889aa4cd460783715cd66a094659d563a3803980b5e9218c5e6f1dbec59fa4027cd05607b5db424f417b3f4708a130d791329962d223c2f90e6766;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf90ac451cad464032859f9c90d759c97e354a219dc02ee2675376e1962efda1bfac5d470bbb1685195c81d932adc43d329300422640f09bcd31521195eaa410830b1c68e6380d781bbc4f127cefafb8d2ce7875dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefb7f6213a81b03f7cb21ed3b80546e00e678a7b0cc49c94de7e83662c664460088b514585787307210f8326fe9f4a9aaccec1d907d4cb6ede3fa95e4a881661de0dcbecc3c72082ce1b79cb1de1c3a78ab90f85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f31527e26b88ff6e2c40fefc6db53f34e667c9c728f7ab08de7d5cc83ea8349f35bd506e5fb43d03fc1d5ce0cbea3a7bd8bc765aa2b41ff7f66bedb81c6786f2f8f202d361cf12ca1b2647f7bb7b286f558a69c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34bbf8cf12eb1050b3694ffc668ac8af8499c43f81877da7789ff63ea94744096d7c44fb8e1977857fa949190f556f913efd43cbddd6306b83b6e6f08ef3bafe5c323a223e173271561ebd03dd52c5de13f14bd62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb604f47efaab3c855ae05871b93739378045593265b3a6e1b13a214de8d1554ee6dc01056c352695bac23165c19456972b214a6a852204167a7c04f0fd5b559015a437455f1f505fe40058dd7c79c4e2fcb538608;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9958606fafc16be1f115950639621bfdbe27afcf440aa47fc325bc05639fdaaab60e41c1f39324965c27bfb333344f50e7a13b91824b670ed7db77c61001ec6ed2e773a6dd65b922a9d23e281b3b87b5005f4f83b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4f8d04d54e3bb548c9b0af8df0e8761f2ae46fffb22ddde5473acf71be37fd5baeb68c72ea35bfc9e35a92a6f05201f35b69fcf749066edc80af29ac0127bcc8f23c7655c3adbb9a8e014ab650b2f7eb46f1ae58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca5d1b193413aded5b051dc2d59544dbb91912645382750087a13f0632e7684aba3820eb374f4b4375c5795903f0f9e0e4aa0f68f4cd9bae76fdfabac5471cb32a262433495313962b1f68c6c7acdfc5568a914bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf622971ac53973aa193ed918813fa1163f2d4d0f34d70a5fa51be750896107f8a8d7a77ee1c021f09089081d2334aa7c7bf16ce0cd845f87aaee9022074016f5dd18d8945bbb241740c6df7ef1d3356d70965d8ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5ae0b24cc4ec79204636597e42eb3eed5446a7b1cf4fb569d914e19882532f492e72e2959aa72e74a8d2a9dfdff81f0e8dbdfc0c933ef67e683864afa50a61f70f8c0c59c806726d297eed7b9891afd5a2e3b0e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he24fc26b74b5967a48a6c688b22d73ce60c72a7e0b77d21083eda68c1ae5f3ab8e9b615785098403823ad40852b1a115746352b708d344c810dce520a2b7b91fdb0ee2acf60d8951e3eaf7d257d3e2da0d7d6e5b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f14f48b4c86cfbbc909da5a5de50b90338bcd5f5fee3f8f49a1215a5c950b6a388176186e0562884b2fdf2977427c24a9f9d364747698efcea86200ca1f5f4fec12674db63bc87d92b0e4f6fc7f3a0aa474e5d88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0b0fd81e3143565730bb241def7b8ef556420681b8cb2eeb9a48ed9b5b3336cde185b808960837680e1cfce77a1dcb9d336dfdbfcb97b95c56054100523b484ddddffbd8a3b1e33ffce204693aa71ae16ae5faf9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f1edb2807b30b31c3ad9afd0cf0032815fb0249e568b9cb46bd9aae4249ab8ddc4f937234ff8b2e59df808effd58aed14273f1d41427505dd7ce314a136c283dce1ae3a50ea11d2989da0f3cc8008707f1e9caf6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0eab7429dbac35c3b947ede4e938b7e9588f21d83b5cc218436f2bd80380cbae6581b532ac456114f99a47bb46b54fab23fe65a5e356ccec53086cae9409a6a5b45d0be50501ca8d0f4ea96d131162298bce402c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4d9f730ec329f573d87241e18dbab0c6efa578688d47f192363a27ec4f78deae42fbc5f34eb90073e730a5db8ddd24c3922cbbd544c64ae0eab027b04046750464232965ec5e6ea64e7216dc81c443c5e5881093;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6b7d854529ad204419204f3a5b91e278d2472d973f07ad801d88092306c05ea850579d974c8bd2215ae72f688321c620d2042488fad810a0d46e40036f1a4e2fefdc7df63d3b7dc78fec948d4bfd88c3f3e0e87a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f24f5c3360b53569ef4dcf3896a59ee5a488f6caa4b817147d68aa829dd01a8904fe81c002da86b38e2d43a3210b3fb0e7c0147d9a6a5d14d5a87b8969be0b1c32afd0c22af0b47501711b8d2aa1ecfcd451d09b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0d95c2a577c9f01855759c6c2e9daec59fffa7a0634e0ff7379bed9575b3b12df7368b00748686de5091b6fcac261aad5a26405fd7cac3edc555a960dbfdea54b04c37036effe933a2b05f12037533992478db48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b65ec2c4c1f2710e6eb1d9cecf1b9f92775ed7141f7cbd23d2692a0c941189be821bcda64617a6b1146a82e546e0e5b2e17093f9998e1bc0ba693f29f901c09d9297260688247dbb6a9ed524050bb411ee01b522;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7fca88e34389d6ce30801f25ed632f8ce01ff4327aa13b3e64e6f43e3a18c6997a825d487f708db2ff81141ba8dae40f14a7b6e65f24ce8e71048e721b220912fd12c7843a3f17941898cac8473bbf7641c3c197;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d754b0facc17987daec4f85105042397f952ca97faf749443b075522937e9475dd1ba6672649ec1f35eb30973abb19336094ff3cf36cd37276b06d32127212f7fd5dcbde852956cddb9e3fbe25e0d0489ba37c2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4737108f9760deb9387517776f53b628c03ff83ccbfc92ccccb03a2f315c68b7245d7a0654b73deacd40c21256474d62f3d37686dbb00ad1bd0c87bed8472e0a0d6ef3a024db8f75d3c1ea919479b7738825b5497;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94ffc6d85217033b8a4b7c21b3e7d65cfeaad8209ffd2e13ea25c659ef7f459b5fa3f9aac3a1468314cdb625b146964f9b22cd7fcfded86a3dcce9ff724f0cb2f1050bf54c7a96c78974c138a921d981b9f391f10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2f78ab1282b4994f879b302dc2ad64a5056f71a1d587af5e68b60eb5f97fe194455ada86e15209d7e1c27dd4f8188c8faf29005e534c285e105a8ee6f9fe850850480daa92476aec35a6c31d71e8f9ede6d51d83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12470376d02f3d6884777811e2803d65b306cac6a903f172e309d37da95e0a10b4e37af9cb60fa3f9e8c4d654410e2a4d001e29b4d5d9e8b9d6e9f0b2bf2585e70419981a88b464b5fe274373489a706f153ad403;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91a36b1760365e1f5b3da5dc5afd702df2690ac3fee39e3cf1acdccb4d5576663dec43a7ad994863c84fdf6634d0b8a094f3a73bfaa855b48ef5daf82b8394dcdf49e9ad93838757faea0acf8c09f11884fbad347;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69991ea464de3f6dea1f08e5f18537e67cca82159eeb9fd8ceca21dc526d840d06878ef7e326861c2d4d276662ab78066f3dd7c45243602ac59c5ca92c6d9f382600f00fbb93254f7075e1fd628e3ad333022f791;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf44079f51f12debd66ebcfba8571b6ef1f50246fb7dbcf5c6c3b3b0bbffd96c454619776deb620f64d0f05b5d049a5a6b95f91f5b9b5b489023b7d09ed2cbf5e4f0d10173a98c4bcdc7d885b78a23cd75fe9b5b24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5d4ca3e84d0b39b4570a051c26e3765545af308365d9b13021d5f206bb00ffd84bd484835bf86d78f4bc6acd593837b9fa5404913d2ee6bbcd5be05d5fd16cc5612f4460c4d5a901526cc4f2ec47978ee256e272;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7964a016970a54e6369988c03c88f86659367a8b30222390afc15136156658fed535f416e821d102d0ef59e9db56e257d7fb08d6cc61d58210ec59cc3fa146f0348555ade242ddc5bae185e7911546f6982509df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf630e9f43527c547597f02fcd4ff17507c45dd12319e315870b29dd28305ac88825e727a0d84fd32b2181343f02264443394a79b1fa40b55e205b02e3012ef19c22f11ab8bdf14085bb77a94a4457edee7bb9c8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7da12d18a52e179d47947398f1c9d6134814c5ba110c29e73b82885623a36fc72c9b530565a02722c43f0b9b1ac1a2efb0f5b33ebe68a50c7c4c913fc68529baf113fe83a63f7678fd870d7c5f28a42f9135bdad1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he54a9e05ddd7cb84a910806ad178a2fd09efdfe1096885e3530cb54210d664378f89bbe96bd1dc9ba26b53402d910adf7ea154c5cf6d3bc634fac50647fdd48ca3c9aa256e3d2a065356ed68eddc6642a5ca00ce2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c1dffc6adc63a735bf9193e8a185e0588af65a208374f01b608075ded96d6dbf3b4b0873de5c32d2d4700b4bea3ab84804c1c1b6338fb286e4b407759e0b90990f5e4d596d2da3236d0832b10a5d82fc72e01ad7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6184ad6758f5cfe133922bca6d3e8e6fe16ebba872515fffeb8e8f9df45e84886336837daf5d1cae1d335d06c7a34a0a5f697e86cb3e6ff5b052bb73a64393849e3b6bcd825ad270e6b040a01466d463332aebdf3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b90b3830f81280b65892ce7a13729af18ab052ac44c3a60a49635386bd1cc341033b376e48f8dfba7ca6ba0c7a940ea687f648d2e957eba84b23054b676d83454323bd332641c134bf3a77dd3e9ef92dece1b2e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9500a9932b8ace9f9fc778eb1bbb24b7934c6c828053e5ce9fa9425056e58dcab2d684bdb1cb6bcfd0d07919a07357c20f2639add541504775ab0cd6a8919f817f2d3ae0c8c703345d787df1292c15e5353054b33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e8a71e10694e3c5e0eaae4a9a59110008515a076e9b1dbf84feacbeee269391f352c9b35b6a09026085b8d2a2abcbe272bd114387cbbc69fa8668b9cad11f652241337677a1724e5464509b26cc81c47e1ada0b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2465ee741f28d061e65ec2c7f784a19e2b85bf7282e53dce3e49e3868b092c43370c731a2ec8ff5ba98732331285e4b5c8bbb79653e7115fc5a787e083a05a4913ad28a42cf85a7143abe2363ae30d157bc125754;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8a64de273f90d513f8acc3770adef28638c74a8e62a587c0ec0641550eac9fa3fe7615a9c73dd64ba7bf6a0bba3fac2b20f77b37ea5c012aa09f3bdd98b5f740d0eb4ffdb108a200bb8e651ecec89364ce428f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf36ab4d910924a8610a26de230d7317367f6c0f8ebe4942e042d727bd51f091ab1f9fb6d0d77eba1e9c3e2e52098986b3e875c13c04548750761fa0673a2b01745304d202f9305171b35a5700b560096f9d86e6ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ca6332a612becc886697d7c9c9a342f67be70fdbbdf8f07127cf3630e5a54689b77f9acdcec8de5fb1340750f938bb1db19ed3e70384a2cfbd6721eb53ced29aeb9f674a093670098769eb7888c7215104c5b2c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfbb3392fb74ae70d4fa6cfb44b058dd55fec79446d465ebfebf80989af7cde89d6aff52252c1f722881629beafdb7ad00c41b42158325e4331d2f469f3700ee212cec3e861d6f539a075d92559d1ae49b34a94a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1932197667b77dc6531fec8ae6173b0e60d01ffb66cb9036ce20e8093f3919a0d4377c555831f35b45372e6b02b6c3eab583817f4d17fa17be928c211428fe06134cfa9f846f6288684c6b7128f1dcd75e5f4d75b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a9f5deae3321c7c0cd2fd2d67e822e65d5bb3ff45d409ea0edf328cd9fe22ebd0fe8dac7e305d34035e67fa6625a93a02443b3efdddccd949b994e7c0c5bd0b0f8c4729e403f9641f93f237bbc3e3ed58920e2f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb861fc4231c2a473c3b0817ba1fdceab82e7509d69d34fd2d225710d7b293185b3f1a82ca6c8ec85a406aebaa696f887c80c53a4a551b13642a5e3fc7f0a2e3400fffad6292f0c2fffa04ed3836a94d6a7da9fcec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h772dbe4b2d4c68cbf5304d7aead97b3db6e867657e07b0a0f4acf3395899183b94f75824b53e0cc57cf0db0b8b93b347f6d9fe8ebaf95ce9c3960c1d804f77902f92f26d00a5aeed72fe4b3fb6cb88bafe8a7b1e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f087cff5a0552b05e8122d7a1ec79a77e60ae253ce8873d5b8d87d5a7d53140c7e8a168427e205b9c5eba9ad1ab8c3a18ee1657159d682973fc07009cabe71d0def4977c05d72007971c1703c2abbb2127e8fef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c45c2bfdee138944a734c869883b3f4e80346e15b084dfb1a123e11264702937d9249569ff88bceb6df63c452874d54369cc6c238e822c176feb0c23691c6f460d8bac5014df5d9a6089c9b29ef68b71a604c463;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb393720d4fd7e671ce08317c61cc05c895cee7a39fad1b16fdbdaf1ba72633a84b2c0ac321e3c42358eb681b1d7dcbe550df32061d657357f134800e81b1d11b5d5deddf0613af86836a49c4e1454b219ed67ce6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9704b9299a4c401b2c5d836b3c585757644f5249bdc3234def51b90a7e52750e7f87dfef266c9574a537d33325c47850a06bfd653c81d2aed1945005ed9980a72b8bbff72f6021b76a2b3bde2e05d6cfec17d3783;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1058f2c60f1d4fdd28401566082f00a9ef044f59e9888a35d764ab0d44732fe0d57fbca9f9878aa2807813da5ec48fa4e7192e949cfc33cefc222c304732326bd57af97fd69aab2c46cb081e956b2112b3d409263;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8cd28a7b8e4f17d71925d01c513087acee7f2d6700f982c8711092d638b4a6b3a7b0b41e626bfff2dd15431c1664aa777842e0380caf56fa667613a08de9729220d27e0d8987433fe183214222b81e3e08f70d40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h248f23335144d5bb5ef9729bd538eef3071ed945aaa3d26557925ba5cfbf89d5d8574342f35699e8acc8afcde2b3cf9cc07e7a66bde2f0563c41faf7d0860f1ea48d867c1c4b93ce2a4790476e97fc89650cfc647;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ed146a03506bbae7f3c1327b53047ace165ba67e0d416950522e3c1f69885463c552d6bb9e56d450d6232072a1e65ddb1babc429e575ddd5c011235793d2ca8d6b5bf2e4ced80ef6319a1e68395a7f946b52687d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83cacc82acbc8cd318666904044132bd5f72156d8fb3e3450254482acd2dffdf57cac690e31220f879feea4bd587c9e87a6cedc0faf17df917a3e0555259dee82a2e9c3bbeb811ddc95b3ec4d90e86d1c0c001e53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b6500784f508c55ea9afeb0a09f9263d4aec0916eae4892566fa4a025d3ac4457c03b41363f3a497aa0a711be2769341e6ccf6d6224a8e18c211e3ea7b2d90260a2b6e390de643dbdb37323ca4bef2f13a4e73ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac49e5bdbbb15d325a75ed91ffe953a128eac5a6ddacd880217b4225eabe38635ee0b901500000598cd1808c6f556b955205d215c942aeed8e198b24582fd92842469b1d636b77d15cc310e7a4e8af0b0e6e3a994;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h263dcac94a89d2dcc097264d0d959bff8aa456b69e3b74df695a7d4062ac895e64bb03d438ed0dceb5b800c06f5034e9b311259915d97d17ee1e19f364691687b89f1310939f0375b8025935cc341ada96a35cd59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h979cdf104313866f00c2e06d1d0dd323c94dffcc7f1f7435bdf22bda330a98d02b6b41bea75f2d5e8b81f66bd75610ecc445a7080685309bb3e86ffaa26b9516fe0e68842dd6fbdcfe008bc01cf5272154f6a74e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18beb200434fab823859d763b39f427cdf53176c5eec35a901d1c160b80fa5e83a22024b4941be8677e47f29ce0e44c84656cc78b12b90c791a7a859ddbcb4d76305d0313bad45e22760b902e9431777224f83bc9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ade38ff4b932b2b68919794db90920cbb2b05e8cc90eba1ad4f869c4c835c08345c75e6a502ada0716ce353301abb676f5e6deb0dd32952418974bd9be9970a3865bb6e4073a6334cfa3144587ca1a073b1050a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfe2e125c4fabd4b4e48e15d966bc2da9e0baa14f8834cf395328ed76f109e65e60d2b29d6505058bd7dcc184d0b2afccb79c6de09572acc8ee7c5487513025ea1d850f4749e4febc84a8cc1a850f8a072628ab83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf180b4844be68b430ea298e25e61c406342f790fe09a8f1f3d526a9ea4765c79745ce419a09275803337d2b6183720bb66a5214e3d713b4d1489cc799bb1504e7398ca892d4dcf7cd14465d482006b110e95d346c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb08b4bc2424cfc51b7ccd195846a6ae3501bc86eba400f870a25fda6b963c3f73fed0cd996bc420630dee130baf894da81bcf9ee9a38de7b4f799010e2bdce83d7491ddeca1eac41e1e713a4ccfc29e5cc0e0a431;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52dd1570bac043139e627bf28cf1764808fbeddb6d5171764132fa391267d5b53fbe5a87b870e2c160c0472279ab039889bd3004847e18025831b7745da6e04aa9f6c507335be032528443571137b7d3a017794e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb924bae17ebf1cf1d3ad9dfc560547c6053d0ee0d3bf0b04c2b9b5e5c234f15af7a1f80dd59b3d0c2ad3d4537401e75ba76574a195c34f1377991c0e7432a38382f3875f1fa74bcac5fcd437a9fd40d569f85f8e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf866b24d98e868bfcb48b428ba946ccac56aa5001a931eebb91811972a7d441365c5c28f9a6fed1496d228f425c70db6eb816b1d77b1d80b3a390d72bfe2f662c169e645d71144fea78bcc2a16511cc264c10103;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74b38918f2d4176323a30be7c12d76f10535559f7c57da582f4d961f600acb0c0c345bf20ddb6b743752c9a9ea03f1efa7e3dde7b78636fca2195baf0a3f6dc4205d64832778da90fa7c61dd07c40719e336587cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e9d31bbfd2cf95ff5fd121b68e7ea2082364d0e4ec73b67650e943edbf4765192778e4ab22fb3af0e53d4577bff29e9c9d86657c99e2a0182ab4146161ee4cd9110bc6d3223958a65316fef50d33c610032f7469;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h500f062539a06b1736c5f117a7df4fda914c59b5e05b818c7952d4b744e75bf4e88caa2a27d45f92908191e62e93deec68d21f74a460b65d0a0e2e46c77fd490ba1112524d9049d3e9675075cce0f0316c38668d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e1f5ea7bdf38b8f351d80b675ba0b2377ee37a0f1099447d391d6992a443c38b68d977f2ef9f9aacfcbe5d8796252110afcd8b025208a4e13c57218af273da258e8db44b257b25b4bc387a224d46070403a42047;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h111ca41163033d66c0ff1078cb5fe48d2d3a49fac38aee24958e53ed8945fa98e1001bae4840042f35a0eaedb81f10602d460e6dd57bdb30d42e5e9145684d4e788e87a9d58ce6720b5c85dafcf56d51582b6191a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f7501550e4d702fed13d0138142b5008938e9af789bac2277c3ee219d74c12f6ef1b0963aef45eac5ef620b2478064a67cb0dceed0a28b973d0f8605b50781fd93a95c6c2d0c7e4953b0bc10df64d0479c7548a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0b979065f03a56b9c1fbc84d5bfea77a0dfcf21f8e5bb9d0e5449f736640aa5ba1e0fa9df515848a4602686b57b46e1d2fc90acb5e7d681af3e2a8cc02f88ee2230843963b53d28a8a862dd7b5bba824581a4721;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1835ac85ec22b7c7c0b320382eb60efa87d37a2bc3cf08f81c0f450c656fae9827405644f0d7c20df92eb7c770a4c9cfdfc06eba65d417f561c2fa5037451a2b9e31bb624fe38cce98bc68da810a71164c7198b64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52538c6e1cbf01ae8e7da35c10790d5a516aaf1ec87b8bb964658c9e9538aba44cf62dfd8c9dfcf3a00eb9d6596c4fad6065be9a1254a263fd9039c037536e399f3cc987801dad2ede2586d1effd3542f4206876c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h707861013e90335aec3d8af49719d944a8a1280b44a1c1bd5f6a31b54945b45f5a588ed20302a79cf0800b0cfee4bc84dc9e3f59227a8f205f58c5cc4e2870a75268eab78a94cfeb5e72b188b5450c60241fd0331;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27916e254d8646da4ae4b56948b52b700b3dcb3a07fb778950631f780efd7c46f96ec4fde9637fff8d63e52397dbbfd79e980e279c47e7d8442ac2adaf6966f75d986463c96d16b5c468cb135d5240e450e157ff2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c7881b4914a12189544226471c29084588f08974084c353c3d9bf9edd8eb64825b4874acd6ff0f49d3e299464fc0619a392ea96f18f67ff1b2eecc05dbcacf69d5fbd0d0372af7147fa5d7d53391976c9bc8e749;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4080bf818334d041e6a20bc568aed8e30cae447853e5444f6c6e46dfea97624a89842e745c6985e4047004175376af3631a88107212379dff9fe00a879228c55d4ec1fb1acd2b390712ab035e8fd6d1c527625018;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65f26c7af80e426006842f11154187c3b12accaea8ec5e3f3b8a7982cd0220a8aac90efdc03bfd4703a4698ae001bd7e7081cb0a12faf7a2c50a59cfbe00acc801ac1018556db840ffc6d8d2e856c4eae2b4b51c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdb4cce56db2a1949b195df43f35bff0abc8f4f27cdbf4adbd3ca87fa54f19f9a922c23075710e4cb06c617bb430b763310d9c79bfd1d3fddc717bcd1ae509b7f9c25e10941e4a7bb5d5cf9d8bbf26db1eb8c9423;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c7ff1ddbde92532587b0e407e9292389f309a14be4022bdf36183e8047a9115384f55b14565d77153edf2c0783c5ff2a14a423b44d331471b45f3e77a5b67e290690da1f274b5d7dd300b3465a6bffc65590702f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cef521b016ecfc7dbacd5dd290719f088e7ad7ce97a2ca7fd42b80af7b29227e6e7340d1414475d56462d5f9f5d6c719eb4d62d5f01d7db70d5e40e7ee09d62f60ce5e82d95fb4a94b852588d6ef7a7605dde174;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf50e4be7741dae0d637af0306e0a96607d91673697cfcbd03c0e08d66583230f24f2fcad86e89b79c23ff50d9ebb091f2ebe202521463d2a585fa6885b6b3e3aee75bfb4621d18a12ebf9c923c708749b9e601ad0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h534b0269d18e22be29d901b25e24c92d461be54735de37adb0c2d039d9a62f474e453a68ab39fef4e788ae834abeb5a6dbe1ad1b2d47691d6e16f90065b87c0cb1ebdbf78cae47d6bf996349594f46360d4bfcd3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d1164e2e29d9e04d282b36402f75522a5654a16df823dcbd253ac9257aa44da366a2b5b2022746f18d9d0dcdeec7d549cf94ccf6d8525c499f01ccdac1af6615e41e36fd14febd68ab8a47e1f16e78bd7b85dcad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h576e0dc8f82f14c2086d6bd9e57c4d2519a4e46be85f6c3203584547a1264c6b92ee36185f51fb4e04a1d00576d6e0e877d17730b33955996b3312a5a0ff3cfd30f13aa6034e4fae0d7e4c63b4ef6017789e8a588;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha561842d910dad2030dfcd306609ba732849a2beaefca8ff76b326498ecc26ff4ce02c583d2e033e88861b5874a43a177a3626b3a939c03ad0710f42be9668db3861a41af4bad2d596e4c182944927d3c9a285de8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe6a535e668ab9df4c8dc6ca89bcf1e6a4cc83d680d87c15083df2adf6a38293aa3644eef2772964a2dce2da9be86463edbbc437fc22e7a497fad4a54f610b705d290e7095c3329525fb150fd6c130a006a34f24e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36fe1760c7d526bba50e8c4b2d9e2c55b484cdef76786587aaa904554ed4a065721c439d22749efd6a31803e3aea9c25e13b7d12806e6fcaa49e02e32182fa1f99045e915eb4d115ab5c8632c36f10ebbe90c4dca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec77de789f2cc695f173836047624dd35b2e836be7eaafa2b5d1de5b558bba0eb96944bd637229965c9acc2d37ff84eaa1ebcee8d7baa25f2266e7fc0f9c27d101a875bc6d4593761103cb282ab0a08d8bd7803a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61f245d51494d9eee5a02032f49db95537d9482da30de606db6c8dddb643d629c16a5d4e7f59b2890adeb2c3ad0af60c717361185438ba30bcbc85a67d02f86bcbda15f4372d74c944f3abc5e6206a9ddc25ca075;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e9c51f018121ab6f4428b8060de827eb46cbedbdce60daa5f4ef4f70cd99bd8a733d083a4a164cdda0ad063d010ba31e00395226cdba6a1937889061576c460c1095b4e270b73f9bde93c479ff8723756f92dc6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3237cb4134249056ac6b77e0d61ba095aa8b5f74fb9f4dcde8c0cb122dcef530b732c7ff0f184e4868f47547ef9c86b6f23cbadee59b81edd081382b64a748f5d8b62f435935650d4a6666e190f15b648210f7ef9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab483d201c46f60d30a290e563bad24db27b9c92c2a0603e4556f2663a80676780faa916b51bf1e0d2aef01e48c11c94cf421e7a7eeb3eee21b92c787a63d37b0b320f025e6e9676a2f8c0a90e78ecfca6e1afe8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h648ee0b20982ec99d93966d06e791e7262642adf3f7817a6bf0cc51217be9b2b615beb32ed2daa09f4a68b52624aecc63860cc1e7b951acdca4149941e6bf2aec7810548a07fe360d85f1d1f7b05e64bdb410560f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h788a1e2aa1bb7fde9adce7c706786438e7ac61b50a3046ed320021190ca847552f8741295d1a7ba1638dab2e0b432f913af8fd424283919a6926a5484cc9979acc733c2e60a739fdfd64335cb9246ebe9060a1ed4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h555b85391ebd8e5acc9f6e05890751b615d867d668b8314e44ae7484a57d4b432d8eeab06e53f53d0aa96c86ce74c84c38452e2b8e4d5a9cdab3b60c24e5ffd04d740ab641f33199dedc979f6dbd5bc6ad306cea1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bdfdeedcc9c8e05e8803e535ba3131128938226073c12aec365261d99fbe85ff22548156734014dcb4a5b366f41c0597965269e6ccc3d2d77a16f30c2389b2bfb696071a7d7c4ae434d0270daf0c9f0dfb4fa157;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba52e089f3480fa2e202e5f69c9bfbcd00ee149949fa8ea9f7898c7b5da321a5c0a91fb15312682f48d5e2adcc032b6ca678d88ba3b098454bf5cfad582ff53ec0324ded135e7fed118cf9494779015ef537836;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3529be229fa03627592f027de8d309a01414080a6661ea8eb0a9496df278e2b3f61504835cb6958173cae312b3f8bf3fbc3f69b72318c56d4feff030a96ceab0a79713fda64738a0f817ae1155c5e161344152ee6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab4a5d26272b36990487ca35d91123d270c4350f289a0db7ae7acbec362082e5980b7f1d2b89ab43cb049c44dbbf9a7d7933eaf7879f55be2b2a4df18cd3a14e4fb192f8401eac38b34a5342c05cfd1fdf9bbcc06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3d32e92c9a0ce1d9595667286ec1808bfa114edd13e270be43cc16ba4dc18471dc0cedc0cf62e0645e3ad52b35081f98c2c6364b09d5accb7cfaedc94284bba82974e9bcd81579aeb9539b50fe13043527e9967a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf627513d11ffb1f9bc2357d59d209aa99931f102da210508af1df638f5d8153c98b03b663bb5917e0c1bffbbabb725ef7f0fc56e34bb0930837fb1f2576a86acf6ca883089edf5a3b65c7db12c8e43475cafc6cbc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11a9802806c9b747643ee47e79eda02192a9ade5b7cbf55776364d0a1cc9f236748db8f874c1b84c50becccef33b07d39d43b4fa1f2b373f12a9ab6df29f052304490cd89f082a64154643b349f3cc7f39ab474a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacefa750f2bcdee99c5c50c52110b192187d9f99c0ed291f56cc927e2bd130dc13c941a5489066f214d9f90fddd7d698c78c4122f5c869aaa677790b92de2e6065de0e7dea458eabbbd7f5553d051ae6c9396591e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3ec4b9f86ee1804d4f83a1c2bfd1c2e19507d13c50577a06e22a0c4ea27b1f6db7263e0376898b50df178fef687f40c6d5620763fea518ea81ec11def8a68e85dd8f9287e4075ded90906368a942cdb9b1c10e9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h475c0ceed7f29283423ddd2ff1088b9e8d0410bdbf28c9dcfa489b771d3d92a648779ea552cd0bc79529973ffe034bed6f1e6107733954d600575414586d72548a60e80459c9764b38eaec0d82553e99dedea9b73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6494fdf124c1dd7a9ef80e771be7b3ece2ab36228b95513a42577351ee5c92fe622d1e33ea34cc29e8b3c64866accc17a7f2b9395c1baa017d9da6f11998e969b87a0c1213df60e37e29f0b74a99cdd22fb34714c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c9063f3f3347abdb83eb6143a8121665c14580fce8a0ffe047990c8bd4e337fe2cdc55376cadb89562991b792153f155db89cb0a30d2001589b44ee71f95f57a9fd5688734004f2df4ff538ac82bdece3bc0dee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42fa5859ed63a91b22f9a15f68b57ef935c21bce540a05e468a657d23a099a258a391c8d3c884dcfbed4382419c8070e02a90763879294fedce1f4eae706f7db56133cd5c54c538e1e2aa9e89db7a24988a42cb0e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hece139ec24d1d6a8d3acaaf25dc49d821de0cc050d0311dd3f62ed4010b235798bb0810aa991fefe20f22cb61ba2ca68b09b6535bf9e2d1d9b4baa4e7a086682ebc72a1d3b50d26ee42523e25d2eda14bb84d066d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d5aa7ef03e11d02e0573b31747b08852c40c8f9077190b71d9b20b936b7bb90bd52cd9d89a35429da8cadaf0364f02f5581348630a41d9120735f91397c3e7339f161aadf09da84c7970031a7439f8c7220a739c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h184abcc219e65ca09054d634efa6b70ee177ec4039588babbc523cc586f43da02bd1827733d3c82fbf18d8908701ace884fbb11e98f4304a91f4a48db83b5659c54653aa50afd9905edce89443a445c30f206439f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4078f49adba7d1f72105fc615883c2fa6863ffd8920840372dc747454529f19549ec6d00e245141c21b6c0fded9bbbd905b0bc0061a2fb7308a92976ddc70190f86124b35d619d13853d5d061d284bc1b1a46211a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fd2cb266e65bd54faa0b9f349ed0c820031f201affab18c109773f5043a91b5e77d6a49280406e02334bf00e6b85872a588c3fd361d5a90c1f33f2dc869d20b594f6769f8053e36c6e0ca2b4a2e85226c79192ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42910065c5f5b591720227611ecc74f6c08730a0f196da7c37ec7696c65538c0cb204cfd0a456bf1907c063b1abf1cd28ff37bb533c959dc6e4851b47a7ef088d6bf4b2b8a299098e5db6ecca798912a6a6af8125;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7158def9dd21eb533ef4cf83f94d79f526424ced29029d64bd3394ae7dab57c0c3741a7e6193391f2b853c851b8d1f258b9317218dace1cd730a47219a111e03faf5547be8e90319d1ea8e4fb828fe4adc04fb709;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a10f29c5329599c91529976f57357d7ce18c63254db12ea7bba5d2ef8f75e41d818e95b3a9b738eadb2ab1ca4f52d760b6a4b0097ed237a8fd2087395e7620a2be88aac43c4b2fcca1b61aae401727e85106c662;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3c4742453571b265a2b793eca4d56bc20c84dcffb873a18211fa5506379f5cf6f111ea5e65074728e658f28083405ab7e17a50c834139722f9b207f488c5ad3e7e00d4f7c8e17fa9cbd305d0d597b9761b00082d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefe066952f313e7207bf9554910af0e5ac768d309efd33b692e71338e8531ea2e850a7230c21d723fadecb538826329f2d535742d017d39259f2151e814209dbab61f535f9f4b0d066adbb392ad492356487f6f4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h196361fa8f4b57235593113e35f0d0aa1a9e9420f4e5a807f434e4fd4e02c4d9b039ee7ed52875051f6442f73f2b95c3329f29d0ca8d561de438ec96a43cde5db4751cb8f7886b77bec0e45cf7816577506299fcd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bd8e02f8d281bb7f677cca0778e56cb745099dad95e782892751816bf9d42b76aa0287ef89a453b9e83bd3b289069c67c4efdaf60f86897f1b36dfe0e4dec7a0f17846a3026488d034150f104943b75e5f138990;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4ef0e6c2fe1bdb75e1bad85cfcd27cff23baaf89285e3c4378a6336e74988ed9a397cbe0c5b88c410d7d3ea544956f983e6ae88a16f6e6edf5e8129c0b29c3396985b15b0a390077aa1ef3e26160070a27df3c78;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14eb8278fc6af3e983c62b2401e84f341128f8f625c015cd3a63de2698e9d2cd25440971c4e895aaa5da9145190841f40ff29cea92d02fc1e4693599e33ad3f626491966c08cf722a090996c9d95dec8fdd598bb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fbac5761963bd05201a583c17a235fa5c72ec8db85ce4f3c292483604491296f3cb289263c40ea5264e7bc8be315c72fdf6fdf9db6314d66f61cb89264e70a00a2689a183b98200e68c18e32aa663267c94ec9a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h772e0a9f31403ba23c9030957fa11e506c8502840ad5d7b45b03224a0c70c036ecfe4cd033ef949d86c50b573c70b4d458453e009bee6dc9fe5cc22cabde79ccf15f7857c7956cdd908eea6af2d4b66c067264830;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25a9660f4e72cb7e75e227ede76ef9cb4cfea662b4bf19cdaf33bc97b2829ed04bccad0f8f29c5d63cd466c05d15f31b27877990a229fa800fa1c68d10a6eeb21cd152ee40ebd017530e67379c7857f64c387e506;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c99d5f30068e30db573bd03ab6e1a91f6536f6b9096c8050159dd9a7efa8d5e1f1342930bb77d3401f031ce60699c3db610ab1e8e8be861f963b4f242223dfe8b631fd4d4da01ef155bdd0c2678dccf3117b4850;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc282de335f8e653e66f05a2631a6d951edb998a3993e3bfe37c690d01e7b88f9bf79987b8781aaf2b8ba9851466f6a3b174fd28de5c0b30011c4ce09627c8129ff66cb7a6fbad862c9cf715cdd71657ae81dccb8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85c6cf092f4c02feae28b2c7a831436d7005a9b6834b9992c821bb714fd78ba84539cc1fc2d46a58a7338e3623f18a40fc0a126f88a4051fbcf5d5860c48b444ebde5a71fed236ff50b0bd77d54501015b3e8e1b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbafadca374ca27ca916084694442a2f36c560b70efd4b69e40b644c41b9b48e38d7dc7c6913dfa092c3d76985e7012c4b0ff339a1097e526a8cabfc6708a3c33355c697768956b68cfdfcee30028dd03fd60c4a6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fd43398184bbc4693801d014aabe2faeb68ea4b27b72df8eea6022546516cd67842132610da292f81aa263c40ec4f747d2412c871ddad36f508a291e4cc748a42b2345b1c1a93ed81c24cd669895618deefe6a5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f64ff3bff55e5f923dc1cd4b1729605632a54193cfe5687ba1ef034a249708f12b26c9595c13c685c16e7889d910d41584a0a0c42f88b25b5d25bb83fb127378a51b975f7f64a1c76ea5c214c138d2d626811930;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff5ca403ca4c4186b2037188107dc562168b4a3752b331660cc8f4887f313f52d90292b54541e9c910c8e2bbd2a9bd300efd949cf9cd3abb761994464a1ac09aa9ce3b27420aaa97efa6a9ca501df838531408b62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd692adf037f7f5111f068c0016357223b0863633979c99192d610b26a7bccc4c0f075616877902fe3e4565f3bc043a5194ea296951f9e616fd7b92c864565cfb9806d993b3a22c371eb2964e0fed4306344e143a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97e05f223a9c58a5374fbebf0432b45ce00eb77c69123ca28ffb08cba9cd5ff92d9cd23c665441a5b99a607f7c7c579dcd5ffb57ccbcfe118fbaa20951586a85d160646d86b6e483be88c180b9c6dd8260a921232;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa94cc31db5700df338af6d77b9f5a13bd77460a372527ef3e85fe56739a28f7b13a8d63e7b3d61f987b8bb118c4db8901ec6e8ea3516c792bbc0ec5a8b5202d55875cba61a3ce0500c32ec593391af0f51d42a7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef4727a6cecebd940f816984367494279a7afc5574010958047ebbf6986d27407024218e0dfe1a45ac8197d6bec2b4e40b3e10a073db2953cbe155903637631d676cb764fe862560973db57bfcf0a675b1488ca20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5d0483c629d2769ea06732112250338331c9dda0b741f6f694e57da017ec05c86afd0f8b08fd97cecdb5af0a7b34de0750434cc572706beaa19faba43005cbc6ca3625fe7dad11eedd61ef1dfdc450a77a4e8933;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf248f9f9905373a93565002938cdabec6664d258bd69ce16b2ac31bac398191d2abe2a67a64ad8f8cdb2fe30c5780593767710edb13464a17223f8757db5dbd7174a913278a1dae932a9a2b048bf7f75a2041ad4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96714083865eeabfaf1d196d3fe92aa2d5409dea7e83c758c5a4481224e726b5e26ae3a8787fe11eae5fad45dcf89274cbe70db57642894f1cc7fa8ace728e915085c6fc5883178f04a757ebe787d3e250fdea653;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8de4ee0f7ac3aa1e20aef917428d8876b86c2b320b88f61665d022e846707e5ffd62242e215466875f233f9bc524c31f5dbbceec6cca85e3b714d35e8f6e795c8ea0b386f4f1397b6533d0df7c7ae8f3dd390a6dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf247c014d40064ff9ff69bd2a3fdfca0b99c9c9ec706608c1bfca578e3f6be4401479afb8fd068de6a9728c3be287f191f69fe9ed16d6066ba92cc8cf80e7d1550b41df270430d81c091d4a0fb31119c10683b1db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd70f45eee48d8de3186dd1d7b788a5eb07c875527174c16b8b57b94d8e182c5d12fea805228997cbd4e0d5cd0c76bb8c19f296f8758f40204ae911627d5f24347d65b01e322ad4cc6ec8a66d7c37de4d4bb3097c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he47e2566f814040827aa76fb92a05d2d30b5079a1e622c6c3ae56ffdb386acf822208d2917b77e7efd69c2ea1723b8e4001e4cf28bacd55cb19fe91c1dc316d8fb4198b5307fb267794d6467c56cdf5bc2c1288ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bdde68f08edad0f39b29c4baab3dffb57ed5115d45b28fb626af6c57d578a3edd0b8c412e924bdbf65d66c38da7a46bf747daa99f3b572bad07ef2be6ba2684dcb6c10a355e8bba9a200b734100c82a2b7541420;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f5a713e25c135e77e4ef01c270a3af38a921ec4389698873e070fc81ce2635c7f663fa2ddea41e91551cca7cf934a6b52fa12e3d36d851f55d58f441947e172d9be5771e581953318d3a59928a8b5140b12926f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he71f64b6f8985517544bad55201239ad8514408df943772bdd55c86ec755b4a5119ba29f6be6ebad06471be83ac483177a0bbf4fa5c205adc752a9804b614fdd3310c2dbc6d8f4847679fe9244497c85b8a93914e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he30c0cfdb284008e602782fbe6307857638a4234058848262a2a60a17eb0433e8f09199c8e07e76c154e622c665f85f6b43173a3dcc6094c3161bcee9ee1d0a520e9b6c3666b565eea0a99a5c01f904abf4ff71bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbee807541354596c1e339ef04520a8527c0a65317fd232cf33514951d846553102304dff61b81da2be385bb8d057a5c06274cf3d4bc9164624f5bf96bfe3ceb207403da7178bde2ab1770948d57bad9569a6747ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7eee2a51fa0c7d37cc3376692598c708845ab7d5b59470a0586a9be778f76b709cc82c8df32bb8f42e56b30535223fe49ab9d6556ec670a3582e22113cedf06acd7a4322cd90d0d4fcb548df9e9ed23d36c23eb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he620e743d313833ed4070a0728f28aeabe652f873895b18a1b6e3f7e17831f4f99d0c1a144dd798f7edb8d91114c65055aa03917bf9ae5b399be94bb945da6465f9b62547025088a73a593c5d12f590595c6207ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e686551d69014184dce40fdb63f7681b3781f56ab6e49f4880a4c6d7f5f3b084aa77711b8da132d09494f040ac78dc436c32199e7fd84b9fb5b5ebb7011b1edaa9ddbee2502f018f22cda3253cf06ec5bd2fb69e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70428cd549febe7971e984aafdb6976a19cddf23683a50c112656db6d8fa92389045c1170edc3f8d835fde077e40f53608e408d6511750c516e9b745a6cd0f4a4493fb9c63f9eeb40756ccee89256bd2f893636e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha27a297d1e7fa2647af263f1d12ca7c2d4d1abbc0f15310d517e878caad7ad2c1fce8fa35f5188f2c20022aa9a36c24adbcdd7df9007dab6668d5fa34c82ad1dec3768cae15a335d86f22a2cd89087d26cb3b8c36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b88fbc007e2bf1ee6e0c19496f5537927237a31640cc366e241811a1543f3b94ea017bb4b1a886e43898b65e7ea446876bcdce8d5769ab543ce3fb416384835c8b86a7f4c51669d2f36a478f3e7f86a535ee4407;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9543b7f27638fbbf85291ba91cbd434f901ac823239a5999dc5b643582700c452242e004ad66d067427e7524207a80c8f1d2eac77344b5c892e62e6ca7835f5fd5306b423005af5387ac0f008c268c9dffa7d28ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e8ca5c29821298c7cf8e5bb5e0dcb40e0883b9aba9252f1679f70e7865eb5b2619cd6bb9cff4c3e7c766b70363cf900579016dd64948a76dca2abee1ea4885b2dcc85a3e3af24e0dfad3d8c8139b9e75d804fcd9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9db4a02574bcfebf949bf024a3466ce960cfd111fa76996d46f94a9b64ae788c037d3cdcb2bf6e4297009f50e6f051f190deb7bf3d47d9e893d8cf90253b43f71c4322f52d52a13f9de274004f0fe83877b5d9391;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea34a5380d2d3ccd6d04acd30e7cb64c52e16fc210c4a03698dd7722d8083ba9eeb8fe6915c891f10e1da1d56181378b1d7f33c796d636bbd47f389568eacf53b074102a658cca0a424c667d59c72e1629d85657d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0b4db0cb6e168c3bcaa3b3719396650efa8f91dd2f27a29e60a076cae94ce7f909cec92d548662253d91a47d56215e737ede3a517ea9d257cf5c783302ab8ba31cefd9942d89a0f13d11346f1b06b332ee262346;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2f3a5f187856c4462b6012db7c0cdc0e6b8b6d2bfc7c1da969cf6a82d358219a8572a93bef3cd19c3007266dcd44e1016f33a8d5e44407f1a2b6e5324323b41e2a1eee7a576ad502695075775fcca26b8a19f6ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe475ac854873001959e5225b77527401a5f2bcac12ed58ce0f438d89b34cc87e90b68d36967a0513c580aaf863f67e0f014a5dca19c3b03f20158f95c5c4e6ca928227f72c863626de729954ab409a46355fcbc4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h467d338da06dcd33c995b9fdb8c51dfec958f0da06525d033e56f67c00f9ec6af63ba5ace67f538c6b6aa32c53e32e8f9e1bdf72b43f40cb30b60e2160d2af5e63f59a61fa60a0818094380fa4c7f6575e6cb6683;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h573729ab799d998702f5461c49cf6c2668f60493d5e358ef4ad9e7aa8e0e2e72555d36ab4f55827acda9800753f1f1c50f11bdd6ada0092f23d5183cbdd99b3a81450baeac02b0826e0591472c04364220661b269;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h172cb7ab1843922919be3331503d8b1a756cbecc1c01396f5382682c5f882acf121d24a44fcfeda51708757a49e2f6db56462382b863b60ee1e0dfd4ae5a2163256a66efb067185475ac8ebcd7b9ae0bce62b063f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he465436cf4e31a443bfb5da445322f1d5930bb863976f8063782a96ced24483d3709b525cf353fda41f44101901c498ca921019de85687ade721637d631a9a52cf5bd76331a3476ec7784ddf92b05797a09c63b57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ff3a138ddc6fbc3bd6d09e52fba60d9146bdd844a93c01b129db4823dbfc2b20fd244a3c23cc5bbe3d90aeadf1726ebddec421d23b1a3990047e6ba63d956b04b99f00e7b225b3a42c54da8090e21b215ba5cc01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32fd7495ea1f376bcf21bf28ddd5c0429e7b8331a8ca8a7f4f2657cea0713c9f1bfd5b115005f42112d0979437a76b5441968a55d709dde25d5466e0bbe55181fef0da20cdbd1c4d4ab9ed06552d516bfc97786eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67e2abde3d5ab71eb14f55177677d1732d760e37402467fff04bb9cef3dc04e9c399e0c0b4a63e34cb465ecdcbed71cde8791196f403faf229d80eb7cdaaf90cce9cf1053ea87f0c8a0833c3905c974dd82ac30a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a036a38fc3f595672dde63e94f7f319f0d54266f4be224e22c308b9ad993f2a379b7e17f9e8677c057f6723ae1fc165347e2ec67ca194ace4f1453bbaf24f47de5d3c67975536f4306c74f2940c395c31e72d2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6375857fd6298ba627c1fb87302af28b8bf026594076671af384d1f01ddb72f77ec2e3fe85d625739091595ca3147e42945d3f51d9767940bd845bddff479086945cb400cb6f0da8b1c03c825fc02cdb6f5a2db32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef4e086b763f7c24c6cad38927193e0092075cae22dc9f526369dfc5d4741e8b11b1b18c4006fb5911dff1f71ff50ab62009fe34ca581bd11800e51af992179fd3c4fb835a8bb41efff2fac724338ca4dd200e099;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9258fd9c4257517328f9f9b0463603f833f9e954b67fad5a08d834b804b80bb4713c443b6f799afce1526671ad7af0ef66df3ff753db0dd36cfd06b816e99401e6ca491dc29c5f9a01eedfc52280047201c87db6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d2b98ebdd03677b1c7ebacb357a95a5a0e00e69bbce29364a7b1488fbd7021dad4dba699835e8a056fc577932158c2928df942ea840b32957621deca9951bc5903c5b58820f74b1df9160174edf15342818dd569;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeac53205db5dd01c0898abbdf17bf3a2d079e75d1c020e91c276c3789d54863314ea15490dc33b8626b19f2561e16794cf5809a1010ba4d33cd5ecaf882df07f8a97ecbe39f8b32f5ce1a0b6ceb07317cf586a84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5162bc5dd6c101304f346e7a59d06060e50c4b190772c922ea272bc2ae7d566491da5d18e12edd74163ef351cca022164ac01b1a91b07d9306d7ce317de539cc0a454033d346975c3e3127472c907122ef1ab75e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h140eac517568013b07fe72635c3bb0068bbe4b09e1c922d7b1c703e6b79c66819a9388e625bd53c7cd7eda965cc1beec022dd378bbccb1c0286e1941f59f96e168e2a11d0f3b00625da6cdbc6131c221563617c19;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47ffd123e6d99314e0fbcb85a1b87106371810f82d3ba5006cac405d63ae661ba76d48e1bb4c64838862949e1f47def80a9e9a505724320be3f67c2e1771b62cb942d93df65b6be7aec947b28bd4b7f5fb38a1853;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed228e553f8194d3a85e16a2d19dc20ef68344b0ee600bcff0b88d1a1aef5d9050b72425e272e0c646c0e5ab62b64d7a498a00335b1aae09d8d0b4512c2d422bc978a0379ecf06ac4695ced221973562026e6c4de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c221613dc634fb4a169edc63ca9a6c27f7e4023154ed008a6c9b4c28f17c18c465b4d7efa4b7eec27ab5d7461846216cacf88969e51091f4a4aeea0e486fdc0415202e6009955247bfcbe3d7f31c3c7ce8566362;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41cb1505c809dabbe16e22280767915170ee32809aec403e90fa7a6a8d44140154f68b66defa013810e1e9dd3165441a12efb45de0493fcabf7eb4deb3f8720cbf180b04e558169485db27d89d93468c34882be8f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f09e20cb7c089b836a7aeeac712e56da60e76a553eb65b5bb439aac0e50b9f8d6f388c73f279bbbae42418d664acdedae26b70eba3d1686be47b65fa1683038efc5bdeaafd5ecdf2a934fbcbf4b99a639c12fd6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h113805041b089ca5ba6917131bd8b8f624c6a332241be45df817e4e251dc8dcb4e596fe0d3700b4b5d8794892d4cf67c9c6b2aa4e706b9a464f309985a8ac2c4bff47db332a1134f61097f9df1a663b4ac26990ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h746f5d945cc3554440fa0535bdd746f7abf778b6720b563725d2611b59fb521bbe11812e926ef4d61aa02edba4e27b310dbe6cbb27dd3ba1db2fc2fa9edbb5129f5ae6f512ec95abf7123d3f1de0c04d6b20f0398;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc66d73fc29847594391792da12a178f9a4cde4db201a63d941397370477e92f591d97f2094f34f87edb64fccdbc4cc91904763ab0818e7667d11141f7e7b2f1e978ea57015e5120682b475258a442ab96f908bb4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aeb194115ecd3c897910b4a84408a39e4b83f86cacf4198f6a5316e62702806fda7541f62ea70c30f72f8c39b0c7c420f24d07c7c7708dc001d41d9996f4474f5877221dd78a21a8aee9a96b5dde165520c6a76e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8dd778ba1d9719041a792f95fb84bafbcccc81136267fcb3ec9c339f41d63426f5a93ec6d09cdbf1d565d16f0ef97e4816770058d28179bf688b288d218ecb8a56308d6eb2e20878bbc7472bb1574d3d4428734b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34c533bcc62f2b7eea7bd20770b586ad771276841d829ef4fff801029033ed3f29dfcb552c1f514dca27bb774257447ee05c4bab2feb3c88c53031806f1b000e4a355c6007a0f81bbc74cb64cb0f6bc82508eb125;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8e913e84083e426e735576b685382ee63c36b64490f57fdd2f7869d13efe982e82415f70fcf8f4fcea90d9deaf0023ba9df0cb4ad8f5c549f329d9d134c54f90ad14b44de92f7c25cb13e5bd61a204cd7940c8f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2c63e0a892ecbff685716e6e9c718da8de7fcd17715a6a0ccc1a9825ebb62aefebcee6432c51f31cc398b76276a5a2a65fb22e861249adf39523518d945c36d089c43cec5839e66f04168e37fa5cf171f13c0132;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19af6a9f3039cbd9ea7a56765894828d3043ea976bfc1ba2f6d74ae950f12421f3f43f505ef9fb9ec3b323f3333937a2997eb5249bc3975f78770806cc7f17b4529b6cd96207cc1efb65e30f1d3269137410a3322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2899705febb06e01d5fac0e69e5b72d4ca904ab40c19e9b455d3a82bca0e9e42fbd1c1454e7a58f0db48026f33a84160ed43a34b27d57aae5a78c746e168103e950382a93e1c6bc8a2e57f7c2f72f9ccc845869f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1d68eb307dc4358836d75fc8c0960fb26bb36f7e604238501dac05720c68fa54a45b3c4f53b585dcf61fcfbf85861ce479274430effdd5ba002e7394afabcf1752ffaa85a295e0518b659bcddbc3081f0e9c6c93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he82565ab06d463964d1418769c29f2fe4c1f759474894fcbbb3985cf186bc8d62b2f077416ba18814dafe1e2cbcfcde36e371806198783344c6ea2286d0ac136eb90413d06dcd163a8a229e9ee594e99a90363eb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bb7972b59f287be6e25d0aa2be8097436b19d189012558b927037f2ef66f49135874ddeca484192da64ff8521a9a5f4557816e1cfbf46406900f17df061d265b9cf60fb0d8ecda748721ea65cc901865255f78bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h246293bb068c5aac5c1339ef6848fa265de96a10820e8add97b580d50aa6972d0be25b9c25a5469d22e3cf039a335728c898d2e77eede19d7080405a543ec0725c47c4ed9dc5570198b4b84458421057ba5ecf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba098ba2cf4f5c1da1ebaad6214c60e4024518fdd8ba674b537a3331e2f26d590d352f9d52e582e283f881c8118c25d0de5787ffe705d377297e329b18eb01efe4dda493fede4b5fa37316e2c6d9457bd5c5dd3d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc26ca41c6e12e190cce1fa242a8056c57791ad9e4e31c6b891a4d062d56133c0748b7edfff97ef9369208744a3d533696e9dde2ec605d8db5d3e5e1d3db7327d56bdc6bf443f9beef8ddea0b2458d7a663b8b189;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a9e94f3f7e3c2ec2f71f393367c087be63acf4ce935f241330d0669a7ed8e598041bcde5a94c0520876945c041b6b5232e8a5585f4c9115b50cd65f536128019e6914f54dd230ea47b8185a7eb288a688cf8cd8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e96ee9ab078edc37d33758b60f221faaed54249271812d6fb27408d53ea7123a847ef1eb19814aa97f17654d2ba37d2a4ec5ef9d9ac982f361777e424fb61857c197c3e06d2165e566e17bbb26f84f3df3cc45c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71ce8741a263918529410a6b098ce54a27b8ddc2f95ba6124915ce9a0cf0463c9e732161f93e0a93438091d767276c4cde62b7916f91f7d4849a9f7e5055145c0418db4440a1abce4563fd92d30f577a1c61faf2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7efb1731e81222497a1c39b239b751aa321558764d5f6a8f1790c9fd245478c5aeba68358e3d947229b8161a5d1a9295f9b10d3bfe88c0da9b1beda82a70cf4ef17fc3789abeeac39ba33faab29e92b0da35d18e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7ec681d3b280e07e36067267f5392584135f06b8afd62a23797c70ca3fdf09e999c0b75588394c77da5a6f7eaf405b17bea6bbde8815be0c15ffaf3153013faa0b294823050d743e904ac45935bc78dba812a9c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf48bc073d9b886107419ba0ab56559896ff82f665ff495282d840ebe8e95ff76a16668349805ad99ded8a50f6fa9382f719028bf9ae4d3159f8deea9bc54796fafbcdd9e8bf923259ae00072076899fa15cc58cf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7710df9690cddba5848af52d27d62d468066877afb5492151aa3310e60de0d4b697c02d7d8a84789ebd547c77db86679724a4630212d79e64bb7912bc46b070cd54072e34d98a5432923dd5217e1f95f467f6f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d335ae4ba1afe6cedffb106737514cd71a2b23e2e7fc40c8cbc7315afe18a958550a989558d488c9195935d85180b4c17dd2f4b366f08e2a2265bebe54a439dcb535e43a5f2abf92649e6b63eeb68dfd5b3b52b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha54d07a9bfddf0beb4f9bcc7648d0a1c43c300d8779f1e397e63f406146b4bc3747bce7d3bf480f42d3f044b9fe7b9994db6d354190872d610657dba8160f9cd02f8ae5023c56cb05c91d987c6bf901ae78e129c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14327ae96f5a7172cb1300abcdbacc0c9223720bec59d3427c49465d8424e07e50f4f4c51907c1980b436c29ba5dc26b92d4fd0f36b26594e27befe9908580c71934eb194c71c42120a1ba4dcf2c6fe39ef91f522;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70f897df9af672aef99bc48ce3291a5b8b9918872c67212b22cf9a940486dd747308c9c8351368dbe74d3922ff45e3e315ccb96e9a4c8cfaad63e49771d985bf1b5a98d3cd855e2be1e37263f9e35e865a20f7bfd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2d5857b6895e1538996210497fa3cd220296a8065ab734d43d1f24a038bc475f81d76403d5672e03435b0c3a93b1c992f64971dae83406dcbcecd991bd999589792d74f1dc0f2fcd5e3656b494a293e37e98daf0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45a7ceea6bb52409c98dc68298e11f798091782d1421093410d91f9306b1428103cf004ca0b192e6c04cc1158a8fc8e6cbdf1745b5eab82c704a1d47a1f6c0a32f8def426b46b221520ce73816a190d4cdf6c6815;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h476e1c495b481d23bfba6573bca19e64bd5e24e2f19da0eadfc838c0c90cdf7ba10be92f9576a21fcde21fabb60f3d8505dec1c68faabb7339c7c534971857d9b5d07a5e16056e98f8db696a65a085088322398da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbc295bec8882347ead9d54486645ec5d45b77648773766404f0695b741bf0409e435ce1bf381b6fe9b5bc4d4e42f39172b8d4c57b8f4a80bac3d70f76625b5c45c4f9f20953690eee55bd401d5c568a8bfe76370;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf23f90dabbac06ae45a60d2753dbe0348e5592ff55039e729fca1d43b29a575d8ebaeefe66d53527797aab70d2db1c074b9ab9fd4d80ad57035b66e5b08ef02e9f077a6427aa5640d93eb61936b5f78f9e2a069a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac9e1e73c644af3e0db555211d95f62fe502fdbeafc4d5a460df0bf4365470c3fff73850dcccfbc571559e800c40f0a820d2a66bdbd1e4e79ff139466d0b7ae5f637bc90d00957917152fc61da5aa509dde1e6caf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b4624465f91ac88a6288c4ad81cb56cfc6537ec439efca8e932788533cc0864e18910082541c0660580377dad08dd2427d86af7040002406c465b5fb9419bdd33d7ab0e192679be82bf8c4873d1b4b186c2a818;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c2d43eaceba38ed36e86b7f1feda820ecd7a6e8704795681e185f978d5532e6d5853996807607f822f0c10826ca9fc0da5828a5af014817cdc37c8d5804714f7d03ee1f74b7fb20ba266d3e6217886c60ae48ae1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h437dc02dfe10006526237f1a504f8b905bf5853d9557c3b522cd0392836a093799c3c9382cac5236552d4447893e3f90e380e7ef4e387135f05b802e1c1dfe7955fb30d7965e352bf202a81aacaa352af2f3edf9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e3ed2db24de19f771ce4895dbbdd39a8b4021e14741d978169defc220e502e682564d253b3a24392b56234a6e6c4fecd1709912f95714ddd46702789f42c66ac84aeeb651c95b258c3551eac8d94dc2b44aded22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h666ac2f4c87938ac6949a947be353558cf51f945514c05563c8d15eaebba4edc581a969af42e216839ebe06b559efa2d94e6347dc04cced89d97a4ed13a7d8abfaf35cd93d60ee6132549a99bf3876fbcc80cec8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76fc02d2a5a6248ecf6d1c0ca2a7935e1b74add78ae12adc81e5e053e565d40ce9cb82acae198d0edfe26f33fad477e6bfd2b4ea76348820cc3525ff2b620140f0a91d30de79b5fe722b79c45fcba3a7b5d6bf61d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha844e090874f3bbc1afa4ef7d064b41aeedd0c6f6bcf14229d696f193c6a3feb1f770282f6cff7d82e85f9d6876d8a8ceade4a3ddd4a869cd38117b77b736f72f2592ef6e4e80ea85ec9c4de96dc7d7a105dad79a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h722c9eb6047d33127b940590d277c3c2a247a506d712a42e592bc2221eca69199062bc909a4a3832df83bb45c1bc3e33531e61245a4570c31fcbc4e02ab7d3f33617d5e036c0eb2607333bc14af7effec3883c08f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he82d94852eb6c2af90f3104905b60ad821ce6c2109bbc61a011308c66052083a13c4b4ecb4f8dc13582ecfdc47b4f839e4778717fa261463653fab198dcd7f83cd12e3a31ce36394b88db7cfffffe2c1ad142e33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ed4100b0571a57ed86b723ed25c510559f4135ec5133b31de6244370b65bb45384a96bae1b6c4f5bde8d942011940bdfd6f20791b8a0faaef069d8a88789de4473a134852ed77fe08d7b4790adcfa0beb9db7650;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb23736601f2001fb7959ffa710f3740e85adfdc637b5dfcb75a6725421d4c2c094c6d86c5d8c549b2e5f2570b8041194caa1e327f4b3dfb6cdefac7f13cd849e1f6f53a065ca19ae89abe6e6cab081d4a8c369c40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c8be5861f9d75a994e5fc8ac3fe9bfbbcd61c5d124448b4b9c95621625837ce9d30cf637fd650a3e093a692b1ac002ac72c58a22d2e823394045ebad51b5e1b331edc52e80b7ae382ddd6a83540935c8c3901882;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb5b908d23948e1f14a659ceb8b4f44ddf3aefbe0b36aae055e12a6d2080283de5b3fe0bd4fd3613b014eac2c0eac391ba2b7ddabf295f669874181eb4b902187e2f8791203cd2ea449b499f5f82283fc6174898c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f82be2353a98418854a2378bec6d9ede2814401370e002b1e30e522327b49e8a80f56637f50767b1e9dc6af5a8ac8037e898b411689b7fb034206cf29a45c8c63480eade4e187bbc1899e811076eff68c21b61ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4d8421dc9aec0aea49bea9b9d97d20b40f2ac1f04079046204dbbdf8646c9656997495bbed8502d351382857f7bdcd5e20c9fbee0175ec2372375f0ba6b292b0418084bf37d817d8481ee4f855575e2978736ab4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d6586e895202dc02d540ccd329b1ca6dc8a1ef79a79a91abd14dbbb9f0b5d43e92620805274197fed51204520696a462ece515ae56a7f96a55b060cfcf2827f26a39d83eb5f6f45fb97834786a29152119c81dc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28603f6cb28096a1cfc3eaf328fe00f86300a9e13cfb1136529bbf3e035a0949ede7893cd1c41322b449ccaf51b649da2ad2664f9fd1badaa3527719a03205c2e22fda5d07fb555eeb0845e0e0efcfdebd2ef13ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4079fa6ac19159d4d4ab28ed0f878be7c1a3d60208f29e499fce0791b80203f5ad88b8d33325d9fb6d44c0c74c2d64bbbc645217018f4d7c63ab98b6e932524ffa97c95d8691c4633cfb70795a0cd881e207e2d95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3692346df3e4803b6ffcd96db3fd23fefb7f17ec73cb4a8ed90580a8e1e01980c46efeb9d69818fcbea0793ea2dfa90e14006a640651b2ad54f67710a5ff26d3908ab373995cc09e185087d3f7f74706e1268c127;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30114a3b7507bc8aaf6e94ce7124029f2180ee30513bd97c5f3a77b837bb5f4fb5f9f5a43ce8c17e8aa3aa7de50d22f35695352e25c4f1646fa5f891e24ba396e31101e5f5da48ca6f0a56cb823692f99bcdd8a22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69ca52605cb6bda3ae1d2fc2cdcf4e74b7b14a8463933d82b89413671838a2363b99d060a0169c9c63cdae13be991e04b56581a60f458379643d4e8ff34c0270a7a2a72301bd0b336c5017310741f2dbdbf3e0a00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6da81e6ef3f1828045896bfd6572cb74ace3b4d37e984815f1e06b53b5cce6ab4f3baf36db1857aab9e14fce811b70363c3a48cd04aa5e880eb966756ed83f953a964dbc353cabfb809d2a8954222364cbc3b8f3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80fb8aab72b5e2b3beb5b3146d0ab3ef3ec3f63327bc0d2752e486877bc94002cb3c6c867f7d059b7439d4aa9639001dc9cdb43a9c960e0eaa0f18028c205e5f372e0378fbcd0ef3ace6ea12c5899cb9e252af895;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5e7de609a6ff0f78f06357106a732db510ed709c34c83b1ae00dad030021ffce5104e6af1d40bc8caac230953b8a11e52452a6921d408073d098f67ae607489384bd6b50c50e6a055091d327338c94ba28ea0fbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb57b126280707e1b40863291db2e21a303d62915a1f2d849224d1eb1e587ee71c2851dd9bb9890a3ec4493aad3cd5e9558db359ee47aaa4c0f59f708308b65da95bf7687d727cf297b1681bdd1111b97f6fabb415;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b09ce488ebd0fa938262421781dd4b0cb59f793557e5cde5fdd09324b22973386222e13abd31d399cc145c17b76d0121c6efc6412f35832737dc35a74f6d022bec40c84a2ee57ca1b6da434a5d87cb02ccfbafce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c502f0feebe4fe1ab2541e78eb904858083e4a55df69c68d9d905b3930c3f7e309c18a0c09241d5a7ac604ccb8e33d7dcc9a31a8282aaee3d33dc9730267c2d90b64b9ff4cc552e9cbe0442518371759ddc8c012;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haae60cbbd76c55670b086eb624e1259e8ac0b47517544913eaa234e2b49e69113410c442396af7947452c356bd88e1f257b4eacb1e30d3d643bbfa45f5c87ff06cfa9897ed4e1fd36130c64aee178d10b6ac6b99b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4be5fb64f2fc6766663d712a14bd32e3a04262be47322c9dc4c47d5b1f1dd504c2d88e2ac086651242198f8376c6e0f24143848c1b4998628f48747a3384ec17fbcac5ac56452d42f1cd5b606c0134ee5d36ded2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3fc9b119596f5bda8b58660ba363ed4fcfade5422ceb94c06e1bf5fd7a04953a5a818450653449661644e837eda31d83e5af0fbf8d4a0830307df28eae86eb0113be96bea3035d1f160b0e96844c1ef9cbe765dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc250f02c4f04562adf262fbb7b1576b18582f222c0b026282f421166a94252d7afeb63a0f15b13f4ff090306610abfe57d6fafd29f7bf4aeaefa9c83b5d7b44e6493d9d9ab2c438fb60f6328f5f9a666272c916e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he736aa34ede492999f7b6bcd6e5dbe8d2280d17a1ac4d67ea1b745a51ed08ffcf306aa9d2e81d808b01cb00c8e51e76779609da1b2fda5ee752ca5e04daaaf480ad454052b035531c7d2ec1a37a55aedaedf438c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc999d0a12385e0efc2e37618079bbfc4b3a76b8a7f1b395a7dea3abf487fc08fc4aed1a884d3d1318fc540bbf8c2a40b7364dab815a78fff7265f54a181fe676b8ca112528a4e389cab19a44171a14dc0e7019c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h968e43be500a9293c702e49be6a140ed3ec373ea7404f2933a19ab3c6bb0e2a011b15849c1976a74c667eb7385b0750d7c5991889d409502199f1dff07f884e02363acb648199a176552cdfdfaa038ec4a442936d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3b94b3186a3580ae5ad8307983cbbd1cb0d499e3b23a726ec8667ab379583e511145a0d4300ff7841280b93375cb67d7d45ca2e436b963475f84bc364d93b4d57badf0bde200e032830a1cb1806cd2b4bdca8227;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c3e4b6ea394db239fbafa518927a98e69a1ba0fcc66fbc757f0e89b2727a88e611acda4875c88ca464caeb0bc5a99de4d3c5bc234c066b15f7cf0b719e859391c73abafde8e33774a4df8a4769aec40164bb38bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h414136f4fdde666226d9523fc573ab901d12473764b255379e7bbb1f6d8120c5266e8f7b23d5b4f558832ba9d67a5d47f3d99c430a94ad338904417a97ea7620265721f2d630359982f9cc1529d40a9e08a6500fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0c5e7011193bd3dc22d6ab45a47cee563656de56a896610ca6fd094556ae3d2d21feefa6cc8258d8e0170ddb4d41481622492e0ad50aa2101d6678114527ff20b4ee731da0f9b3eeb705c2e3a69308921a21e542;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ea6d0a92229180eff89938683d9e7a6aec94a7d16473c119cfe106880ab6fe640f976e597a1eb02343e22228139f4394697fd1e5d3eb7be830d57f1d2d77ecb5b643a40c01454b5adbf74cd2ce8df78de51b04d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4452af2140b92b638911fe1a3344b16c1d39c31f603e71077ba79bc82d26c97648711728d926632ab63f9ea893457ee51b24d08cd68b69049537e412d59e4c86a9521e50eb6cfaf569cd09a1c77c64b076e4ba433;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dbc50ba0cd6334459504dfde78a90924a7417dbc5ce66a65499320447756b88968918a7dbee3b098b0adf58baa8d72b44c3010cc16f8d2d5239cb7611c16022655b4d6bd3c87cc201afc8765b5c7260edcf780d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb770a02f8d8d07477bf361f223147f9c26b4d355b8fe99c44f3cf217d7b84c53455f98506cfda78d72a8ba49bdb7ff2c07fbf43ab560f5552f0864c2d3a375088a97039ce1c334980120079effd4d5ccdcfbe336a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h966b8f00882e1e171058f069778ff5960502f1ee93fd2e67a2472b114f766f1675a4cf504c5a677718885e9206e2cc1ca029e0b076330140b6ac3c8180d9c7be06e74cc8aab92e30851f2d7c3e7833054d655cdbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h373cad7a84f65408a50a0f6af871a758bb87faed35efec842864637ad83cb14d3f9c1315b9689fe203e59e83c9698bef1cd36d58260aea6b64627112616b4d1c3c62bac9979006b72c00523bb01aecd9e5708da8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67b4b8c2dbb3be41fd0c0801c9c35d198b1c949e00cfd71f6de2f3bdd4b54e6de1138faf6d0440b61865e32fdc7496922b2ae5f0cf9b0764932a1867a32baaa9a028ab4cf44ad33ba122048b368026e1dc28a0e16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d070e53b701254da619ae08e602883162e578bfb8f75fa2b232fa98829ea36e6e3374e166bf46cf44fbd009622a730c2a6e8e6fba9fa3df2f6850a57c7fac53f276eeeb073da6477fae1a07b5713cf11c2c62e32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf974eef368a8de67c06c6e6b18f13e3cbe8e696e59b770f470c3762452f08e4c9255a957f4d43fb91aadea4ac706559e9d46403d1e8c6a6c1c84bfcdf56bbd7269b738ae2e76cf2702484f1c7ce0339dd6e993a67;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4cf2570c3da3ddcc7d9c04120877f3250b6d85d6d7dd9fc66f2a5b53e51de7c7f66e1faf5045da6ef8f8bad9ddeda1c4b3766478bff6764b31c834adf6d50fb317d8f0bd8b1255e94a9111a1f05999d059cf5401;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe29d8fbfe098ef476c976544e395630a1b0f895707b9f741c61d5d8f8d8b48d6b8c88344bec31b12156c0208a856759cf931e19c6e94fc364259e320ed9f37baca73fccc30a730d93027960835e0ee38caf7980f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64da53f9d214cc2dbc25005bb9431e3df7c9f3e44b395f38a3680f3e8a48ec5a876d77ac0ca795392084e8421c8dabdfbb2baa0b5eac1f1dc11059dc18c1888631444841d21fa0d1476342eddeba7a5041039f838;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe1f49ceea8d661cebe4aafbef5a107ac9fd576c939d6150773317715c596040f403e208207bdc364a4c73d5d22373a3ce7278d784ba49aeb65d425ba480a104386c16341d5beec49c56f70a50bef64281ee9e652;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd13ee3c849b734b20fc6a5e9d11e45e8f9be554118d1cca4d2cec66e0be946ad264e83b6d843482343140c1ad7c155eeb3f666bec480db836f6255ecfd55f1eaefd434ccda771400bf1a26afde0fbb6ca86599d6c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c22add7b9725c9d0fde38488c93dbb3fd0950901ca6dae385d096a3c433c5a645b13fb7319004f74b08803496bb2993ae93fd0e037e3d700dadc2f23d128466d78e9a65055f0ffd7b85cc0bf09cd5ed24f54b930;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cdf5edb59e6ebdf9c308b149204f49481133f5aead99dfde0d3fe5c22f5910790cfe5e2fcc45a8cd112a8f38e0dfe228aaf3853f7b5cc9b5320513187c2206baf7f12458d61110128e0d62a95d4a6647947dd26b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbb1b733368da7fd3c0f4c3294731c077e16a5922aa5d47923bf5bb08c7dfb2e9b6bbc9b013b3d8fe47e0b17315cd5e8721e30f4229f1690e24ae2fc5c31c2cd57be53ff7125c34791abaa49f95d9a6c109c03c9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c432648e1c07c783893362c339dbca1a7c50760345b1cb1ff05c3e545d85c5f318a00437dd2ed76fec5cc3a226f21304c0e4744659cfb22f5240a5017a7c3d66b2673888c6126e8195e4967dc9846ad123a6c8e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h464ac45c28772a8ef2109c3994c6c38641fe1d026011902c90c821fab8817f684c9238bbe32d0ae28ccfd48d81aed47074f7cd469498624b28689b4b53d3a4a523a8b2362ee009cb16329d48e6891dca717e956f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb062b65f5410d7c65a2a9d368cf540c1c66a5e614e5a25c29ac86e641df84e7c515fd91e553e68d23be8be5b1e8dcebca5620475141b88d9d1b19696b1a83e1eeffa6d87c2bde810fcabdd3ad535395eca216ec8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bbd3c2f820eca5026adaaa2dc0229eacf5e3da47656548722c8874f768b03ea5ecb671cb378511d719946d9ff04f04cb1d0c3e186f8a44346ac3f191828fb5960fb53511c89d7e58a9fa636c01819ee02addae69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b2cf13c291ef271165de61ca77a71e004fa0ce9f593f385b7f740fa9749295b371ecb1c082a359f04ca0ca6b68afee580b478e2ed3d0f5f9bf8ab34c1c78654abdfeac54f9b660bf1e2c1c37c14c375425b10fc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec285cbf32172ff09bb30de101d842c957eb6eed943205f42015402cd6443327d668378636f19e7f60061aebe144ad71681eac29a9f8f6c477f0345ae7eb35e16c58dddbd26e4e9d1dcdeca27ab0440ee18acc4aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68c76150f67e8206eb665d461aae8dc9ca6ea6221c83955bcd181c5227062eb0b5d91734fd1e878bb9c6a1e42ec3289e96f611e279d6cfa4ebc63462fe17193369eee3810fa23c5b7686eb7c8d4ccabae58ba12c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d641a04030d43144ffd5731ced190334e9968df5d930ea6a2d12e51b5b7b96d40800e29dd5b64276174b5b80657215960359aa3f1672d46695e5c83ba318225191b8071cee457c0d81dd43a194a90e0a9b9ebc4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e06b2e6c31a6b8b96952d85a2137f4f58e25838302f8f9ff5011d75a877424c3b5e40a861de4be6be0fa895cbe695dc9f2cf05c9aaf11f2da127cdfec42aa5016cdc8850bda72483b3e3d8b82ea8ebe5fd968706;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32c33d1a2c52443e5d39920d72a303d12c0b5b907398d507f1d0d91191b9d8275cba913fa2479c7d8a9e705ac986a641755be32929cccf872e2a38fc059dddfa0ca52131d728c056c157e571a62b134a798acdd74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2cfa761fffb87f2e0159a402b8dd2cd186c69f6a3d5f15f2735d3998b220a59c287868c827653fb5deec2daf900aa7dbd1b985c0a5571a0bbef261962204226e8c2056411e244635117337cbd60b569e5f2e9e17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9a3be6c0c19c2dafae149db58079f5b7daa3c2d3163336a0e1419f681fa7dbfc79c69e88dd8dd9cb1618bf58e95ddbe809cfe1f43e22c7f40fdca2c8aec9e916a0690f390c3e5ebdc6e2022c7f30d5230b5a8428;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e1b2e17c7424f6b96b499a16179da8fdf6e42cde50a4adc607f883f82977be104a86031f2ca6faef9f7eab6c90d3e63d8293cc5d7180f8d8cce8a9e5c3cd2de745b5880139ed3480e3fe50cd809abac5baca7965;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f13c0db0e1805c96f07fd05dbf28f0b3a69096bb2c53ed329560623300d37ed9f5b0729212db5a6e71c16bd511a31653aea623e3c7b2b77fc133931e0239396f47ebbdb0127afc8d9f712ecf6397abfdd051253e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ce62ab1279920f7fe69837afbd7a00168e2adb552f6ebecd14afc6b6ae560f16869db3c55d179a7ffecf36edce919db9f24517e9a43b272a4e31826c2810defe9575ab26d7c21f68c4e9e17a5b6113cd744085bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6582df545d8242bf2c8579536427199e73476b5f1f3da8427c88e4c655771c59447ca9dd0547dd3d4d7847e464a0eadfd6195bf9a8daec3cfc4dc14cc282f00d34588399bbeb5c2c386da37bbc266030ba08625fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ecbc6f4002d50dbec2d5c9960777552afe13e8df613ef6288610479b85d484aebbf5f4b2fbda22084537f9693d73ff718710f3f8cd4c093e40823681a3aa0be0f78368c1957812449f3489f56ab47d1a4e01a66e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb200d68ecd74dfbb08ac28f2d394d43363890a7efb496355b21a7d8008b1b42a2693ee68e9da11c27de8c71d1c849dcedf7e4296ca3d79331f51511fb2ac58840f7ddda1ea9935f2d17ab8a87338a850a5dd32225;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9b0b3dd86f005c2d6b6744c931785f0077deda10ed4478bfd0789b0c74f739672881e18023d8e896af6cf98424d01554cfda9b283d3049b700cdfaa4e00a6a3303856a75ca7fd87c3e981d829ef16e3b7e267236;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b2d7e2a405769d57fa9786df7bb4ed4eac53b78e201f83ed66088b95af88c24434acbd1ccb1166d03737cb8033c95f6fa8ea0f95de69568b91184b73bdd09246bd6dfe0b95a3651eda199b4d79b6af10624417c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ce7a1d2c3c6b84a89cd040fb1a8fafbc874e6dc683157f8fa288e53f6a70c74db5bf2574243bd16f119b82a445429db319e0ac919fd3e5a1bf70aa5800f02c009cfafc5932dbbcbdbdedb0acf90dd097c8880c3f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56809d0ab5019bb4f94e867bdfcea383e428ff1d47beb8fa0b34b15f45a80ba4705151ff61ce06af9c412e5bf21f755afc23a17188af388916a0fbd129904887a333211abcdc00c67f809c8fe5295ff0131e1fe2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9bc659dc6629aad72e6706f662371653aed1857993a63a0a75d97831787c3eb3281f05c31f48a72e2a6def8d43529d905aebd55cd2e9ee573fe13b61c71f19c8f6c93e5360d77931b982126d76f5ef5c60ccb111;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec73ca613167fe7c52f92dcb20006c603547a57759cd7cffdeb8a19595f270a10b126e0db9c0cd2e9e54db16a9206449a455977eca3ed0cddd84a629dc5659b7631116ea4dc61cf301cd7ed8a5b13de02c0712272;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4976c1f19075cdff991529696bc4e1c08392ed496d12901c7ae4d017dd7bf86652829de8b6b9e910ed70f57b3a4fe61fec8ceb4e26ade8de44ae93b912ba8e30ff44c391e713530af1f46e3aa84b66f1ff52b227;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84ac630b99183fa73895f06cf68284dc4384b33cdd38faea6752a7ec740d880de516833c44ec0bc6f88b9227334f7735360e31e90584ca3f4ea1e91a4f4c99bc5b52444375ea00310e8192fd3c45483d682de5acb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h752ff4900c30b93d00e141e5b3db3ef0a7980649aa9b7ae0820722b7e6ef95b9ff489d88134fc3bc4e02d151bb041980dc992630f4b40fab9a33a9ae3bb59adca2d192250a79933d70f38d7bb89d5cca26d240f1d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74267e719897d5c5cfd6aca860a2be7e52a4c940702602cfb66cea6f535ba06244485db5154f24b9f27a4af5a2cfa997877d3164787443b7c9d3775895037e744a6e78f1ae91fa9b7edbc0f3ee940fea91bff3b41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h411e03ad98115a5802e747e55f8183fc5bc8fff188a9bc50d4d38b2a293493c58447600aafe25129d28e9c85899dfefe2e83f4505cbd0a450c6f1c31ed4d5e419aeb3377a94a3abb53aecabc4ce17bf4bbd29a414;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40a88e1aa0e06a609b0b9276c304e88683ebf9eeabeaf6826d916007f8d25c1ead7a66f69ecc44e87049046c16174c23f6564680f1c484cbe6ff09b29863546ba1bb9024fb39aeedf0b9a46d48774264db1c099ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd70e67175428ebb913a051e965703818a4a3671e68d15fc11fa815ad299af0f3236f83fcea764ddbab5274d0659cce840c11aa3d83c1f9d3589c45a42a560b791ffe9897e22d78de7fe924d70c47f8d1187ce8ec9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f83d3cee883f9fe9b7f9ecaa513a7ac7fea5cea636e7776c86ed989a3de61236a2ab8c6d33985f4e678202a1597bf617167a6bb7339574e9899f75dcc90cebcaae00ede11cfa2fc1a628bcadcbffdea97dce9ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74655a02dcaec986516a6c4da18fbfbe5afac08c1a8778f54c637de82a104613cf224e5d41fd265df497d836f59820de9af489be8e7545c63406b8060d0e7050703da4df9cefd877ba8f2ada11236d03de21c5a17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9b565256afbce9002ce83d814335ad93035daf65d344dbb74939aa17a2366f21bd20c1e5a25f3702d675972a12f9e1ffc88d27f47b0122942455cdb883a6037d6feb239081c0db62c2ac16e0691b191170d5c5a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h601cd1603af9ca37d827fd9e05c62af47aa08b5b7deb9ebda900e5c93c19e1d59be939dafb9667ab1b1592c3cc9d6ed693f0479bf25e8e5341e9690ecee506c45044d407661cb67fc4a6d4161ef6b4f45833592e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4fccf2c2c5513d583007b6e940f3b3211145a3fc92f633c0eb6fe1235da6ab4f22c92700b39a587f82dfc82b5fb005b99133ae3ceb9a85caa0a802cf825ef8d944ab10dbe6126f10d247a258f8d2e6cd04aaec02;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9d3394ef188b6282182e94c8d4f233eecb4ec3c062652805594aad7f054feee8649cfc33cfabf21dc3ff1aaf3d046ea2873601111b1b65964078b05087932a8cefeb678da5c03ad4b1ed4f5fd7fde66581e28e56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h627bc96549b3a4944be7a310ad351d1935b794a8207475e83eb53a2a3cdda5f22e4fdbb885f243a12db9587f201fd1fb07d7cae3f9293d0bc25da4173fe676a88ccb03ffa589ff3fa61681bdb220b33db75938b54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h258ac1c317a2d0508faf56da3f5c51a9c53e200360e3e48a3fb7996a112810a7986c19f38f871ed5823909ab62196fb82ce58e72266667f3aed5ae6ead8aa040d2452da6d84d9ca7b721753b178cffb3f87d94647;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h546d515a190403292d95465f13e1561a7f7f92d477d17c185df7e34d17c1d6523927a6914a323aafed16315dde92361b22a376d8624b82ef98e35f077d3f8ded656283f59159a4a11128167020bfd4af09befe37e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaa3dc6bf02542fd584d924355d312e612ecaeefc9e7db677e1ed5c9c2d497f7f1e2444d2527342d672a2635d351f33ef60cca5d5a2baeb074dcda8981f5e922e16e01a8fded233a62ae4a4f219f3bc590bd4da3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h893c42baf5814671bc1891e481f2cad422b7e8486a3f3b5da096d20e56b2b8a8ed359c29d68c7631ca87f7c61d0cd29c5131e9e1610fa1dcd1ae574ccb2e7f2b7d1e27d20476fcc70591b63957899060b465434c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he36069bb6dbdd43b1e029ff3e21640ef14574d13434640789feea3eb8ff484e4db3575362e54ddecfc38134031eee4be0ed2d1f368d8ec82bf7034d50917f5eaef7327b48f9378b4bca90cf8778e306963e03e345;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60f8a945b4fcce6fbcf092d12ebfd12f9fa596d2a6ca4411702f2d612d117e592a4a453e56e630a40b9504b897581878ba63d4678039df4601a80cba4917b4103b9cec67b69b1c203491642241b0cad645126713d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cc139ee9a8b1f84e3d23c91b624347e516e6d072adbed183aa9a8a9b2b7ae29f1a54e3400336c9c142290e5a8416cf882433e965370341ea7116efdff2ce0c69c0a885d377fda3777490aa6b02dbf457447e27cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he882c9678c08f43bbb336fc513a09f80e9f8d4cedf8109466402391e09bb2e92d7d3d178037649d15cdc85d7a951a47f6b1b085056659339cfcf9195c4e63c4ae89bf0e107091c69b3775d3641d47812e00f98727;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h522e1616dfa28c58161c8360484060dcdec0553467e663d2a546a9576d98fc475b227f995881ee14fb791685a8e0a78c8181779e08d66cc4c8f5f56278d7580224f63fbb10a358946304a7cc2dc79c7ff109ef01c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha84a3eb9a1e1e94dcf117053bc0322e2cc39ce431dabf9361edc17c1c1b9c44e9b9fbd081cd6d730ad7ce5b673743aa14cf6a9e5539a127bde8be31786db825b4591880d50c002d4259ffc20b6307fa33da1d4927;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25a0377493853c204cfb132d69c737859e2196ac75d7d6b0e964971096d4ad13c9dcb0dca0a0f1a36cb20c84c799ec461fe317f2987ba1bc0d025e0fabb300c274163d0b82c0105041bcfaa76beeab6c610e7ac4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22edf1a8f288f5d7446dec71e6bfd6130ab1cd59a0db759e00b8cc53e57ca6e6be6419bed9b5e64cfed97126568fec0cfeb55012040720363a58a07dae235e85cc8b4f2fa859e114dfc2aff274393a960d80572d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h225dbab07bd27dbeab1cde727b5684252dd0cad6ed0f7bf3618933647485bfc22107cec7774fc6de653ff2827c8d07d121c80abe022e15bcbc901c45c72fa471da064f45b20c868eda0bf01e6c9dffae8a3b0306c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8523e65b41c83a3bbcf7def675076f6f7b47e9e1fa28d9671de1ff10aa941b79b8c2a6d10aa6e738a7eebd630d4eef1d1bc19b6a9a3258c73f6d3ed4894d5100cf3b9af6e006a642df4cb3ce7c04eef9e467aa983;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84b3ad272e2e0b3e22917dfa528cb38e4c8ce9164d1814b9d5e6e18fac982942672bdebbfceeea2732d1531feccca86592abdb19d7a8b74f734f51e9791773b87dd6f67a2dd1d29e9b2cd6c0da88cce1cb816664;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3769c1e1af636a7b3deef9399825044b71ca2c689aacf17761d4e67770fa232447a3ea3289bea54c193ad8f44548d139638820992d318d1feb47137c4fc278f0e74eb451a9492293ec85e2eedb76aa78eb534ffe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h187cf9a5624c758112747d2d4decb8061475d219e52574c8e341c6fb70426598596826af88ff19d16b577dd13088423b26cc598810c8e20f18f55c58be90a992174843e4a7e50a4a46ead5e817bdd2a6599719740;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cfc3aa7647c4d98ab961b394a25540bcf3008b9df5e7e36090e16fe2e0b819e94a5d42e42a9cede4cc391602200c1673922848df42c20db4cb04d37bc4847ba0c0a8c735024c53633435c9e5662b8e0b4240b939;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha57ecdeb13a97842ae947aa8113d5cc3229ba45edd0abdba31abdd0a36446ba95733bc894c130cf1ad8262f64ff4a084364b3b0648882783eaf70ee0da07f5eb8e9c27126b3cf4b233fc37899fc7748c3b9176541;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cc6f4074c35ed06580eece1cac987cdb4bc37ba0c5fc4ad6f84c49e5a39e9d972ab4808677e9107ac4b05b7748bdcb9706afda31228b992d63f52b4dcd54ef03648176cdb33d23346e7715131297949017866a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb0bfd51d6e2e4a8e2994894ed8b9204d8415d80b21dc37594ffd482163f9b2b1558da12ec0794611992cd2b55c821c4bd534b022a2c0cbe7660484856f07501cb88f395e94127ffef9d1ea978e3b285ae1b6cddb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b7756f64c80c77daf997c091df6dcac1819c3b55e0075fd60cf767e2c0dcc8cbb82a165ff98c28a618bb1ca2076d8011ac08dda91b59d9c3f9c7681b38eefe7c5252bfe3a244d738f7c5a8d0b2e884afae4e839b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had64ee6821276e43b073eb545b99c48541d35f225d09aeb3f0565401d97412b70d1143c2f70fa0e21667e521a9cc3117a5eb838ae0bda6ba9248392a3800393532faefca0e4d362ab08080c43f54462c01341b051;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69ee67ac93491314201a3b378e2a241e6b6af8a11ab01ef87354bd188684a0d110e7440a97e9930c9afd02b4f37511e3e85f9a7411a94663697b193721cdd49f16309db929a19fa44626faaa3adf28ff58903f815;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a9fba0e78bd8c164bfc6439d67ece61edc77cf825c65cd93106a7304904899445cfaeee82e5ee17de456785f1bfee9dfa5c1eb8e340568c43b1f4d73837a59fc5c533d673bfd5f2ef9785ddce093c350e7c0b8c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a73d817d381753c87e2206a5791de8e90e7cb774ba668bed22b1b847d3be07dffb406076758d7904c74445ac206e99850aad4b96eb3d53a0ca935e2d45de4c555556f24b03649000cf4cc9587676f7bb2dd07392;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde7fda94674e7a94641ddd9c22999fa521623f09e0558fde6d994a8b5419f66897f9248e9464922cf0cd30d1e99916b19ee511f7d51a3c59fd5eb8fb7a183ff5eb551d3a38a6ca2f4aa9ceffe9c451a765c60718c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99eff8e3cdd5b5877191c7e6048942bf6d7820c9550f6c47c9cdb675b5800b8d494d3796e0342de4786d012d895b7a566fa5d1eb95c6c0e300ada062fd2ea3bf569827b8f0cb4c7e310990f5719f85666f79f9831;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1764feb97a4114163ee10c64c8667e94396eefcfc4b2e8d1ca10c583e4a920f5aae1d470e8940e14951a7feecfceea538f5fa94709106463d27f1c328f9506f85153ac9e041c2d8ebe65802f5e8d8fd9013136e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15dc139eb0fd777f2bcffcd61b3ecad9c272096c6a69f90c3b9e4eda07eb0c8d3f5d4a4ce09895312bef13fe26c002518cc27e30fc4421341032e05fcb6f222058a677eba7cdb47f7c3bd572bd7444110385f7a5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h529a39aed3d48f1fcb9dca1e9d55e2fdeee7c572008607d46bc8b6de9c06f7ee67475589218f58dff6a2b5ecea45f27b564f0682b105c1c91f408e16b92c8f062492625787ef6e6accba2236e0e25e4c91c59321a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80d5c27027defb0108d59e8c7f7898cab23dcce8b3ad346c24ff63fa9ba21f84f1312936944b745721765007f3a1434934df4355a1fb685922aa3a7e0d8458da4b4231c74e1b66452994ab08348cee5d3b6e0b6c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e0aca713fe6062a62674aa8e691c2d2154d970a3aecd833203f564143d8ef425606c7fb0d9ecb52af468c047dbc8ee375fd8ac15ba79dd28a6ed8fd4fb076c87baa6639fac946105051b48767d12920655fd8a4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1db8a4fcdf9bcd59fa7fd2b4240d0681aa99fea4a92ba7bc5148bd5935923a1bf808cd75cb0fef10ccb2e67a5797f4816f6af50bfc9dd236f087d0c628cbfcf27da415accf5564cebdb21dc7c85072570ec76ede;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26894088f1fca6b29dafac3c564981e8769df65776718f9556687c515650b2b71eec0033dbed4be60b817b8ece2e5c33b90802305dbc8178be80183bd739321f590377ef51283250c7baa7d592434981c8284ad64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b88db87f5dbe1a2d9138a316b3e4ef210a9fface543cc663d6a0587b7477d13e2e1df4772fc99cd780d92d0fa93042b510d9fb77b7754503fec241cb6b1ca79823e86d625b9f2f8c2af28461226c56caf749dba2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4d363422454d6d3e338e95e37857f2b18371f508de1758391228eb56105d22b44d953585340a3bca6c829f6bab8acaf1737e58aabf439f80206e30b427645f485bccef4034cb85c3935becac050265e9635dbfb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88ae019cc0a877d9bfa028fb3c364aa32775b2b3e22784c7f9293b4db581fc9e21fa4d5e433a1215fa87fe1c98316e3ac82b2969ffbcbecdc26e11d6b36e306a08b08d9b0090e590c54e3adfd3bf93fbd10aabfab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5327063ed7bee503afc0ba671a8867b3a322e642bc684f9d7ee6d97ae2c41cb83a2913301dcef873fc4a44c9d4fc1f81083ce09b21d78cc6a6e0eb6a8085b824d82eddf026d8a940c7e03be18bd8810108dbaf17e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed70e7de97397ed94d57c88453d93fd0f05d3a41a2a418f7cc07d8540f31ddd3229f14f4d899fa6b3101dcda4b4bc79fcaaa8d0337bb39c601fd0d26f88ce7575c7a941854205c1fe02d73cb6df3ce7c6eb8f80dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7082bb42b6ad6b88f0d64567a8cafedf1fe89e76415801c8754b410592d071498186de94ee50eba45bd9f17cf9feb0f7c782e8fcaa6f148192e8bc99641f066589381746fb22643f1d85ca50d775e8693df3e423;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92b16274daeb0d16ec8789c6a4ce6321e4acfcd30b8d3b6be807073ee64d33808490330c05aa493aa689ebb37d58fac58b86b3f401b0e7877a2b3f2de1968e2befc2a60b23d4d1583caf1490a1183961d03429596;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63e5161d9e175a8c9b109b298eb5404a577d77ccb807e1988441644cd01001ff5a34ef4b740691e4b5765a774ff316f0f4831b940cb14b922d271ec04d94dd030fce5561d6ffeadc9f9b2f47af495117e19f8714e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd5914b5fe3d9cd678a8419a177c6a4e11869cbfeb78db68d55f07ef4768a0ed8a7dacf677b60017947b9540929bf03fb2ec54f537c8890a690fd14d8488ff4d19a80fd8ae404a6b579c22a7f22e2bab71bb5a15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc44a69972a97367de2398c9bffcdc7b74f3d924610c25ea47bdcf48664c9fcbd295df8870c2f72974544137a8c71e4aa7bb1f2dbe24b7a4e6f8e0c52cb5760d6de9a4de3d359923b009780506b53695bd40577e4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5be68db8d206c2077f9f217d5d7ab162d1ed462ce7690dcbf61d805ab2dac0a708135020c161764bcf47c643f3c546632c83bdf633b599a691be464ffc38d1ac2a609b1476cfb03974b957d1444b798ce034dc323;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h469b1dd450893f76509b63fb8e9ccf9d2443da75b59916720d8305d4353157a386a62b6694d346b473befd3b255bc8faf08cb0c9edb5b0790c01fa4d1d9f07cbdb92a1101c84e5f8e5d06615c571468af74dd31b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha089559ee9d2d54345728f1367b91646558fe3874709dbbf54d796958fbf6bd12dbae3fc57231ce72af4f372d6b609ad1a91659ec623dac7f1e782d00e632a237580a0b261add8bdfb0cd7afe8fc0515d1ac8161a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9214e732fb1b1c6c107d685eae794ed1007cafda0aa56df3d66a32554bfdbfa579488e74b11118299c5e3ff80e25ac68d15d2d9193c1917686bb1b6dbd556b47d89e7509616524f88969edac8ad92b5950e2eec48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb342fca29b41067477f0e543b46e58d83abf4c81883fadf4a31f1d7bba6b5e20b2baa2cdab1c906f0ddb42cd8c9881c2443a0415957583e8097aee993ca505cb1b2a8634fbca310e288d56a96b836e14286d2b2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73acbd16a91a93de48108a1e985c518513cc650cb454b7010549ce3ba719389f8464a08a7caee5b4ab71c4e9ee37ad5d92d9f9e59790faed8a3b1d9e11b1020afe20d9ddbae0d798bfc52af5d14002a5abe51a9c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d83c1790a7062a9ad33d18eef6c5c1aef7e13bba33b90aa645c628e13fef1e18172c9d583abf54a98f5ef55806fc3b3618c27da8de8fda641a3d910b9a0b9f24d6883eabffa3856136084983f6b316a5031dd7fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d15b413319622951ace1f1e03302ee1cbb8d49561f1a53c329116fa4832f62a90b09636cd1f25dfbc25bb97e02f8248db6bb9ee5b3da3a064c07c84280401879c467123c51bf41078ee710c9f84efbea81b049a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bfe91e69abd3f2fb44fce1abb283eda37eb04e674566475360503b6e70f9067796903f525b8b2ee8693a17ef91d5464867b5c02bf2e849254d7f72ee3248e867021f21c7d4d2080163ae6871e54b88f336317080;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c3b60a416570581521d50638f458df415f857ad0d891a8076f33f35f0dac976831d4bc9f4371d4921397754576e99032c76662757327924b6d999dfbd43ca14e14629e0d3ddd004abc64d5d502bb59d648b5cef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2810400628dd0aa3cb3f67ab0c72bb49f688178109528ef7b3704c89c84c888e303da4dbdaee8932f9b125733c80a1786b7a6909097749fe95e0cbf616a0a0fab648974d5ed43fa09ae04ff040151173724a50bf8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeb2c10b17b4a503d37ec9ceae5c20fbed2fc5293152141e9dd7760403155d5daab292bfbdc50bd894c5d7abadc1cda4b317acae1cd3a81d5523d26205a9da9894043246b04c69d69e8dd5f2ce6542387b613873e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb39b54614e15d7c254338b87bbaa51d59b2706b15f27fe380184b1ea34e214a36255eb22af3eb65fe5248769112f9abb05ec9054561e292c7c6428756d7a55b16c59298a42871aecb408df93e0ca51ac4609ad7c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48fedc36e33c2da2dde79ef4890f73e90c302a6fedb5a795a392b83376c9671fe261233952dfb72df1946b6cb7403a4a89f6cb4b107393d2121d0066f0a96abd4d6a0dbc3cb2926313b0c856849c9ca8ecfc00d1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ef7c61d788962c9e6c616dd3381fc8731327b5f15789aeea8e9a6a5b547a20f812c3fefd4b7b7fd3aab0f05fe2590428ca8cbe99a8afeec8c96bf56e9a5544295a7c23dac2263bf0952fe77013197d5b2fb604ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5773bf421e6ed87c7b0d6d0367881f3b661ea5d86d2834351dd4300943ea4267951cefe705d8cd98890a6b5ab7c031f9471eb1c85648c646b81a4549874e965b9a8c4ad8337ad91da1dc2e5f81340a77e94dacc6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b28f656505517d38cf5298428b4cddf5792f2943ffc63e4ba9a831ddbe7e92f751bef4be67ccd4385b919c2fa7a15331ac0138871b30d3be490df5e51ac03a99460d09e93f2353bc833181e35f8e546b0693523c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8677fbf275b965dec5f077490429732a5eed0ab984b33af6ceac1944113781cd36b5f90d93804551f9d56c883e44c970f4613b8ea425f2c2d34cf13a63469d603425ef91b767fd25104c000159e06e4cd931ab057;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7b7c03ddcfe185d43a7ea110d9a688c671572b79e3b929bb6de9676b9977d39d6c026fac3c359498469f255207a88c36be117109d092f8a7f92c8323ec125b11e1196d02553e27cdb6c8760b7342a9f5c5fa9c41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33e66caf59cd694e2ce6706f7aa9e8f78c8e2d9ca4471e87793a4b6fb6a7ce2286eafff0c3eeb935b4ddb609c2963ad081b1e419198e1c812104afa6d500b3868ca1de611799931d26146afc7edb34967985fe04a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h478f1a19c89412570cd252219da03fba201c9ee747c967a3d5b4ec52754c8e3a56a1da368350df2dcea4a0a4d87d69ea1b7abf8777a893d635678f3537cf143c9070f9f5b5abe6eeee8f1bda0f185e4e060eaa1df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha316561bed256de766bcbc407d2b2e29596d1d65b9566a9a78e6196fe830442814fbd30e2317a4cab27693eaaa4cf548304dffffa883d0474e02bc681dbd013fc4c34e48a23980eb83b7d60572c8272d6bab728d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb24056f6eac7c0c53139417874990f57eba59c577bb75a87b7d11b8b70992d1ddb7d191876351197deef0a1a2cb60697eb1fed42c6ca9fcd52ca87b74951c7f6f89822277e3de69d53707e6f2457910d042ecb51f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdbbe3e8c8493b5c0a6c765cebfdf45bd2f75a7f2af4ad7d6e25ecaaa8fe7e201de6d0eb872858ea7dcd3f9f4688dc24dfa55290403c7e02c107d196e01cea3eb25d451fbd5a91c4ac9140ee1fe255f7c2b00dedf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28fdc57802aa1a36995d26acfc7cf5f9476d9e8475205853716467afd75c5bcbe36a5e8c7fc14e8a3c555367e75f81128fee5384b968d1f2311ecdfcef7fffe9f2608772ad7f3a95084c2f99fabd8e89729b1b1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a630b7c1ebad5cbef87af4e21519a1e07808eae91b21ea86ddde09407575b0834434a20b6ebb044bcf59bb12ddcc58ee378e2dea4ff5f9954f7b8d4e7922af5bb708f9968309d2ff23aaf434c9292efa59c6309f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce30c4fd3c05b237ab2bbc960a04769a6083ba70e6d63f79d62076f03a528faf73cf69a5cd186f9dcef366954b9b5235cd9ac6695958584a008e162b16de91c4f6a5d7c63cb7246c61462677f0b05ba45504735bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11fe355524667483488f8387a9abb740c94d701a49dc9da6173d6a1abbc138c598d22e8a3ecfdb3e588ed065d299046b814997dac0fd31d51a859c56468c4d8da0dad7ecd93e5a4661170947b0073b649ded796b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h746c8b08012ea29a680bf63e3ea684f98c56c9deb0930425ab2eb2f7e9de71c669fa82cd96535ef1571c4723b8356a55090782c1a99263d50c2dba5d6c12c6048220135ad02e9d76140259593f627873b055bc4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcda1b6fdb3dc15c0e810cb03d9ddcf2d402763e42fa001531428902ab29c2b904bbf2e9ca66c884e4828ab830ff383c350a1589d332d2c30e5a306620107535791b1799c1228c42861df32cc04942519e6c90be1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f7686a038a2f7fb4ea15858d966db472684b815a4aaf145eb61a6b9766e46091f7c6217a272a412ea051f6df35d462ad50ff6da3ba64e9414c3c8131f8b77d2b9f28d38f76f5bf36250cdb0cdf9f360a33ccf4f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63792f88cd5cc53bf86055a6c0a1d745dd4b75288f3ecf2d3f071cc5e683ae4ac78ad644216953c15462a88862919577dd7b20fe815146afb0b149a1b6b252cbcef8cc97f84e6a3facbfa2d6e181ccfab95865466;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h591d572744e7b72c061617956c1c1511741a54decb96fb24b0b68b3899ca5595be1ef850482b0183804865f47144ea743f52f3d853f57d2b69d00cbb13e6e1f3ad86db5c875a4dc6b2eb028afd0443718075096f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd988d4857ea7bf8e999443b5338790e119e2d438658bc2bc986e8f323d3d328bcd4a0282133a818eff3e62d60e0e61bd6e35ad0372c25652bbd7081645bac920244514e9193d8a43d92c886f672e9bffdbef71a30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e88c8bcf5e04f520ad16b6e0795f9ed0645a1014af812c3d96a4c70b03177b8cad3d45adefa5aa04d5364e395da92a79ad9ef3be961fe75c0b6ae0a91cb9eeb23215d237a24860b1a5fd571293092ecc6e4b1888;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe8524b0c51737d391eef6f17cc8ed66b714695fd57e0aac280f20100a954149027ff53096591a310d74970b729ce662d3cc8cd6249f783ae2f4c27c8da30c7690a2325984f18bced86bb5004852a9698510b0318;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5bd9f9ad521539eb1c155387c4b06b817602573927c23edfc0d576eed3b57334b38e1b31227d4c59dd5566153e97bc5d05e6d2fbd666c4aca9f9f780e51b5c1b8e3b4a15fb61b0454b9bc018dba5e2b19d45e0cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98d697bfac0210da6512a0fb20fb432869f6b62998011ca8326d5352c9a0509d6370abb305737ce26b3903b40d6b82c3c978e3cee7512bd4260e8a0793259d11cd9a8b734fb789bf38498dce4537e6aa47d05b5b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h129a5e4bd910713b64cecca79412a227d201a366cf2e04c8da1b52feb1b3d0210051aa299d3d1bcfb2a5499081b4f924f0e1a1db7c47bacccec9adcd2298b7edf434c93891f726013fb3f1c8d2be72e1da8f1ab14;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3337fd3b7a1c805163770ca7fb5c25f69c86e049213d75b598ff218dbb5f418cf4b3635c00fbef707b3abe59b0087b4372292aa9ac69c583286acfd4a17c2bf6533f4dfb0d76b1ec9dbb50655cd9a5c23b884c90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc08b17bdaec396221e2f0124897ea21187a029632a49672fee54e5315c803a8bd352c54cb6dd08943a45cee6e6f231d452b6dc64a080c6cba5f98495bdc7e89e3a71c4e8e277b69dcf588d36ffb33794b0c6510b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaa3f65e65e589fe8957c2a39d9801dd8f698a06aa450e20acce1d1401a55018b2a53ab1219eba3ecc2be1fd38054c603c71990443080760aa90d1977f08f861e7ded640ec5dabb5a4c751ffc21219750b79da77f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc339448bf1cf9acd5c6995dda77be5fe6ee40b40f61028d92e3099212d9003fb0e2840ee5cb5d1deca7200e92f6e135738db6856961a91e3ca6127b63c92869594ec44e38c7c86f45a4f577e154094fce1fc7e431;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4667970c0151e8d8f40179bb0cfa400af005fd65b226a8b9e928afe15f67d40f3b4d77adfbd371f8d561d58fd377924c77b75808a39e33aa1ba46304fd35f4a9fed77cafef4e4d8dbc098d83ad4599a17fd64002f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e545d0a4befcdd0de8d7fc86d6207781a80e1bb9619e95927e5681c323e4dd5c86169472796e1fbe299b4c94eeb4f1fb03ac5c3c97a32219b3a6ccb2a1fb0496ed4161af4d45847bdc079a8b509a1727c6ef5779;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7323f8da9c18b66e929f256f1c50d3fa431222138ba02d89cd626f8883cd91c90f6add67c52bb874e83b67e9ae1fb278891157d95e7aad54315ea3906f3055bfe472d54028b28bf574f15058bd782411f28bcdcd3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24e78519daf5b7ce1f9549b0ead56a7a093352c6be0004e7dfd5f782ff42e8398f386a34a0fc3aa141fade3d1d7712a90dd86833fd26292be61645f0bc686074c41e37f3eef88508c5b27f26e6e1f3355f3087899;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77cce6edd15c4d2c145848dbda6b1e52aa1405e2719e8c35639563747980caa46568f7ac786081a978e7889b309eaaa937d1be19abf8372a70a85c41d41e3576964bb393af1871c5d0fbb8583114d28d7e78c63f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48b892530d7034636c02d0a43248df58b23d9239225710f3912014bb65275a1fe84215ba9a551a355883643ef32df57779ad78659188e3acecdbac8ae59fff90fa8a003cd8252007370b957d662bc9d4a338be0e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d01800a63abd4b739295af7f77610d40dc9bab5e63e77f8540a22dbd942c636b9e4916ec521bd96edab3adb6329ae35cbb5f7f2916bc252b1b0e54c2a1ceebbc3d98dd2c984a570bdc30048764d8fe8c0d597ed1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd92b086dc0060804bd8521fc0b175bac28bc4b1160be582f8fc3282149f55087fd9c03ff35e31ad29c22a24d53fd7ff7d2a978b751146d583af176f928c56312148239de60e2e6f16175772851d04624397d62a4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h488b115e2f3d03bb3c1b051f53efdfed67296bebaedf00a6da1cb7e00283753fe76026a6428f045ec8dc08f8c3f01ac2b0674d42896bd5e9f3ba5cfee4f0e41ba2f897e70b5e1409dbd020993137928a08061c66d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h425dd204bc0c6abb588cfbb59d41508f89843d6121b1591c36116d1430f339f2d1ffe860c26b6a68f6b57c6d521786d583c558cb56ec702377cad9cf9a4840ec5808a9ae3bb7bac10a792ec31bac5c4e241c0a54c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29ef2bdddcdd73a60208695132f20f46e5779339eb0c8b47675a1b323e179ed858fe2f834032c140cc62791e4c639b9efff34f733641c7ea5eb602ee318a5864050358501f750a4ae7f8972857b65c483937547fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0b20976006e7ac810cff0cce03cf2cb735adbbfd61d83bae2e1a900440ffa31c4de9a10c7c75d4ccd44b36bd0bc2654bf0d58ca111c62004f9107f36fb0af36c7a8fcb46cd8ef446b0f1594ee7bb6d375006865f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbe7dccc2eda47632ec8ace5e67e7047d2c9f2a0c3c0ce9195c8d5a5311b9571787ce76646db707cb6c0b9a61e356fd678f7fa3125f073238390a0398cc2fbe0277fda4439dd0f249457bf76eaadd7c093c270649;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52f6b0feb9863c1af3f1a0d8050bae184c24f34c0649c31e2d640dbb0c8042c71f10ad22f5a49fe52614352a9cbc9427051b8b3d366272cf62d499b96918fa2cd0432274989a986a00ecd751d8af36810948f67dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6583d4538e4fd4481f68e949022b18c4a50a279d4baf79d4b2313c6154a6ab7ccb0f158c4a2896c453bb01a3dfcdf5afa39b00bd56f5b8785c88f178b8da1c56626095dd8a36a9e877afc1b42d4826f3707164a0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h339638200aced43cef6c1e47f480c6548a193137332b4b25f6ad98002ee1f7ab4e917dd032c3710500f2bd291e0aa374815554bd46c31ac25ba5a42597727e812bae2ae33184570f8b0640670b44cd9b266cdd2ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd94de914d6751db4d12d8437731f74a6ec94f4e2072aee43dbda75e3a294c51d271c6b2e900660540b6d5ce320bf2c77eb6e95a21a1cf0e1ecd992740912415c4a7e84d7d3baa63637c2928017b30bdef87352a27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c68187e59e2c5328d9c9a258ac90cfc55fca077129b397b36e5cc5ae7f2ac176fd57360e2c5fb6ea2ffd50c62582bae7394cd40d67bb32f68e2bf232d11984bc53b0d61f9428235d0d2a88bf85181a6af57528a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30664a72f16c9d0db4bd7fb4624ac3ff9f0281e9ef18573bbba4e2e8d16431de167f30410515ea5f4a5da408898d5f36a9cdfd2e08ac6e854bf2c629b904f385c5d57d19476fa109b23e539ae0a14f922937c8a1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54164688c43742ce4900da5cdb0668a02b6dcaf4088ee978d82e75e0392fba47637985ed8edec752cf3fd3ce292db9f3a0c8c6acb381e4ce63bf31cd7c08fa1c097e918c95017ad55421a881b04e072f3d97f26b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab33f33dc9ef754f4aaea4226ab22788ee3521de5fb5049a4b880bc3082c0e44c48289e7e98ce88cd4e438e4bef3e420c60a6da5b4104e299a0a75778156c088853e568cac45f904d1ddd3918c49340c76936e1ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefbb00976da603e545fc8e424bb934e6ff90a05d3b86616cab300780eefb5931667502163dcdf93e3841d4198c2a075eb340ea90396f77f2e1df94b79377a47f78a9ee2d3a41c989b05ae273f105ac11300f33279;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd5e8f9469e2bef6125921df7d80b67166767c9ab84c955accf8622634d20093882a2a2ea79f20fb177bc8b5eaefbe6d50ba5b944a15afec60fbd29d6af4f1a972e11c9fc5217f5aa538decf9311b75fc1a3a8121;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51d45522f34386085b94a6c1494cc612e4d4a19ff313245c8691d06ebaa4d11f432e24df78a0c7f671ac1e941a9f03a9719286c0ba3c61749607b08554acf531c592dc185bdc377ae9a20bc162c542ef45e7463b0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf795d8f2bc2463a199f174581735742e381e51af4aa7036d1fa56d26ab19b514ebd940a4e8a41ba43f8ca8e151c44bd316bb5ba6e3d823c1492c7b2ac9d5d93a9c9cd7b829cf406776de4653200c8904fda285ed5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f3068ce2666b9d84183a3599b878f3992f063fb87ce72ee2a9bc377288c9a4fd642653bb0825f1dc01adb9ef661a0afe6b30a6402561dacb1d168592dda05bcb458e10c306ecbd2b6250c601624479384262870b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7bf92770fc5462a0039b553557eb4bb451894f5127b9f1324fd75ffc64b681ead910b8a99ded3c20599b0019752d4c87057945b0bcd2101055c8d894f75f4a36d8e4c9d372624b4fd186ecf52f57b39c7972e92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59327ae2dc5e19f86e15c60c6997970630cfbc0fd752ec78d40a6b2657e9592b11c6f52bf2239e9e4689fe0123303fe121ee39ae4eca58b7741113c88ca41ad91089e83958f46820aa167c7bd19f917e2d0a23188;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6f37e87cbba4db3c7de3520d0a77be804d45f882ec8a1d4ba6f50fd802edd9eba6de6b55a342c4b71edbc30436e6e90c4211ed5feeea8efb12cddb754c97756945886aff4d6390561098e4adf94517ede339379;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ebc1c2819d32417a862d5228b09b4d791d96cbb050cecd1df5ff203064a06b6995f91a8e469578587c86c4a8ad9a3baf3d5d216d911cbd4f7d61ca831b528186b471e9adb879d17ffa1de4b67054eef37e3635f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc45c29fc79d9a650d8b8799d65256a4fd4d83d5da747eba9c52ee9d51115f64fc75326c78e03e595560cb3580f59f758c90b1fcb0ae87a4f87a10da801888409e2fb51118a6b930f8d6aaac762de253ed0a592f10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a6d71db9207b8ef5a771aa85993df2626663eac5eac098bacfb3ba6821d9073bbdce918b1e9cb6937ede9507d4c34ab53f828c7c7f77fddf055579ad96e5d695e622c8a0ff71d685a6ccb3cbd9d8bbd1d3ec7bbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h599291bc7ce81f8cc8a27c8690bb418b2825b317f9b4db1afd146833ad8a05a320d842f62ef5817f2bafb940c68a9bd1d90e9735df073d6670cfc0810f2ddba69cd3c2da29a2593e367c8d50d3dd6e22b3f876e9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d7a26eb39302ea921b18677d17442fa5f73faea5d2740d2593056b5faa540b1a71826fd4f324b93285bc31a59b72886ac527d2a964c1b9c37e7ee8f5449453521a604781f2a05c488b2d909fe93451fa164041e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7541033974438ae30b25da82ab745889395733b823695a5fe0bc2ad7a52aeec0f13b0518785b44ab421f6338e4b8ccf26f83c000a819ceedc5d437df2f0ec6d59f7ddfe063d2648505450491f994838bb35611ced;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c9320d99a49ed6609511fba8eb248d561865f79a3d16aa60709e0b5b5ec5185dbe503b01f29661c08ee56b8b3580e702ab5392702ccfc66c65b828e2aabdf5ae5c6a4e1f5c413f5e84133e64f35e4024e3ce232e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb46359b136092385afe994307f709ea03aa84a42f329f7dfd62f0f1a51150ed7a4794863964f17578113b9640a7c36e90ac15eb1aa45f8c690556700357395afd63e8b367ef630f64bcd01f129028f98236063b20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94718c1aa6cc2c88f37a81a9dbb2e96b318d08696183f41472d6194a5c39356e7f20bd8f3cf1c3b639f7edcec8d1b0341716acd9bf30356e4789d8639727b5e11b91e75abefc7d81c80340b9f4f9338252b3c5152;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74ba9ba8144356caf029fa06cd029c9a069a9f66116a71311b65288a7843c937cee6ca1ae4308f313b758d4a22fefeac089b51f6e03536bb997811e932ce35c9ffe096195d746891ef12e8d051f70e9723f4e9ad7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3029c42007c4b3dca9fa2937ea3a0fb988fdf9691c667f4dc4e69de0f572767b5f5440b62d2230a4d3e64f026d622b1bf92283f42c08d8e70741d056f5ea6be977d9ff66880ac66b112cf39e408b203b82442822;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa227b9eab3c4d6a593fdc9ec8d59e094d1a5be10ee6b3457d9fe232b56188435c594dbae77d143dbdf53c06cc285af6957e4201977307d98352e4ec5c2148a3ed7fe19e0d8b060b5f3c160d9446ae5e128195ea3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ca6ee9e25db5ed1a0ddab006436a5afa5d8c9fb614aeebaffdd8b577009d84cbfe178918ed0d000af98bec175b77907a00116b934c320356e9973d2805a4423c451cc894a087bc569573fa45e78cae0c92d5a9c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c16bde2bebb0a829aeaff437b4be96d2460e6f8a045d60b0e75f9a86f1e063a8a57ce93a63b9330b78010191859113df20863296a00b59491003a2572a0c6ce79e3668be28472e8e883925d75aa29470032142bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5eb77a667bea8ab5e7745c517a81553b2cc7a25588baa7d1c8ddb9a8ef6a0ae6b7ce37d7bc51939e06fdbf09bdc7d340bd3bc91c50b7b49b08e1be87c8f01eb9be6f3cf9d81438db44e6cd0e848e8c1b242f6b91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h973d40b9681764876f97b81e890cf183b2d0b09e78a9b4fa5ca5d12b190d6b31f97ed818c7cd7c506e6457821dfa7400dd890495caed2c21214e7259ae661e36cba0efc82a62be412a6abd06a64d49f10d4523bc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h478740945c5714254304367834d933ce4ee5488eecdc3eb6b15192885f65084670dd0f19fde903a07b322a857f1e733f869099ac5300b4d902f2aa8920f7b8fc7279fd5c44cafb760a402b76d88a5ddb390a00d8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h876a2a245fe026b8e849de55679db5c2244114ec49bc37d4112606c4935e5db49bfbc1a556ee449343093e9fce07753807be92ebc9278ada6cc6a87af1ffa081d1a570df87bdb45b5e7d99fb38c95af8d47c90706;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb470fa53cbaf725fa04b79671f165d982019c072266ae1d075b408c22a04abff2ed4db1d182919b481988d1ae3f7405a8c79fb7fbd501dcbcf0d58618d53d43a3fca220e0980972abfeb06e33acb6c1cb44c33c89;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6d4761067be6626811485ca3ab8eb81674820d7456a0e4f006fea99e94e0be924c17c01825cd7274246ac7e1b91eb2099458c1be47802382f20d33040386952a6fb681a1d902c1742bfe7d947e697e3503827b16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0d68a556241af48c3c8cf08d5e1effaedebe11f6fa0ae63ed03a76ca8326f524e997f87e0c08cbdb17d2cc23147d14b610341a51d140b65cbbce9f542a9c0fd0149efde47d67def2544c02cd9da0de205a61227f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9b2014c4a5709ca3e37a7716d90d06c2c833694becd1c8cd18f6c49ab932eb19dffa8a8d6d541115eecb134f59fb284959ecbda957e97584979f7cbb8637efc58ff1e710e5bc7b0e90757e1b234f26655f32dc5f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f1f0e9d4aa11cded64fe70e81011f3080fa564d25c05a466dd52b8fc8eac9af7c02d69030d9fd25355b9fd7138256a7463c434def70be4b8f95ea1eb664dbd79862a7ff3019b6fa173a23268db9c527aaf358c22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h304beb5aa360b1fc05abcd9066523e4e90a758bfb8a53ac6b2606c4efbff45a6b7fbda0c4f0afdebe8122b8756ce3b3c46973936a57f76d0c82ef54f844a5f5b3c75a37e85a8d9f3143483c4be05c6df2501b237a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7b5f25e8b2e33641991476a885eb7ede4ebcff6bc2cdea9040e382d96edf22ebd8bee849f585be0d0ce7c3a878333a37a6b69ff6363701c4a5c7afd480a9790626146f5211f70e2734e7272eff97b1ae9c0ccecc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93d7c3eab71241f32c04b7d8ddaaff7e340c110bf1ddce5429038b18281d02ddfeec1c2bcdd7dff4d12a1ddde0e62de627181b3e76cd6e1fc92918b2d2e422ad9c00a455fdaa9ac6ba5fcd6da9d739cd072129640;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43157427521e5e12338db021e43a5e06ba0632fbab7d23b31afc8d7b2247c04b3f9bd20f7200e734750ca0a03cbaeda1dac55ccc353059a75489bd685501a72db7f5505f73ff11a76d35d73b4f51969dcfbe7959;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b9005fcd83a9b9291cad36c0605630f0a5317b59ba44dfea0761e57fafa263d1c2c7098a4b1fd953d31c9cc9b97812d9287d07dfb727d3f7017c455f4d5194969fa866fbe8502cd9d2ef6808fcb61732fbfa263d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84b002ceed6b2d4ec3f520ed0e8e184be8e96d90b79a559095547e9d82ac73305e07686c13851d46a706000471e74a8f1e5b2cc09e44c9d8c487fd7caf48990cd43dcab6ba1f9b1c010da2ab801ce367ce37425bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85d2f5fca1efd5333c7c47446885e72ad2f058dc457838c5009aa20ed1f0ecbe2587f39dc9ea131182689376e7bf6f6be4c424831d6b011c09300a49955fcdf0f22483ac49d6947414f82425105ee0290544bd981;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf294975868980e737c2309eb2952921cbcef8730fd8046db32eba6ebca479b37dd0fa18dc1130366d2e1a7c230e8358fe136b9a78143251042db254d070fb4874038f1f1ed45d99e772bf5aae8a6ccd3ae1c05aa2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63c2db210375f41c818edeb816c32e3c037794c79df016606716bff2c7e0f517332551a862c49f484f2c1e9d6f98ac8e0b2171c97e2836caf2a76bcc003ea4af30dc0e8df9002d7df674dd302008c8436b04a0595;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77060c953964fc9bc34b432df87ebc957186ab34e48ca66580475f763fa6daa546e145467be0ec73a283e9c331ad552a4c54d026b559b05b9b28b8fbe98dafb37bb5cfbfd93cca9c91cf15021ea77ecd73aa49e89;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h264fcd38a6adad19bb4c1d96ba621516f30aadee6fc3e1855bed28869c97fe14f14cb6c745ea85c8b0f23c7856dbda593d99513e14808102938d79e7c916f0e291e657cde6c22cf3d5ae68ecb6f8c062fb2bfdf20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ef5e44dafae123e536224b6c7ef895b1fbd404c6079c1dcf283e2e909940bc4ac8a9918fb32405b756fdc73b29e99fe1b9d5e8e3be4a59e292410a9add462daf16995281a1ac515c0d54213b1e83d159721fa29f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31d06413aa40cad98c860d05746bdb28d25167e576afeb5102e62425f60e283d09116bc1a4c2825f113a64b7794053edb870304acd633c3007f4c7fca149795f3d7ba59c13fcb41a38f4870c39b9c74bed5ec5aef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b2a9152749591876dae4779f3e3c545f06256965077f3539a6329c133e46cfe89d15bdaf82f95df33bc1a0e2ca606a60acd286762ed19f8e5c86c51bc34ead488f868d4d07693b7a3c021160ecfa35e381ce7dfb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69ec48e225a990acc206b9ecdb5489558f7b18b81700144acdabdeb59727c623ca2db2bc3036460c01f69093e6c92302a9afc85edaf0f938d883113b8ec62a06636257282a031668a06b93077a227716c29dc725f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcbd74ae26ea239be003d199d5a0dd323632093b83c7d0fa446f0f7ae4fc301f0ac79edca34b2b0f765b28183fea3fb8e36cdd9561f7a1bce45f6f275b0decc8ed61a43914d7fcedde07894e805bd5de201657d33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca075c8bb087b7bdcea25d4cdff1dcaa1fb3c95ee261fe3640f1e94a33066580a95e3a5382a67c8365edebede5ab5f0b0adf1cf5da5718c29e19742b925cf77cac2dc3ce24e44c6244d34f3efbb66227323f11d7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a941330dc3198657265c9e2e80f08aad211ea5b6384080fb5e92f2ff85064a539bb767886d5222a60e26c1ed287d04b2747164408c5c0bedbd2d96be56f5df87d3145751637a99edd593007e96a3142a17f89aad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e9320dd236a07fd747f7641edea027a3bdee61561e8f1daf5630aa86a257b938042fdc9ffd67ad065a5baf25143b714e745bb6f55b00a605e29db072131a2c479f26e0dea692c46720a05030c8c794809fc29edc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha25c2899ee2d417b47403ec74c40cdac36d0790489d9fc5ec8b9a0f2166f01c4caf0f2fc09b089da8b7d439010b1ada6aa2f2b90adcedbe50d5ea7a62926ae76d1c35c2b3f2ac5d2913a5ce321889fd84c09a74ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85a2b33c89562a31c8aa1694bc9515e56ebfba5fb0945eb94200d2bcfc10e2893723daf8d6ae2a0ce208a1ddc90ee75b9c22b8d74280377da47d1efeac2f9b9189078adb327057df9ac22f56ff0ecf8fab82cd8ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h284aaccf31c8651dda1ee4465e9e8e3e5c73067486a33d12c8b8da5012f794d39741d0a66eafa0a9b9cb6aa36680524cfb3f9c119c1bd55c36f213624bffb47ea584e2bc44a543f7e103baa424d3289b6601f3634;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h673284c56e1afee75967eb5799717499d8b8aacee5890cf4a4c506b30e1f6628e508c5420aa52f92bab272824df4924d12ab0684382d13b35d1c166a594cdd3610e477dd04d00a734cffb72d97c6557a494d487ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc78fe7c50ec5fc228ff5cd09184efacaf295dc774e9f33b2e81234afc861d056bfc3d2ebeb1c913778f17031924fdd737fd683ff8dd13e84ab7e3284e109d3c12284123069c0655116143796c7972a10ea2e6d82c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8451b841f770343e147b6adc28bf52415c921ec6bf307c6489ebafdd786faa774f6950d95f3aecac2bf172cbf0af4226ce5acc7e449573b346592858fa2ab6ab977287cdc4bf7c01753caf67293e0c309dd1660c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1483d6379dbe5dd62654c3d3ae4aedf0b8c189c86b57410daa94657136f9b1699b72d55e03816ec975f27bce1e4435bf00a0db8827fe305df3b11f38b04b6c7571e00d26f5d44f48de2a54f169d69a579d70e5a6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a1c77ff2145cbdde5c99e40493a2be7c2f704a2469da3657ada8c6a06ce894d66845e890f07ddd1afa2568ec7203b6283845f3211faa1f8a3a78d2986186e5b1851734458589469eaf2eaed1c34e5168d2187a70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fc30d7817cd642e7085048533635614687e9771ccdb2b19ad6f7414fba6619b845b21d03ae52fd33610346c97f88af99a81e8d65d458a2278ff71cef79a3ef3fbbb778c49804f69da988ef47314b8aa9b7dcd6ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd301e05ccb455ef85e8b14b6b1bb8e73977d944dee73c066b4455c7acc738e25034cef8724b9abab4c0b60fd0b1f4af46383ea8b0128f7395d7a8468b986dd6474acdd5add0ae87f7c54ce6540d2312e50a400567;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he27d568c9edf4206ca471a27ee93bda5a3ccbc2e181807974f015cc13f20c0e48e60f631c9f48d13dce05ae4cea5e4f302ba733d46ba3607b9ef070096ade547fd3d712c232e931298f99ff7ab5c33fa23b915003;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c295abd40f13d6596ea383df06ec1cbe37246c674e56f71abebdfbfa073a8c37bbe7ac55e10947945c9f3348fa13cd000a62a7e9de75ac133a351d364858cff8a45555224c359cf550746809298f574c0d7de6bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c80b8237802b51740257d637b1c729a5cc6b83faad53994c9ac5be1d4882a78b7ed7894f2e2bb12284e974bf2c3f775f70bc73fb2c316dbf025e6b267ade199da5df2e78136805adc535c0d5c08ec6438790ac03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c22b3321b0708eb721d031aeca63d729896259b60e7d30a71fa5f183cc2fea54d7570bc49013342dfdfd66f17007779c6e4bbe430e87431aceb1ee5449fa343df75e1114a25225b8aafe1d6fe223b9c1faeeea11;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf7f67c95764063659e8db5902776a4c4cb6994d4c20d00fa854b810bf93e606eb2d0476729532c5c0626c95cd8201ceae864621ab027af6ab6576fb447e5b33402d7139380256636092f1e10163287bb93674232;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1dd46e586aef521272e7f497c868ce65dfd9c086a78e18c61814d2dd93f00f2ce303b7efbec4c453aca1ef901924c4fe3af72f25902af2d85b9b5aeb22c4a9c442c7651c97acd86ea82dee7bdf830a2f60d68a2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec7566ce4898e5e4530a4cb94a7a09668892ff90bc700a7ce9dcb537e1f5bbf95b8b4d1ef5d1f7a5b30a97f8cffb0f01f4d8c704c0540e46e1f5d65e20f0a414fd87fac7eceb491e0be4fc1fc8f39085bd7fe7951;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c4c32909a5783fa9ee184d0a545e613b868e0d66c0a2ebf96eb48e75f7699ab9fa1c0e655ab04ac669741f8f3b0a285b4bd16c9453ef7b8eed3b304aa835c25bfe51260fd6b59fed6381c75bc01bc5ebb0c153f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc69d613483fe7fa74534c2b44b3031c53e8d1ff72a09f1b0a9be74fd675590cd583037b764ef080048f084867362f41a7be32758fe828160f191109b0c27b2e9564032bbbe91229d017e41278eac0b7cef8cc34ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h625bfc34c7413eeaa92e8720f541c19df74029b331d541edb8637615598fa35704b18482a474720191807f212dd95c23c50a7917d4007cdb692ffeb42b4b3a29a750127ddb0095e9c9c22fe6fa1225a4bd37b1e30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha65642734d352daeda226a18988e65086e4bda4f84d1560ba5f248548d6066472dd3057cf991cf8dbc99101fd85514e238852dda165d23d8e4d149ed2d052c86c68d7977654c8bdf9cbdffd0d3740d3907e5c8b30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bfddd25137a3d511a8c48c2dae3b099ef79f123a815210839f2ee6e415ee56c25c2039af8c21488ccbf3cc5f0c42f47051ff8dd54bdc10871f80850cc3fafc669fec2fd9dbd29eca2c3c273f20ed259bda55b060;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c8350e178bca7fe6729a01bc934834a39d2a640acab997a0f24612f002a21ad6ee55d06c27c61830798f01bcd1e425e795ac32835fc25dd52660de7a70d091f8664533dea915488741b2acc225fd5540e891a62b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaecb0ae3d436deefc77943b1b20de44721bb75e1e3ea9f5ffab9e12dc399ebe89067bcd5543c9d2cbb5da19bbdbf0560cfca754dad6106a3201c635b962a289e747228c0496ec42f56dcaff468e181236fedab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc759c078c4177377765259f7f7a91a0582ddc5874aaeb5e3086b790dad12d4865e4e974a1453f9509c61b99111de11551773fd225b95f6743aca235ae6b20faa3b1d197fc5f73c011d1b29108ade716f93c8f8988;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9053efdd2b250043d854f295d79b2b791054cf2be855e51a37f989488d2800d537286ffad6c7a6bc357861faa31a0e05117f13ddf0fc4513903eca22f99947cd6bc134d958ed6ccf84fe67833cc5f555369b59e6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7d9a395cbfe2dc3782ebf14a45705cc61672f0ed5300324ab5e3d5b5986695f43fc91ec57d396c24991b925ba07c015d17d5c300bd7653eb0605a06173a7a241bf35aa42e2cb7fd7803d07d7bf41deabcfd33190;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8339512a3610a937146f8d95195e537a73ded2ca1c03237c505157cf1d2b69617a21b155e2b42752507110f76fb9ac779ce7bbae88983890667be37620a2e8ff125fccc8f1d6aaff2125b85aa2b6631334e022d8d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5d8ba1e77ffc1b5eaae8265b718fc4c44dc901174d3b5d01d4bda25b69cc3a8436b103539f39ef17395f52bb375ca117bcb0d1c8c19bc3b6aca461845b942f2b2af268018c79f22a0afa30cf1027cdd05f119952;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h505d1afc055cbc55160525b3a8ded6fa50e3cf284ac9a7225d9020626b4d8821db4f9b2f259a92dbac2ff03c765c8d9cf9ea3698fda61ae24ff877e6780d3df08f9729069d961f371c17106ef4507242c306f2439;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12a88de2ddd03e3e81116a64ff1cb557d5b13fe884e5b7734da489b358724a5c5a058662937a1cc50d86694a21f44d0d9b45d88cbb1b70d434d915ed385e29d0555a7879c34605c453fcce3aa8278eadffc1f0f9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2583285cebcc715f20e6b7286c9418154090aad4a6dab83f4e793f5447c138b4adea60e1f49871a7a858fa1f5158e6f46798b1f146b31fdc6954900bc303018c5f0f7a74e291c3f9ca8aa933c52e78369218ec7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a337330d75bf26afea4707a7346a5a25a5fb8757693008c8ec6307d716f47693c832c9949d084c3e7f0af13364d74ad7e7a375b357910b7299f8731b00ddd2e87426ca8ff87875c66509c9bd738f2873042ba48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85e29576fb6035ebcd847d780474cb46c15d9ea75a039ee97b7f4c25620f176b0db6abc1ad7d4e169fb1638e3e270f7e4b5354955c5f195412a4057b832a9cd2bea381465858d146fd3b0c0211609c7080ae329c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ea9ea66f303e08fccaae52be4bc21acce9c0590d335c84e1bfff5bee05615e7a411d7655133f24e9f5bc23903804002c6a1aba4af08b774b45f467e5b91a26fbac8ad06d3e95909544bbd03e54c677dba426f105;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbc5e55a3b0103ee14955ee20a77d8bd627f4d6102ac43f0802541ca1040e8c455456800818ba165f4caf380044fd41c894af29be446fcd4e53f12407f4f5b5c2452c3f7f33112317aa35e60fda1bd39ddcec7663;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17713bbea5839117038a48c6fda56510e05f62ee9eb3508948ada99ab969beaa4e6e1c48ee3efce5258c3e9aff4deaecfe1b6ef9d85bc1f3a34fd3854869855c7b9cdd7551a96500757a9f65f2277f6405c922268;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49ca45e71a59992a39df4e4393c09f3b1b77bf1296f80fa25c6f11712476d751fe3c3d4917b3c0647c6cead6a9473a4ee2a38e5653efd096825420c0ed286754b1835cfc82b15b7abd74099f0f9a19e89c214a81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef13aec5b1e1e63bf927055ae361c85828b7cf957d2ddaf24eb7e7b6b21b7747b2da554177c99811da186e84f338f9fdeba90af361e6c749a64095173aa70cc010125421440cf8a1cae844ae3171911e5af50c970;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd65994bf8b737a12d87700876149f75b94655f2aa938fb88373891ac8593e7e0cd6be4f4a84596c4cdb4f7af20e414f4d267a43ddc28e8a9b2b0d720c2f87fcb48f980f268466386a611685d55d2728c74358aada;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf7b908164ce925b6fc67cf75cb53b5b6b62501877ca951d1aa09b68a5f4b6b99e3bf78268cbd3e0d40db779a9b2eac5eb9f6d8ec68b4858a4a1d6af36c49efe4d06973a39f5e9e49749ded18613c388138d4e973;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha63f72f4e5106139f3950ac9dd3508a61391f5086dfb3b4b7316834337496b733966dd258487207030ae01fd668c1af6bbdd65f65a64ae1e1ccb08475f27951f37684d4bcf682c0226245f5b5172fc8441bc4d2f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5384b880c36a29f8c7d5a01c929b533522c066e3ab0f5ffe2862d5170a16236282fcb5bf974a22703b9642ad1bf8092a289b921b98e4415fe23339f99b9fa5b22281f13df75fc93a658b865a405d7592b93b40f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb01bf82301e4e16d9dfbb935c702b40de112ff0c13ee8cb2a173e8be04bb87e2b8151659f9009a7d14bfe81587155c31565aa105b87a50774bc400fe947761bca9a579df48e2e4c89b69f95783781661a2a8b07d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55f7ad8ba4cf60e1a97ea961979d5c6eb42e8065154c4760efee9399b1384d13c5f16846e98cf66f8dc4a07de8913578955662333a6ab398a1663676b3605d3aeeedcfc6ee0074da363fe3095754c9fc5c378e802;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdddc15c9a147b67e0e998cd12683844c5236e5bd5358d9915dea839cf1363a30359dc2243f7d7a0dfb33817677b082f047989d02a1088abc1bb8f18a6250d18a5acfc889aafb401a4f9e0c8816f5f5e9c470a02cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21d92c9e7bf58b13200b08b2d3275011b3ceaad5ed6b9a2f2f391e7e2fcfae41fc270805e0e3bf19d07b9522ca87ee69005d850cce10fb86f6d9ca600d0a3dc95ace68bda8745b60d995c1d8e78eafe3516a5c43f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h753881f658acb767cc57eaf5a20037e1441c200e17bb7d6bd14d6ccb76e439dda3e71e94aa817efa880377efb513a3bb9759d0643d92ea5496ec677e5cbaf9c1d9f42b02c2c663c9027598b7531aa58818a534474;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c5169ff862f6f8bd90142d0d771b4d02c327e958a0d290e390013664c6f92511c01beb6761cfe5ca51cd5bd166a1680d74daad48fdd6318403923b797408a408e1fe7a81c82c8fa6b58b792bb4761a6968e4222a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf3bd5ef6c7130cfcc99d762661bf9e9e663461ece85f46b2c4af42368a509cbe72baf49f4a6c0df74dc65a7df12dc2d66794aa97a6eeb580d23b4eb6881523099f3e9f3b4b3894afb06118316b556ab1913583e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bf46b908bd4cf2c46ef3e03d078da4d6c8f73c4574e0f33ae75afaa35fe4156037866368d2e0a43e96573b1c8b6bdf951bc5da0cc8233aa377905fff0f8e1e35f091d8326cacc1b4ef61739fcbbd50f370cb3cde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cb7473e87fff16b1a69438f0bfcc8e972a552d1f2b755d1605f4b5d24762891534f6b65bbb421cc2df5d601cb404ea109ae75b5223fee9daaaf576de486596bf0fc26910e8499b076e5a94c84f42c2d9f14b57d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9451074f5874a3a28c9894e797cbdd9d37a944f9119e69e720287a161ef845c509230ecd53ef2634a3fcd33dae8b00a1405290705ffff8d15b0949a1bacb5d0ebdc1c0c1f723a731cdbe0b6c727b943e2d6567abd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34b3dc367978c8236f02183277c0479ca572d39dce4a3ee7713fd702717ec3d3ea38cad2b37722528f537b02a35fad3af4194082071226ae0bad5e98aca28c5b1a7ff378f874981c6892e3a09886867d4dd288ce4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14a144bb04ce9cd97cc6bb0c40f9bc7b9ece45335e0354eb136add65af816086d29efd056d50eeb80364b3b0bf7d5752497cdb341b34ffb55bf2b2530ca3ad0c0a2995ffa00862275ddd2decdfb1261fb76f3bda1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9196e28d958f101ac91a723ce010bdf06f2ecab2015d3e2652e4b0602938fba6eb658b7f31fdc5028e59360897314ca2fc6315d4b802df4feaab10081002185990a3aa888133345a0470549bbd24f42506cc824b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cf081ec2722fce8c0c3645db7122ba5a4d33447719b766355f340db18426db637e7b305c4fe3b7f1573f5f724e38a8abfbec1e6ed8956a0a06a1271d2ae8017bd13d6ba4fcfc06d9db040f34d62db21fce7ba902;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60249b0e057b07469d913f59aa5d93256603a81589d92183d98737410c8d29ba3ed53fba8214931156b7d62f759a1d415ac5437e400e52ed727d127eb3195dd1ad11583146aab9d45b7eced2c7695fda3842e13de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf5808c78afb6ee288140d1e7b2ffe178270ec8e2f0559dfe889cd03c593e5be38cd4453398563c7e9bdfbbea0b210d78f4473c7034ca4298b6b703f2248fdf906dc2a7dd6f13e0d257ac128bd58c7e092e7f7a4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6342a4028eb8eed4ec2672bd0b1d3c2b60381831e9b85d209766b6394c40ac6c4bc6327a57be80ad2174887f55eee98e587ec5fec699734d218de8d038e11126c5e10b0f2c02b140ef5cdb2a20176cd5ad9ca00ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1dc90eb472a4c791bd0e946c59d7098a50e5b74e17214586a69a7e305e7165960053248d177c9066a7f20cb0bdefca7700e13bccb7d701cf04f7604be29e3a13e8b94a01340d90a2765916827b9c406bb89e6632;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc83e4d45be4b1656689aecf5025eb36f306218d6ec5f8b054f858c528fa257f8508d72acab88918d88fdb188fb9909d27c74cb873d06e00a558d8bbeb4cf37ca3a17a804f6750134499d19b9e2c7dca6a9b0fbdb8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19cd65de8e32279ae7b01d52451ad7dea3a0e4221b12559c0e6a3cdbcf820f32c71ad7359383a399eee14005332e3b66af36b20fe474f763ebe9e1e836f4c1ee0e9d773842e5f7070609ff2373ae1da8ae0ac7b3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd470c99ab706c4e8f97131c39dcbff342fdd2fa0d9b6072355e24056335d09481de8e640f50154557af8a995f67718b0c108856359f20790ff124ebe8a9cd1daca5ea44914a881fc5b90c1fbb8e1834f3ca24376;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8d770cac1954005315911cb98b54959ec703df2a3986e24cd09eadd870e902df4e9470821f3467862ac1f2e8f4962066657974c8b16f6575d95b86652f30b7866aa3534844a5ecf4b9be367757e99b80c04d752a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3b6f83744e0618fcb9dd144bb5aa9843ea2d000bbb2df6617695cc231980bb6eac5c8f292d3f1a19b61b61da903a76b10a960aa06cee4f1a6cd3e6570316bcc3af40991b62256676487be6e02a6bf8c6abdee889;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24e778e74e432bd47b3775f75175e17ced0e861a466b2ebf33ca6195fa4a4d7f259bfbbb70bff49d924854ff193c0633ae84fc57757abcd486057a81d467674bf46eeb117ed661ba5fdaa38f49677b7c1280f7376;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef4f3bd7d18c751c595e2d11439d250f79f27511a46612cedf6d8a9ed33576d3a1d5b93e7aac597aee59b55d210256f0587b3a15b4bfc6ec76d6991a4d8380d73c347de1f8da36f5fa49b8e721afb5ca3035fd6bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b74302fc2acb2a18ec8666580ebb088eae561c18b868f3db0f89360aa3580a18c5f5d81a4665b98fb814066e7d9b065d7f9d49affbc082e659423a08148454d00e083a9890f9502ec939a1a755d2ad852487ee82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a0db16a29fe15f6b4c88fb6a75b8450a86cc86ec3416e30be949ef194af7e9ffb8e2cdc45aed326fb3ab7533a55cf962d72d85f113bef0000f295a2b5058004c6ac4b3dfc136e3c3e4a048caa74695c17789a19b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5125db4bb3d154cd60daeee0e2273fbb395590cc1e4470c76a348baee95dc564ba1f1566e643138ff83335e703eb132ba153ea4743b11f8eda57119be7960280ec8ae25a0e674c28a9218c0199e00a8ef2ea13f27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedc27cae6f07480da9335c5034a9b1e337614ea67a6fd31027bc54c10253c00baf09239a1e0b7762faea80f7c2fdd34f5dd39e74d88cbae097114c18b0666d9abf4cd30e4a9bea6044bd0847849e49b328a06b10d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3059194003fb6d88f04fe807775da3fb76683a9fd69b7390f68fab242b5fce2bd9f6b3440c50948c17aebc0e4571e9e7c4de3826244c75e4a11e98c39c7ccb79ce8179b5c9a3e5a6f9ea87d34acb183b91198deab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he744a69070dfc6fe839d01a5e41dc701acd2eae810989bbca752396f645f4dbfc478d0d0d042a97683abb93be5e58a5e4313ea24cf6e544e5fd3c284e1f2f12e9c039b3a3e0523e8393391290fe52b4eeaba8c0b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d8e0cd983c75733a2816b9d68e57f10f5d3f0ac3245116f0de746503f1090bc0b306f35b4806c80315bec2a30a15a2c868ea80c5ff533a753b0559f85c09cb1e53ad83b0f7b21fb776112e0b636965c154536cd2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4b9654f86f2b07cc12793b503028c8dc89c8be6c187f1dd66b9753d66f32360397868bd158c14ff667121c506f302616cfb76d441e666e29bb3e39118727fc0cc0877833e249ed0bc997eccfeb1b615ff0349517;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f4480d487b9a2c5898141ae67dceea08b860a0ca1f082ed31f6c41780dfa45ed1bd57d8e0864790c458ef3c7c55f23485fc9af58546d6fc78c68954b192bc1ff6d23a7c63bcf95e60f85fea4bac0611ec4b4cf13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h945d77e1af06b8bad8c1704bf8a0c36c3f4df5359370f08cf681f59a8ea0cfb8b8e5479e652c5286eb7d54edfced120f8b23f53e517725724d2d70f0daadf68e237027533036b3fbbd2de79065e1db99153df6826;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ce7c3799817930e4114173e6b18adf2d4b6e442317d3950ae551010841a3868ab5b6128329d26502453ed80b3d05cf9ed3a9437e522d0ac4a5adc5f21c8cb05e31738dfb228ba48ad50071bc8553c1f0afb225ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha169f87579d26f0b31a9db7c950b055cdc2cda3012871f4f04af8d3bc309c864cb59a02e45f947d38dc1f8a58f8ed40130e18fc86bb5cb85c8319d1815ae1ad175915e850785fd13cae078161e219ee8461c7c361;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75a0b304e76be653177c0bec259c3b3745b0e7a3bb658cc643ae706befdc2c3301c7175f586a989c9019efaf6bca6344f980f4a0335cb583dfae77ddf38b95e174f47e41dfe7e718909f5d1a468456acb1fda0d5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b235cff9e18cc5df4821595f6dfdff7d910fa23a140bcef20bfbe2c6eedb68624fe99dd2d0e2690939a7064e9e74b84edf4c51c322e7161d8b7f2d7eddba76294c6931b6784fa449a85f2087602a49f64dafd826;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0fd9cd0fed83b5378f7bbd1aabd465cd7927dbf549b27aa0701e23713157789a80f165b7cc5f46b2126ebe46a968eb804c1527fa53c9525c345bac396d834b88a154f4f7da7db2c8594a81f7de923ec21689f3ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50e58e2d4ccb2c467512aa60fb759101b9c1a806431b9b7d02e04910fe2a34e0fe9401abd9d5c229ef11d224c770209ea8728806bbf13294281c18581b69f0bc32e267cd49935a89f4e0eea04f7c90de085e63dce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89f0346a38a3ab00fc8f7f734e2ed6c9d688db644d3be6d329bbbb191b05d6d1df4d91bb7608148730a38442fdece0692958ea1b076e0ecddcac07f9327967cd4d5eb3a1034206279df65e99c21d552f77fe96406;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h467cfef44d278b3c53612db4987bc480fd3ad1965c7d9fdea1315769a200674eb6be54118c085581700c00ea24d62d7ae5def648203493730274d5dad01162edc22e7aa19a527bbba6af0e85d383ba9c41c4e569;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb7b93bfca603268091cc3142ef100d00218549c5f89bda13d17c0cad340941e817bb8b68ba0551c069ea46607bb22b137f11113958e210fa133e498ca637b437c7afd59a69aa7cd8b05f6480d9809bb716a74f91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d0b049f0f7acb88e9884c3d8676ed65361d8b38ae3f60e52417111211a661bad1b1679c5f55475ddfad5744bec36e99a814f7eabeef2e8db5f2734ed6eabb96953ed898f04f1dc1ef8b7ee3a0f3ac4322fb83f74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb82d609c97d12c09cb7b75117f83c000c1cfc93dd83936b423aa1c3297418d1016197907e4a0f16c959749703c4bdd219b0413624702e92f7ded86a96673fca8066957967a89499eb02e09ca3cde34bbc3c08b7cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51f4ee31a90ba8a92f0c031d34eb6bf2530e4727edbd6e50932198791183c08d8610854cd262c0b16619aed716f0725931e650b4e6c0dc2f07ef6d6db2bfb1f13c129a889a35362417817b65247c00168bc659da0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87c8897d7a177f9a5e0c8fe4d243a46d6e2fef5cf86111369eba5c71d4da7fcd602e6484ed5963da57bfb72c92391d147a7d068728e123a68151cfe5cc78103a5007bad9f06fa88d5199fb908ca99de4b94244313;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9ebfa9a685442bdea2cca8a1d5b98754ac9dabbeffc11c23b2ceb5d2748eb23e19f7f56a6caf76cb9512491346ac1dc61724e7867e735153b5606f11f7e33ca96189c2317ba10c462f7d5109695134b4a84076;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cd73a4d60e1eb93a74a778a8c25a416d09b677fb10324de6894049bf03621ae5063e9ee8cb5f603da802699777be49e32419099c98ab8484127cfa98958b13ed57886c01319ee6f38270c47fd0c37c48feefc7b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f726d14a166c4930a202a7655251b9966643f749e41b114e603b838e22927111bfdd68d2847db42da02ca97cd931c0cf94155a03875933313e6ccf5667837fff0e4e915cacf4dd4e357eca94122242221d68e56d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9223a60926ce5b72c9868a318c24de4689226b6b5e7b274904c55806948d1e60b98b535f36664d95b28caddcc25a5f6b8ef9ed15fcaa3da9b78b9468f9610c1a5375885777df4b19b43a092de7400385fa95b685;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10908716004373ac3f046cbebe8626460dc6bbe5c9ec4c1af8b7c65e0b58cb82f6ec89a48f1847ee8000110897d865a4622b4f3b46c30003d06f8cfb32dadd8822817ab31ce179bc1d37580bdae14586a9d54d60a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28542e81989059df7de9d123becd204f6970d98393b11a68fd10e84c5c7ea802d272da6dfcae4f6ba365d6705b3486b192db8f4677cbbdb169392a3fe90814896f328749c80166eaff6ae27cc6b3f35ce7440519c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc226f6d8699b286443fe748756783c44d2de25e75f3395273500412ef22cc4261641ca5856662e667ec1d2710e139290bfb3b7866b96a3b85263b1deb81a836f7bc486940cb1d2e272e015aed11848f4319cd33b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15b638ed20e8decee877c9e1e3b9384b69f7c5c8fb3e0c1f56dbd7714ff9f29cf47d0da2e4945df4d7e6ccd515e2154604efd0f18c28a767d10c8219101f81c1b285d4ac19280bfffb202f171f7281c14d7001e7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf831bea83cb0a6c0f36bbdac515752e7becb655073baf2161c212150493a0251153eb98b1261a61c14544d1ccf1b11a38bd7da1bca45d9aa933f25d0213c329db61b7c1b173521014af37743f5856584799b71690;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ae85ddb5d0187bdf25235fee5e15bd716e6be04aa69756b69b3b9888dbecd771e56818c2bf9d3219dc9a84a25d37b2aea0f25f160090d4460540ca7ed4ac04e2e94a076fed9d6b529ddcaeeb765a6e5a870bf6a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc99a32d7f1793b8d67f784e7c2d72226d01b686ebf0014cb9320d9a7c424127ec13188eed8a445d54d6105383dded9ec21cc5e10647e2fbda834e8ce91633abc3b903a7122ea4155a1fb6c45badf0975be75f1e05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98cc770e534eaafe6b7aff7a8c80fe75515fd94425c3775df61df1f1370c892d0225539dd74eecebb0291791f0705be6efb598d8a3aa1ffcdc27af449470bc97ee61f7cb847392925d870bc5d4a49c3341e9a4687;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb66756d6d02f7a099cbe5bdee980670449e4cf9cbbb2e806274cb1f4f60cc00a4aafba2278e29a2ab37d8c807d04cf8c5f5df837eb38bf0d261f4d9e3d5d889b45f4390c31d4fa60be738572b116dbd8e4dc24775;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99df292a93c2357de7fd9f9ba29bd28206b484467e82146f06e338a840794b5de62e72b205e3a6c42b9b54c6b106d3154028772b736ba369df7c964e89edc2ed2e2503e74d584a4a022046f0c8378225eca8ee93d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdf8572b81b8feda9b650633a9d6e7cedbbf7709f6a3c46eff3caad6abef040fd023772c29c3397df388319ec472c7e3b4234bddd47d29a4dcd63dcd03b83990034146bea9ce00c13895be102e9b26e083d16d2d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93f72d663c9180bf5c63428406de9b4528b05f250723e746c47c56176ca74a5bae1c9e46d4b758d0b63ae2d7db0c4c3aaca0b00aad8c44b702f0d3fc7e7536c08ce5c52dbb13eb1124e572f60cfd42b09e887145f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3389316991b5b85ce957bf5300481c10b1cee41d7be19d02944b834a4cee084cf313a370762d9c9b6d4b60bf383ae99f542a70e1f25514dc1de3bea30e8093fd2692640df58e5905bb10e8c69628a13cbf50c228;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ee96c90575f6d87ce98c7e0868eb68d7d00a1b3fedf57c52faa9f3719bc214853d1427e235189cec39810c4e142ebf37b45a07c1f0aef5fae5387854e20d718f5c7cc4019e6246c2e7f7e67a90287d5ba757e10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12fbfbc9f62c494d3c52a98c14787f5b53fce817b9d7e573bfeeb2f543011f6c44811c5189f9a81ee442ff0c351fd65dcdc1148e857405c97a656093f002115327d75a008e1882e0f81598b9e66a5a090397aa432;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4d07a93e15c0485c9ecc3d5e1e441da4dcf5c7e84b5833a75a7826b90daa5733af8a9e4f89057e7ccaf448053c65d722ed7a1ff0ea57beff5b6a4eb5c1e7e0d96052001d04ff0064b44c9cecbe6282b2e4ea50c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h753c0e3430ebe19f599270f6052970d1fc94c5120dd85b64a5f07376d7da520f287365c038e99f81fcaea52ba44c62f72f421d04baa36c7023f568ed745e999e9a12130bc6a90c70a1b7a8874345df7440b0a67d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcce44bdb0f48131e634b21a75c618c9df0da88db19a486db91db8d4d26f252dc05fa34c300024029d3d2aaf4da5b36371c16b3e79ced2d6afe2b4add27f7a082f80182da94d9e3223aa62b2bb590dc9052ea23b33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc95fe2db7fb48f1675f9300bf0b7411b9c2f617c927a8a97cbe786b490f2c62eb2b3693e63baab976821dfc2b3d738f2c56f93f6ea978ccdf05ba5f4478bbeb2b284cb66c199217cb588adfabcb5a4b8536652d51;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf224716159d3575a7a11faf7e4dfa37b6b10cc45844747617fc8a96daf49f3df1447f5807fc77c24a06cf047e4b195ae1dfaabc30f5c71af962e9ff15f9f3a84ab75ab52d202c095c2fa77f6742ba1d63d1092f62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5924bee2cfdde9c5b006b60499d744cd43a753713cad792a93730f6ce42b076587c1816ff80164511e66888eabeb33794750148f903410767a94aa7f239a826b8bc5362ced4218462625048918193739de3c5d76;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d3b8ef921c8f7f6c63b4376f5e7bc24b3df79aa771610b53b4e0c2cff196c249a0b30f5f226176b1d1f5425dd42c15034c475e640cb28f5f186f2c551c3df37798487979c1344c449560e4bae1fe6cd3182207af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6259b18125476065c5a424530b1a2a4d9916859ea750c6c43e1495a610082ab5a052d1dc136464229d99e5e3cf25c9df04acdb82b3fc4d8bda6cd91dbf53ff89dcfc931a66a833cfe2dd0e5d6d1462ea7e9e307fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc23fb2a2fddb098f3372628ec0d24c4612ba9a80ef6492b537c2e1614280c7b8891f4e5cca91d14b7c18decd6b67784044c62288aecc69de1fe00a8f8621ee259a3d3feb4361e1c5acd47ec262c688c6e5d5b12a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87778e2289068aaa6cbca36709396b7b3622aab8f46901c3f724e8ea74db6e36c23f3f18c461cf20c5966f6ea9193a0dcee139fa6df5ca7f1a96db4e2a03ba54ab2a28991cbaef42a8dfc2f72e9545742768b3dc9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafc08f5036ee0bcddaf9f883244d86bba00b29e778c0c7f289bdcee84610c67660bc69679c6b00028323a99038edf7fbf145d02554e72febd7161260a1f66be1c8b946c23d8c3fb1a08721380f54645ae7c36a94;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9b6f65a8a722ae654cd8cb8872a86a049e4f94ee787ca5db99875b499b35e3e536bf2744d3ec3c6beeb211ed790e54f05d108a203d767063c50e70e1611d95c3302370a2076ecd1c42df7dfcd8890f480bdbaaa4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he04149a588dd721306233c6555a707d3ddb6218d34cb57c43c29b75f0d4ab09dd93780674cca98c2a065409302fd565743fc7845c8f04978f7586d7d582d873a1fe8e3b02a899785e2c09948569a5f4d440e30bab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88ccf2bde33df2c17347c9807bf505c0534d0844993d100168f5da3854d58b7a723f90c34be973c8c157e51a4181a6bc04b65637348f0d40be4cafdf582158362413128268fd3efbb08b16e1512bb3a81e801f17c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hede66df41295b9f33354ebed55b9a7dbcaf4e139564f00383a8b2384eacce129a2984833db3d253f5c9274d404724e4db7fa86bb2b948580f280e9b48db2cf712fd5d71cb213a4e9e553a52535738dfc2212c6248;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bae0888b36b29d1031e0146084bb3ff492161ac8dad04ca4e8364ea439599860c44bbda139018cf148b37caee25b1a1f4d8d191fbb8cad1d46fdd2ca9c96f5b46cfba28828e440a092f54d8d69cb9392845c74f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c94d254e772c70eff1a38c0198c4646396e3bcf47f9320c0e97993bedfe09579dbc4d93bac2f1e4d3c7777965983ea3d9e045c21e8c42f69cc24faa9f8b50ecee897481cbeaefd396919b3588d18fd6197338815;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34e90ef0d17e865356c3552992137a91ff4fe393a56017098bc5fa36c252e41fe13bba2491f051785bda28aa4f0ea45a9f10a44c5373b8ce32037db7c36117366cfc1fa3bf7d606e869ec66d4f353dd6e87c9ee6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha913884a30b5a3b0a6461bea8d4679179e9446e9a065068e8c3e6cd5d3542775b5c487d84e6b7fa46c877d7940859ae9366549a52e367bd15e5747bff24a8161447fa78d3fb838d574e63a82ee6dadae75afc4841;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63cee411225e471a03f3f847b2822a71f9ff5932e25a4dce947b52d5047a1a57dc4037ffc602067a0183a3ae60bd1649322e389e1bf8a58b2d0574e903277a29ea5696e599d9ab610b85ed8700f2f3de0388d31ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc35dbef9fd0972216fbafa56560a8a5d73ecb62f6f3b5ae97a77bb783b34dce3978a206c9dbedca40d128896a17e08c45e1d2b110b1254377d501ab2b4d65d6f21a1a26d33b7b90772c8dc42c99bce988b5ac06bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2404d298ff244d2d5ed7e75f257c280c8ec1366769b027d087ddafcfc01e7b9e0375ee13fef13975277d5ffa3132400a1eb5582fcb8876c132c308e6f3efeff33a552d7ceaaf4239664c596c512166d758fcb04e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe154ef26bedaef456cf896ad6cfaee0ca0b02ef8dab9a42e4eb4a2e5b862786a70dc8e863f0c6ecba671c54b7570c5af315c34bcbc33c88fb10e618f8bc094c51e158987fd7fb9f1bb5cc99bb9ca00f965e43aa9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70a80b4de39d0d272d31142f6ce3151684d0ea4f7c912950cea845bf19369579d8cefd23ccb044593d9dd6aff0d0a5fca5a8c680bbf7011ca253a336e661c17673e62e878cb5683e60f190db2f3ae24eae7653842;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f3b196a712bd22dee797586b1e6e720c973665e8fc03ca5e218ba366206b1183f121a1cc40678a91a9b80249c5a9460631fe0c364c03926f9eb34e32db6de73324be2fc40f03c5b464234f3a6946830f1d42df9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7466ddd0b26009a2d1af41cb658720e5eb2baf4b691f6cfbc10493d3302d5d797c50483a710dfbd89695a8f5df9150af0b49e8349c7459142256c25541415615c4176f56e1807ec10f692d0fe6834ab43f746d1d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0ef017fbd4d6f6863e3d8e10414073108344eb808d1d8bee1bc5a419d267ed7d294e5ce06c6a2d233bab5e5bf32fb03a8ae74c633aed0e2487ffa094f87ace1964bdecfdfdbf194350c2fa15551c2e127083d0c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff10f10434ae4c700911590fd3cac10e58123700cf5f3487294ad2fc88d1250b22e57c909dd5ea67076c180002a18b48d5046067176d1642beb9c4e4fabea46997a1ceaad3e11d16c35d75cdabd2f831fc6574954;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e295c15dd7b9985abe4589a45bbb5794b3f39fc405f105b9a7255493ced406efad15cc63aebde79ad48c9edab7d9ee0b4908a1fe0f9a02e66c0d6a689cd531407388c00985741c7a113ce8b25425bcd9ed5d6885;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8b75908964212204f5696a4dd87f1fd213846dd0a01093b32630733ae0225fee39d73043dd4180ca1fd7cb9bc33e236af91c53292ffc152022be41521e7e0a0e0dd6e4283a8b9322917a2388dd0f25b95629313e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc522e25eff60f7f31fd790a09523688d40a51254edb794840549b782216012440be2dd5cf14f5050cbfd7098681e6f068355aeec3edcdf1df5ed185a4312a4262c8d546144c4614694148e53470e92196cfdb09c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d439f8a5473c9f80758d865e83c96f0175fee9bfc3a13c1ea6649a9d8478f35b92c034ad3cc3e7a40bb0314e700b40afc1cdfa500f5431672f514282768fbc7c4cc67d3c048001dcdcb58c900f6d1cca43c4f34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35446d06b4abef25cd8a1356fc976d8169c88d26c71e7ff7d7caf64aa7b683fa8f17dc8b614e18ecd0f83a13370edbef9749483ad6ed5a2319ae5bfa14e3a2ac224f3d2d872ca94dc0e2b2faf40b25d84d4c195b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8a80e2ecedc40b1cfa7c6bafead1da4d74f1737f35c6abdbf2e5b66d588efa61985fa57483ed9ff361b1c6e0a89f32f7c32a70b6097c8edc36e95212a5a908a2553640d21f518d7eed5d68c2be62bc60ea555688;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e81288b6d36dd611771eef2bb419b8413afa17f02c94157582487326b5e628c984e7e4bf1a8e84d6a8a25c9c8e13a15258062d7916a8c5e087bfd268a6ec47dd156fed7c2a34907b38610c05dc8b76e5cc30b28b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3df4e46b9a89bd96e32c809f7d73ce0c604a35f62d6f9d93a51f7e5f906e6d99e5f8b5bdfad3f0b1ca1b71ea633962e2ca92c9fda5c6f79a2c240339d7a102bf7d6ba4965a1160d6656a23b6cc39382cf7192119;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b025613876ddd5fc139b069fff39c05d6e12075fde46f8b73231678a0d9cb203128cd583286282bd1514c685002c41209e2d4f8dfe25cec393dcb061f0b7ccc99cb5519bf8513a44d81024d02513f13f8e6d16a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0cf8bdc3fd99297e43647a0165dba34373c07ad6ad62ec23e6527a9c35195db9410210790b9a6d5ea5e27a8e3c56a190619e1453edd5450fbf8710af96fc8cff3499394ad59d2ea630f4629e7fcc46e819d711de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6a8fd7f9aab7d9ddd92f670bae489b611deb556784a2ec6a0d4cf4b46357908c31931ecce595afd702c22530633b33cdb23f210e99f8b0be46f5dc09037dfb949d25ea2d8775f2b9e12b07e2b1c0a6d8e6101862;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52bb9e9c00aa6bf970ec111c363495167197cfdd886337bde503894b4bf59cabf5916cd2f7b1786c01ee7484cf8eae6f64fbeea3d0431ef2bee836e4d0996cefa96e230220ffef089c73a2d0c3aa905ef325d4ab3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdff4136e91e34799e9572dc059772c2a87abf6bf2e298955b06428fbd1723b58da375464956e6f555ec4fd7577c37aefa40a073e03a553933db54757ef320296f55cc0f130202ea71107e726f20c826a9f91b4111;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2be2434e779291047f7714874716ac8e1a0c2213681635bcf846980c76fa3d1d63d41bbd8de61e9a67f5ced8884a8fe2992ed94484642e40015d6468142a939812a8a25e2f4ba867df5944cf9776b3b11b88921fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0ab7d01a36652b0bf7452f014f221c6ee8d96581efa47ad0a4e4fd10e2d099d9b30ca1d50ac7886d3c14ab4c09a1f865d9fa46e1f515e1a98a431bb21d91deffb02c26a66d9595372a52659633ee68697a7d2dc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45a8afcfd0716924c6b16478d8b1ad690cdc2025980eb719651c57a52465021c44d25aa2d9f39dc08ec1768671a66e0f1e8295161bb0d3c332f1b3ecfd4b26b16f06be1c7330ac2b5ee7b69c25fcb7af0261c6fb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1774e99017bdcca949161a33f0efa54b839731be6243cc868732b408417e1cbe2ea342376d2b482f3cdf33e4874cd4fb236d550e14d8e1839b3bbb0ec7fc4e2368952eb0d1d1acb7b363cf6e9b45b931c4f513e57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa9f7ba288b6ad1124e105b3e5c310c4cd453c141551b33a5d60dda53df7196c6564f69a41d4daada6036b51772b44f7ba4f3d5ebf3542c5cd1465bf27a2f767b7be03e1f35f29ea8c801d4ce228773777a9b3215;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8905f5f5d55f22e0fc15571a04513a2667616d23e97eeca12ebe4196ad535b80bb68d4772e747f2fa14e88ee3a967074f10cf38e6ffddbb2be40201b4e0eb4cc189228772ef70febd35a298ef3037794adb4a9a2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ab2fe8453e238cde1e22e4109bb96273113a294788688aa10a2d7137b40aa2bf3472f230dca2e1903428a1bd47d63a40ad1cb267ff977d1cd786ff056ebc188ceaa3f23caa9f92a5aba86e96069a0453ebd1c981;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c37fbf050a748b8503e5326a18c91bb5f36d0f825e058154eea8d9a383e4cfac7b8db91c13cdbd5e8249d5b63dcb06075ea48b2e3044cb613afb1bf4fe8825035adc388f61bde25c1392d15963c598cb0c4658ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4ff397c365a11142424c8f8acde7eca36cfbbda9f1d9d36873b07705bca41e19606428c5b1de666be5eecf54c62e2091c6eaf271817db0d6077e856e96692ae28d5630bcff69dca2dde6da4671071f99dec8d33a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9b1be5217b48136e9448a436d8ef2005f5e9771cbf46ffc6c541b5f17c8d25fa7d5fc64d2a39fbd2fc8c8f885fccea194232ccfc8f296907913c8fa1395cec911226b58d6285edc0fd5c71f6e4b9e12a7061fea5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5f66973071398e6d0b1a7f92da0d7358035b8bec9472bf0d4961374b16885da7f7032634f68cf68913e3ba46f96e827ba28b9e9f27069be67cb9fbe53f56310ed756be9b47aeba8a08671287ca5d3ffc192285c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8023bb3a8cc16a1dd2feac84026f41db4adf89d23842273a77256a29d26b6591340f26915d2ee04c6669081f62cb5b2ea6f0d072ce6dabfe50d6ec24b0ac85a2a9746d431adfaf0bc8e898ce999ddc028a085587;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haadb39907e1ca3d1a71ed285c0de3e320f4e019ccdbb9be3e6032443da4c0bf2ea7bad698e6f363c1733c8da4c3d0fc0f0050530dcbea33e086aade5e8098493fbd65ff4ff755af28e610ddef468dccf2bc8ca9db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda349a607990cc970c6588178195e4aaeac44b28c72d61f82fd89d15c9d245a784325abcd4bbd35a7b2b1e2d171dcdf422addbcaf17ab2277fcb6a323e5f1894eb52b43ccbbc119ac128af1d4ffd323f4a0d895b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb51fc5161c4a6735db01f0bf2e350c93f73a92a982bc2e11fb50ce6c47fcbac35079edb24ff4bbbabd0396c39fd9a3aeb130d99552dbce24ea8da05f14858ac0d9a40312de7230efc08fce2daf05107ba883427f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4772ab2b6d151fd2cedf2cf871589811c623305c1fcb605af1e6c54923c366d056568f6859bc66ada7e40f2661b380fccbafcd0e555b300e7a04e4e5b259e84650a2158632c238449e9f97d6f38aeaa1c2051e49;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3eeb9229155ad57f5ee89c4803884fd02dffb581a57a26b6e03e01f76a788ecb3d0f483defcab230fbe96d6b4df733acbdca4c17ee6ea2b6c31a297d1a85ef84d216c5b0edc6a19cce16f79720e8c772abf8f6f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef55f50af4a670c8cd692106f33a104aa07080d8b9804aab76ab4a350e592889372faeeace571c493a189869bf6c9f76993c06e848a0c0958c9887730247183280544004bbe5810c5686a390de945f800d2cc9f31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec5c21465bf67e5e66915f67f8ab545793b28a04830d50d50a59a91dab2c2a45c5316145dcdaf708c87b854573fbc1b7fc7da50d7839f1ff9cdf854c5b1b25a2a7270a8649db37a8cb992f73adc1b38622eaa40fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb340217ea6ea26aece7dc19a046b0dcf743fa25f3173340c037951589a8da0da278a64859cefe39a95e1cd80939cbd113753060c72b57425394252e363e5ddd784f616bd897995447e723b5905b18a0c3d6d79696;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d128e9bc2ce2029f39359eaa31778322aa955ef285f71012d0c707339f4955d639f38eda988f9135c18b48fc9833f5c63590030ced64e6e4543cd1a1c902f5b0fb217d007177a95273c124d244812cde34988476;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ec2bd19e8173538e7b9001e49524dc6c48a0a7f623388fcff178108ec0043fb77301bca5188e167bc21a22378b9ec98ef092ceae22e0da452b951b5dd1b2f1e152a251c55334a55ab7742d51377cd8f1a9366fd0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18ec1f49fd63f9999342ac98a6dcc9fe61aa38bae051c1c5bcd1531b9018f88a20ab61bcb6054791b534c678d24f15e7e6343960ebb5a15a0c2d2cc9f26948b54178d4499282a7f6e0523a8712675a7b361c82b68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb48280eae7825e9bce9c94a9861d2c1566634009278434aeaa8d0f9b6c9154cd83faab84541b9f129cc66c02bd64c1c3835f9004b1816dc2bca32f5894e137f78f6ed0089d6e6a9f54e59267462951d1ee032b346;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50deac907a75a2682aa57fd8b7491b821f45f8bb25da0c57a0be5751d66b999010f773e5fab8e18a198d4c31122c46d159360b8bfcc7c5b454a1ca210da7642d000130eab9a1e13707533537c0ec8605621fbb7a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a4df7e0ca5941f6b5aedc749787ce574b0f860344de9a382b0e0ae1a28b831e7d923fc16c0ae45997e814b88375bebb6a5fb79a03d6fc0f1329cee2b276cb489208817f85dbe5728ccf7c8acd788fdf0a4f9d015;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cc514ab3c4b224115403c80af83b4183fc632bbe4a51afa4c51aa8540c797dd85d995251a6b3e694b6f28090a3cd18bacb4b1c1a981c27216774acb9dd69d9a91657de62a2cdcb18a96fcfaae18e3049fe128275;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40d3ded70a4ded24dd0e3b3f04ff8833365022e0179690ae8811f45e2b94e3884f2e6cecbb33decf8dfccc8bf14b549650761071db1eebcb3d91b9037307469d849e6a5493daf43577752c17d593adeaa5fb96b4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5097a42daec47d33e09bdac6bfece5026e431aa80f8ef68cb7cc8047fdc80460aff577ce99bfdd4c3744d04e018df123dbc904578265ab507610d8df0669e0ffd1d8725ebabcda9599bd384bfe06b9814a7316a5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb254eaee4e2db1972de61f678c33f9b534e2491d6223e893973db4be3d1d944b325dfe414e1c930eef8c35b2926df4289e5aa00e01f038f29c4bcb820c96951dd1666bc6a7d427d7147aedbe5cabd51dff9237ed8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4232a6e395eb060e68ee3407704ed9890affb695d2386e5251d8dea2d4c047fcbfb4a6ef58a23e7aa16f9f240272a05bba03aac69fb06494ddaff6cdefc26a016a343b184bd9487a680e41a76f486296309098f25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha960ae454b9353b44719a0ef69df259b6468ac9a33298519539a21cabb0da28299c411f8bf7605a31f919fa971903d280fa34b80fce2a291f13825d264ce72ef4aeb3d499d6a8e7f8639f81998c24a190f12f5299;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h743849693aefd281e4f6df796927e35bcb82e6236136d92bced95852bc78876dafce908cba42a5d139e71843d3fdf37f5bb64303f5bdbdbcc4daed6b72c2f3217e15daae1f020ca2cdae63ad7db5002d1fc1459e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43bebddd6f8e6e7ef0969be90b11bd9fd0e19f69810bc223811df762c727fa42d647baedfd96f16e6019c40ec4e2d0bbe534c24f8c1b770a9af44663cef5ad4529c628bb2b603b5ee33dd6a458cb487ec785658f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a3325d9460ee4b24320b25d3dbbc1a5015cfef7c0ee8d241074a9f91c61705525da1beb4f2e7ee4c954f82b7675d54cd42f1f7fa37a3e8001ef941a9baec718a67748ef1931cc8e694c30b4de9af9f83a4b21407;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f5cbf3de84b5ca6eb396902c5a575424e6dd859ae18913e848d97075f0a0b8a010377330028a8ce42d77598f3643b960d8fcf295083b33c5751e569a98448760dd744b0bba11b49b368d3505e544cf18dfc83c99;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf842a6811a56614b761da149f17ccdaf0694ab8df3c9b8b95be9725b596dfde7eb6cd0cf59167276f2c6cee59ee949aa2297b803aa36ff2be33f8d76240ea1b75c76cb176cd513d38dc63b734052ebc06f9942ea7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b44a803f8b47924cf6fe6a0e800a9aa6d320c6d81f1a61b80609d56a91ac6fc293790fda5a6dc16a6d2741dc89463384491dc114068f30073388a8a8a5d97a709f703934a8586c3259db9db0b39715801d860923;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e4af576f5d6f13fb31a377adc8b8f3e76d6ec26fb32a26c43ed8b4540eeb6be9c5af2f2046f460378277efc47c1ca73fcf7c47184701189c1cfc8767f3528b6d77c80f408f1591b8653cc9903f94c72638a323ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee555eea0006fa5cdb54d59c436c4ad6a8861663880302eb422d0f9ae00639a7e88f446c79f525967c6d3f6fc32898861899a48ba5e3a9104607c74eda1852c4477921887ad67581d1f0284a02e0315f7887b2abe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31c400c99d18205f853cbac03b6848c5d6a2fb48bf4b0750c1dafb93b2622505173a12114133507d806eed5728de74f326fb3c54fcb31e95b0b4bd724d59987633c654681a23995a67e7fe31c8be9ee706d002ec7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb738f592fe2cdbb598bce8ad20a41ff98291ed60ec2afd8342e93ff27d29e97059b37b7fe0e43217eb6834146f4e40448fec4692db00fea40daf3a39f5467a4268b1a53932acdfb768cd727e42f67b581f56a9ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h864683ca8ff3b590a5979614c550b17473d578b01a59c8b8160adcac1ce6ec32ab5c3ba3f51985dc71618a1fe74c4507c5da3365a6da27fee3809056da30d2077e6873744751600eb3455c026aaae82e61d4cb7f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67a32f5e65837a47e354119673b36161429016e0b937d947c021e0972eed6814644536fe9f517d3e3110d087968f3ba4a7288f300f7e15985ba5dfe97034aa64a5e482700473680c15d999d71cbbd2e92921daed9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2765bab405cec92f5ce551ee08b61eae46704e72bf813f1ff5384c354240dbd87e0aaead6a7a7f59198bb799cf822e242c3057319973f70917d430cbe25bbfd961e81cb397a38342ea94ab438326793c4e8ea791;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb07249e3088e47d824a858a95be74c332a9063dd0a9748f394fb9ed40361983f26236595b611fca9ad166424a9f10b67cbb947667ca327ecd15f236b7b9ecda478fb2b378d57e49246657aac345ab19b10fdc3884;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44bc76b60c57cfda2fc9d147a0456a52979bea7f5f07a2e1d99ceb1aac69e8e3e76a9cc2815b56da76300958c4cac0451fc2e2b5365ddc11aad9e0494467becca1470055871da19e78c06d1a4e8cdbf178ab458a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dcfdb1b8c932bfc303b88638bf4e192670052f1963491f427ae6a3615177e0bb9e4fb6a28843c95e0bb18449c20d5c66561721119929142a34e43685793ede492ec969be9918597a47fa3dd914707b689a40e7a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12fc35137f62872a1f148dd16a12038b69c14641cbbfe76138868d8d74d35ff3610a88e0de43c06a31acb4722437eba395975ac7d34cc4f59be27e3fcdfde73770904c7af8d28a8e4a51bb24e12d751128ea12ab4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98702e4e80cbf621c9606499a90f6c0b1f04edad4e3673e65be9585dea2d147728a6638f6d9b4a858ab40537428312283839764c83f75d88cf4ed87a71da01536e3876d5cbee9b7cd2a7d7f5eec477db5d48f01c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3092f022d5dc0f1e412d493a3c178d6f132b3011b10146a9d66b792a7a074034f3ce77318d88c3a9dc04d12422e3be851426d8bade7eb5050f656beb967fa6eff4893d3c8aa5baee4805c860fde0ea4ad2e8e6bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7eb46acae470a0d887c26326da638e22299ad8e16360652e0d38240b767048a5fe79dafa8c5e72a93224c393e2ddf168bf13f716e06ccc606b20f6370fd961619daaf93141268a53d5ec51e7c084ab76f055827;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96398f94e603bcde5ae07ad04e51e20e19130315d618ea281d7dedaf15cff8e44be22c97b52cfe0fae1041076ba7b1f46eacc470d41062574d29550fb9065757f11472c14e509b9559027bd5b667c7cd3f5bd48c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94c010c031f83b9050a4fab846b03d03bca9a551066727b0126b6292f19198db57f7164548b01a3640be89eb3c2a4cd63ee5db9c54e289da20d37ead6c8095b5e80784b9e6da9225ae77f69591c4ffaf09c5fd178;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a8b396e1fa379e7d83387f7dbdd6346c25f0ab124f0bf6d8b72ea26e8b6ad5dad6db814ddaa606fa50902040e349cdc32e76a66e75d18a0629e83eeb4a2907a82e30d02f0a75d4f0f76634eb6f3bebba5986f2b3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h486f73e6da33a760f1bdbfd378577449266f385a6b58c0a5a1ffe55c03a8c2d5b84a4f727bf06141cfc04f8f81c44ffa8e0d6fdc9409bd9cbc7c24b98c56e64bf197cef532b0bcc7f46d84c38ae3827a27c4b2c3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ed9475babeab4e7cedfcc67b06b13efb667b0c621d2b1ea919e03bdf07cefea31499cc27660cfc0427bd99afdf1b06855a0676930d2f8b2b9f56c09dc4933034b04b252b3a4846a1072a68a0cc66ef32b0e24db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a56d5538904b0cdf3507c8d8e3a91649c31d98823a994381d42851905f2a0bad98cd986a54716ba413d62cb84400c5146c561a14d270cac81ba13a426a2dae174f479a9fc7ab5437d9cd2d39034955d01ec96fa4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4789e23da1ff4dfd5d38b72672d51fbf8fcb273871ee67f5a99785dd02e54e47ef26e2bf9fa642b04fcbac514bbde7f08ad36ed63c64ec186191f0850dd3b6fc255bb0f78432095732eceee968a4963e11a1f81f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d1ac409d72f1df51322c0a21006e1e94454ec09b64e039a081316ef42f5cb157782dbce77df096ea8041d97796970472543a4f0c62551e6fd6dcc12e2251fadc890ac3648655dd88b73459ed8912628a6f484929;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9eee8fb65573e64e11885b623906f6d848b1ded1dbc7d030142447bfff20353f31bdc1e495c7250114f309ffdcae3afc7e94cddc392e88990d982b360853755f91310b48571c58c1698d5730868a0331d7c801e5b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbeef48e5148991c84b8115cf5dc7bf5264b94576294a61878111415a08411fbf8826d74532d2b0005a612efaa25ad8d7cbc76810bcda09c7f7978250d2ee041c1aceebc361a1aeb9b24916597e30e127610dc13f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dcdb628bbc4fa0f7e0ec347d11343ae3107fc921328f38caaf14066cdd0d1332033fdc2d2b4965f1280ef6bdfeef54090b8d99b8558d48240d531ed3cad89d4804220fc2e4b59317b9d3a03127515951833a024d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1db26830a5d1d119b6eca0c17e12a8ee4ca0c9ee7fa4e200cf40b48f4f9ca6eb9c75c32fefbb45bfe705316b561401027f7374c8f571a12d0aad81574d47ac94d26d4f952e3bd73ac49a18e78f531c261cad3e4b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e5ac4e435ee7059771f091ffcaf0dd35c7f8a0946046eb86f6d7d7578e75e8926eb2ee63f5f3b1f3af3fd4332096b981a70ea064e5c4834e5b6733f12eb320488ac9418a5f6038a0b389d7e83dd45e2d8089053c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h670b6ab450e1ec5413dcaec7deda08f8bd0563cf0a722162cdf00eed577942d36778b12bc952c2d0631467abf00e7a98965317c6ca6a28ccd1916a7c62a7bbca85f663fb4ef6e1e722497631b5f5acb60c325233f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7603d76b2dcb3d991a6ca37ba7b8be5aa85ca1c8da9ad8a00b32f779b750e641d6ff9c362a6ae5f154cded68e633efb3d2c127e4d7a51f3e161060d052d63087ac2802ae56207c1fed2b2f552c59308155b918581;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64ede57d5a8ad9c2180fc0f5b5bad83557c79dcff759f59bd2125fd74f5ed639d85ae2eec0ab71a90cf2713a9bb360d6fb3f872d766537df840590a8acd38e1a196db1c53a53a35ff9bfbd0ec5baf764124ae49d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89b152c8284195601f1b5b104b3ed9911b06a5d89dbda5770a361276162953a0a9acb767cb5bfed0539abae8fc6b729f047108e1ee826c967d69ccddf82187e85811580273800de601a8a058c8751fe1fd89b8b7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h310506c153c32db63e2472b298b5f7544bcf74aea5b508d6fc82cf5115e816f63e45ca20ec1a3be2b05f0ae975f8510671ba4f05d0bfce28b0ae6348a0756f1e14500b1105e20038fd054c3ea6a644ac12650646c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2627990f827a86c33c19fa5cda350618655d3ccd8a9df50a910e3c9a23e6d8b2cb76dc81fbceb32d1fd7ef4e84d07e37176da1b5f0690e386874074355b646e1d9e3fc3ea834fe5f4716639fb0ff55c6e700744c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60aba9a0371412884aa3df454ce5053af2ae96bc2e25d81d7bcf999884a766eaa975b80bc784650dd59004ef7905691204d8db93a3d075a610c61c79ffef76f4e2c515226b5caa9a530aa7003635a07c8461a58f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79d055ff30131b525516c87781afdcff1f8e3e58a1f0903aa07db6f279ed8db5ef0c37ac0ffdf7cb56a0ac04dfd1ad64c2853d63284b01e52a51f2ec684ff33fd216e59e1c9b472c4821919745d9144bd6b0456ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab8e3d028e7e38664b5737c0e2778cab9e12dc27a243bbf8f02bb906ac2192ffca531e123d12a0a0e720d52a5a10e6d98e4139a340b1644a826615892b57674a28a9fd0868daa088f21c4f743d3dfa00677ddb322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4290e2b398467c5a924e2ed64368c11f9608cf57d89be9056e840b78e33a4679188f1fbdded12018b14ab4baa86a126a661943ba15d3bc4d0d68c843928fb0d38bef9ab195dcdfbcf0eda7b07d8dcaa66201d3bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd99bc4f03687ac1a6d23a60c898ee155f26e95f2ac506005005e0071ece0d01a263acfd176335b574636ef097eadffd89164267ed45c50039513df5663943f6eb7272899950bb49e4aad74b65f42cb98a1e3a05f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c0b4429b88032a93b1410917240e5da46e18ab7eb0463f326663f104be2419d567baef7f1a1f45b34a49c3409ce848d9ca6b8310819c7b7a466bda8f5a5b37d23870424c9de87f60a94784901b888cfec0bb0f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdad1dbc190c48ebda4b98b5f51919ac67be4381ed975947ece38def161b0027ebddf969e44d1c97af219610ef7090e83fec3ef1c4046c9f0dd82339c20a4df45087d022745c59797f20cdf37bdbf3b193fdfc670b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22b5140566c05eecfc27ca32005be9b258f9e1d75ab2eeaa78f1bfcaa2b462b6758983c457798d072cbc28e975f1a7ad3105c88c308387021c3f2a6a7daf07555f9acc9c71c34e1e05142f73057a363ccddbbf4f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2b2b545a59d29d73df592b785805aa17f0093e9be5c364d9ab73eaa90d666fa020d450e2b5b5933c1e4e556838ac7ccfe861455846340847142b866df70d774cab7b7ebb95b03290e71cb44dfacb5cbb4798a321;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47f81d4f8cc67ac2e554e984a38cace84df3389eb3a28b7cd9444b91bd62ef3eb4d082861239ec86999889938292a2c18a2f5010cb66f7a638db07b52c7683277e58767972016bafb0400919a2d1171071723e91a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3fe600bde4ef7f70200487c261188bc4d47225b9b4a813224afcd0db56cd37013ce7f42ed4ab6bba1c86cfb0e90b382f3fe95e2eec55ca201787d0e0cfe3622125ed9d230ec015695eb723ea83d41d77596d5141;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa5db9aeda7950bc29414d8bc5b561cacdba401ba6e9e903e5863b4d6c19ad750a005cd9d4958cf2d4ea8b16830845f0d2447e184767af12d7e742f1915aaa801b2d82c2b4a0f3baa46031a143653601b272a785d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e38f562da34382c3411140e09eceecbefb366931319450477e29f5b182e5500d9b59365b827c580033a79ab421a044bd5a4a409fc901df0fdb5807b485c8742d0c00337efdae7ff4c209145472ca632eedc37104;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c8bf80a47855ab0e9d30ceb0c88327a965fa952781864b2692b8c1f7a6d57c6e117ffe575dffa48e3edec14ee1383b5714578e9d773ac12571b911a3d223e611d01ac3c2a7b119e8f7dd11dfd7d7c382e210b0b4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb639413fa5e39e31ad1862234bcfa28020a19bf05ea87576da33db45c2f6042068b61dfc5559b52bfa31c70c604592122bd700c2a2e847039d9b1d562a4e3a83699eead71dbca316031fd802f783529f30bd6e68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73059674cbdf8fe5e2af68dad8a662a064679b652a599b35751c9b94ec2d5125e48e64990af5c267327f43934707cfc9f577266ba06794db7446f85216d6a0bc6ca8a6af806cd8fa8882cbe1efbbdbb3fb3a95191;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc80512751a5d31f2f6c6b19c0fdce0efdbbade6325b92f19bbb30311e5429362285a0d86c6042575b1521d23187c915e248bd634d86547eebeb8c4d3e20c9baca4bf17f8fc8de5aec3de23e913a82751e99263036;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4766519257bc481594a3232ea78f6220c2bc10272392eca9852d726f4b2085161e7bf9e2ebe93f1f9bfa8157883003be7671e2e89d7e7e81743cb51245b2f5850dc87c9fcd24656835f4c6c76679c723f79e2e04;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29ff776920d3bae93583855900ed2a72266a66d76708a70ce5795baebcb6685d9c61d977eba870d8e8746acf288a69109899c18fd95f5bd2c8fbded9351b4c064a6238290cc56bd7234cd81dfa863ab85fed14fac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99dc6fe5f90aa4f0f2f62aeb964c38b6f28702422420e7d48861a267b6b62931edc218b9466353ae51e81f5d4b676f31c1534fd8a7e18e9fe0de5294db946a3b988ae3e9feccbd63c1176c57355a8ac5a5ecf67ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf98fd28d53ad9fc6c670a0f78bc75b3c986100038b2505253ee5819b1e2c5b40bdb0565ab5e4c06f316debcc9c3f553163bb4bb27fc1cefa4761fb2d9a204afef3cfec049363781431ffb23b23ad41091ea9e018;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a8d9e25e2d5d67d665e29660d88001cd701c65860562928cc4aa23c5f68f525cc6b4f3860e658e939ed720a1926711250711bd5499c24c7fe5f26018b88729ec318432590ae7834fb49175bab2a18c2c1c43a1b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79fc71f91d7acc3c6bbbbe040be98a35dab5a471eba6a40e0d74a21d689c2a0a616d996bad56c3e1de06fdfd8aefcafd3713ba85f51acb64290582298da70a7f672ae1a1434e14f8cea6944f0de61a386ba50979a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had1c783f8b2a6171161c4e3d20c236e4d2866b410a5ab70e437aad7b0d5854119e2ac9df76582356d473a6d9aaa310b56c73181d3e3ba18c2cb31479c35b2c2e492bcb193513b4816d7dc070aa5e6e36538acf07e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87756808f55deb6df2ef4b57aca2702a35e15ba7412c9570c5671d3ed2d4bdc29522dd52fb441b5510a0cfaa16c58971bbd63ccfcf8d273189cd86d3167d919eb3dffa1f4a143cd7ef99d4e7e2a5956d2b4899715;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5e084c30ba9184e02df7467eaa97f267781fdcc902cf57b4e7e600396a1019f2c033cdc37e3bb47703584a609aa408daefd027d06e758719d4cd0d8b7750c179a1dd65305e4f8703786a25975984a5856c3d4eb7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf46fad0882210b739382028e791bd63ba3ddfe99bcc0eea2bbd147b9e845674b60a3739d8934cffd4d255ac0373120d5175ac48f32bb415a43cf9ba9ebee3dbb52b4c31a418745351026f60cd0686931b07b9e971;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h870460fba1ed49c4de1dda90bdf12ff1d893018ad45b4893d2d521ce3216a0d02efc9c69d0501f27a588cfe5e4f133a674fd5caf378fa1154e02638e21d5c09f8d3968d1e7758fa557d7705be152357d5b4284fef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800c551ddffc078f808f0ad237c501f29a645a7efa619e6ae7986ddeab1c0f91725647d014c7defb8074fa852702e8ed2fe6a74be6fe99ebc4e01b63141251e2470dc262b299b1023d7437543bbd389ce95f4373c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb865f71919ecf9d2bb9ffd893b1327bd210e2f3b8f7b8ade9faa298b0a9ea465ceaf7b955902e04c94513c77c70f25f6e3d3854af5104b139edb878c0d5fe827d38afaa8ee250e54ff719be16dde5fec16573140e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62a30135052e7e54415dfc39dc4cc05251754fbd2762437307f1540ba776adf81d879e14c587fb1d02dc4dfe04aa9e7ed67f304ead49c2b1242368043f808c5d708ec7bd978528e98fe57ec721a51ab83fd57335a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb5d58f98da4ea7d536e0d35ecf38b2cf6c70c71a3d96002c29763839be1545d0013e08e067d57996c64fc0045c8c5c23b364ee15bef9c252ab80ab765d3b314dc65ee0f23d0ca58a2468046567538b326bacc91e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0b4ba848fb88ef2f619a020ebf1d7c8f7b1942127aa265671fe104183aaeb4634c679d2cfbb75da8e4657b8b15c225b565936a0fd74986fbe8512388083952937a9b478986fe255f6a01f603e394eac7f42d7b43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96d99051a12ab7219241feb90344c9bb8b2cbc1e9f392e4d78402e90727bc2421711d00b372e864f88452654745da2354c8a797d9b1f00ae47d2bab6bc002261426a3f2c5a26635f89e0e0115fd2e40284a8ca825;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4887f760e6870c140d77f5541a767782b3a5c3334575ec9648d6a493b0ce1d75be74fbd90f443b794144f104fdbe88fc769f25630088f5fcd9f465cedaa62aa603648204d26477fbccc7e70ae3b868bc7d64212d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0a93440b845225a26f527dae927e1515309a89aefabd7c73d059b984c36a52877f9ce27fb135cd4b554153eb3813d9ab70ab020242c532421f59e4fc5324aa41181db394a08713ecf14698e8070188ec22dd87bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99c3b9714f30975b8f90985f0d0ac1857eaea68c1b69d3d08f1a6ff86815fea9e5ccd28fe409f0d08e9d029b52e691ba9aa438c742578f482770f2ba634f3e6603c1a35ab471fccaf66bb456e104fa9e5cb0d2c44;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf4330e8b611ea901d1eaf210aafdcc8eed263a8da7459a4cecd07234b78b3dd58e72fe2bdc602cb57e3dbd879633f70e4ba0bc9f4b69972e391a2f43b551b778d7daf50e7a01ab75e9a38f30dfc4bda13b78f2aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd14dc97ed7dc7e396e2f3a41abb5edbf2d2709d0796df9052a29d5311954e32918e22f4b25bfb6d8d0f419ca64784336e58fb07f0369028c8496224518c7471b26854f4d5ca5597f71699a3ca21b15c9b835c4fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69884347f1cf7d48e21d14e6392a3c71741aa15b40199ef72f81816536769b7beecde8db4911e7b62c339a37ad60aa7bf9e45bdc6dcfbcf2585d9bff4af063c169b2106cb20c848ca6aeb9c49a78808174dae616;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebe6429d8a58f2a2c9fedcd88a54328e3c227f2a72ea93cbdadc45a2f6efd5a7949ca11913eeaab8dea9990095b2b2b7c2f16d16462a4e9ddf739de2736f097f059c3e7dc390922028bd13babab5b54206c71e892;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h127cf61bcb6c3411255985d26561583c17412179de508e1c59b9a8e4fa105a3f0b01d651fee88921ac0957add9b79924929a1bc92e4a4f9dc077c2fc64e3a5db2ea0fd80b06462fac8ebce2c8dfcf55a12f571339;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5dcf92350f20ad09d3fbfd6f0826691d28ed1c48f8815a08462ad99e25556a391828e098490c7d816c04c6673bc383e38951e91ebb8c22ea011f7b22da490e5b8c5422fc3b324311f8f207ad7fe287451bc405d32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h532ff5126822701b8e8af8b6308ae5183a8064759af9eb3021170c9ce952e72c7b9223ec1fa8a3830e4dfae3da32d7e7e488d3a31b46532d36807069bce5cbe5c36b1675df03032b24c6b31397c89a00503ca38e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc185653d397c68613c875b27019c6be39ac0e0426018991256440835eb05b6e46df5a11a743b444dab07f8dc7691bbf459886452bda131e4a08a71071b1b0b5bf54e3112592a88650fa85be9e31e004aa5366d2ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb2ddeef785877ad4e6565894f37ec4a9786c66a20d889f84ea09690124fa21ac507a2af95e7e65a60de3ca28aaf9b0984b06bbe982ab75ea711ef6a31b261e03bac4ed7240a57b6b1808438552dee5dcd0fb2eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0201ca88ea25e67d44d7d681bce51ce67091d3ac7ede45f78d816cce0140c31f7da81f603cc18528fb70545f3950ae0c1e8cc41ea2f6f3e12c382977308b5d07ceb833367aa335a30dde955904aacc4db77763bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce1d02d7785dda02174ed5dd4d75aed934b949a9eb875e6bb6d70e3e8b2a6b9f4013d7fa58d28fc3e4d6f5d1c10ff01e1915c2e46eeffe8ad8c9e0d23d81cf5ef85d129519ea834e13b59c6833d718c1d88dc7f13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1a7c542a21fbf0f80287530587bc1fc0f9b85ef4f1b88a5d11a6b377a83d577e59713266beaac608605f8835481b7a99f5c909d03d9bc5880db1412d4fd4de8cab2c8f4594494984a2a2bff6db3f5aeb907a278e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h275941768ac9f2db5bb9705ade8b21be4d0ffaec5ed6d46f82bd9946cb8cd5d6c8665da0e22add70516f97650dfa68597db946c344530c21b5c10ff1e4ba43cea1afd0e2978e5f97e12bfb6cf91a62ef0cca5a3ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h393c13aed5adb6f9a523c5dec6d644de169753a73f405c17de1eab30cefc7171fde922aa16312ed5a398cb473d0ca8f9f2cc8140cd4dde6e580c195dcc255bdea2b84618c5b0d25fc9e148286378d954f10f11ea5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7cbe5883ad62a653480dfc7c035a4476bfa3cea16d36267a455b153328aa54b084b19eb83a9245ae850aa05f144575954753998653652a1d3984452eec29e837235224fd460589d49d451fd5667d1c52eba50aba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc48056b1e49b92c981b415e716514f3b3f5cbf7fa71817a9f630a8adc15fa2b633954bc681c6e3c9c49366734281a160d440325fb48f963a25707cf98a263b3d35ddaae8e83b7f5cdbb0d22ff78d0c05e070cabfc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd94a359ff68be52eacb6b015e3cf9a192ce0a5ce3b3b3ee4ce915f09d49379b5c52fdb5e2a9c5e4db3e84c0703ca3c3e206a53ab5426e6b6c6c0ff01c2f33f783346cc187d2bc5414311ec226f64474712c3e545;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fb5a7415ace0e620eeb58736c39d1c240020624599beab8db14b27243eafe5d3b0bc79d72b9085c13f5b735d5bc7334689f631e19172d2ac99faf03c12bb8ed35b80db58e6ca7be38b4525b19b291189fe1203ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h902a89e93c204cd950f129042a7bac94c64e353e74e39ea19de18f4c8bd3f3420eb92f55d0e69c65e1aa0fecd6da5a8e86e9d95f88aafab6fb1805c2573fcd99827da5d43619fcfbf676c06b78a8b829efc1df4a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ce9dc0afe49aaca0a85688b23f90be002debd3a48313e1dde09d89ae34f4394e5de82db63f24a0f20571378ce4d5a143b6203ec9d6a16f6ecbef60fa95e30805dc5a6b1465334c9f21be4787de97ff1cb79bfa98;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h485112ac7abf304fa070fbafe4cf77732636856cc3c111f2f53329272535424e98e3677e8631012066418889399812adcb70ebf23798e31ad0b8f6bd3fc605f80aeb29ea93a04d85b74425a9967334a84268bb527;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb170e45399d3153d6f553918c17539dfdaea7e6996a4bf23787b831e71588300b3141bd3854ef770b26866de7246af9f02a31126d29c4b17e1686934a913c38cd7e759bede81ca1b56b0852d9775d32e6b7db78cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa4cc754d9d406d7be2755f3a0e2383886f1a4e345343eeff7a266bf91c36a266cf64c5d4cf81a93681f57e6e0eb5712497b0309e2f2278c84862248ee58419adc313bcb39d758e33b65da2dbb0b1e1f9e4aa2f2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebe55f135cc6da9964873f4f627447c5fcf59de3579cc63bccb866cc831f9d81cd2711ad3d262adbb1c274942a0ffaaee4cc3768518c0d585922c80fb72d80164b6da56060d81b8c03e7e7e1269c73f71c5450d06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0913f2775613c9932edf30155b81eca0d293b01df71f7f2c43e113da57beae6a19b3120e510ae0ee20eba9f9b4fd06a4efb347f92f41b02a4a16928c682b25af779fe6b6d57076d2a1c0d9d572dccd51f3220029;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h531363c6868a54066453eef1bebd272bb5148ea28eff44760b84b185253592e9daba8e8b5ea9fbbc3f9e7f62c5dc3b8aee0dc6ca9ac0b4369a3069d3230385a8417f7f08553ea074c5b244f610a4230edf5dccd29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h537a6e9c6eafcc603f4af797ecb3758ac05e8c6e87dcfa52522dd718581686b169297f934b16b2abed00d00cd1cf4a4207ce0aa7337216dffcd28a4a36ddbb304481411af766d7b923b7cd6d94634eb30cc9999b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1904352410e65e28f0b6f90db4aff0d5b028801e392eed43c7913f9fe009451ee78c4c1dc23ebe8af9ea274a5e60384299dd74c289bc66e763642ced80a5e3c80594b8429514881d9b2eac9bbbfc2ea0cf0fbab7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c4defdf3638bdccaf0bb0f3e90b57d994f3cc27b0e381e032f8784043868e50bda7e2a91883b7c327f0f9188410b26146e9614c5f441790244439142c653b675709a3d70371871df5cd4ffd118fe0d2cb2198337;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77166afc987a783a439038d213528e9fe66590d65ca6ceac29142d0a37b234edee396b8201d2090249846100bf49f92dd56ff1ce3b02920be910b4bd38b1b4dcb76c749d99eb146c7cf4cd94ff0d3d7c0f42c25f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha066a25d54beb43c1bee8c3d5dd4dd5967417ac3e2d0846a20198b82e06caa8ed9d4ad0c3d8f2dd3a259829d32c80d30c11db1d267a15b58e2799ab1655f1c4f25ab2c89c20244398420c290a2e6e192649ca9655;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h620c54c398c72ab68c4536d2374c4e25d64562fe99ca640ba8a88d1e493db2e4b749f1c6d3138a3c37a6210188eb0e32d6a81a61bdfd95f1bde5cb76456fc65ee7c3521104ccacf66133111e5cbbfcf6844d5b0f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d8044a49d2d0efb4bac4e98d3c0bb126a2a9fbd96c3b2b98d8ee8f8be7fee96f07ab6201045df50aef745a37a385bd8e2f75b75c3a1f48b78caa4bc4bd1a9f78c13c6e90ae767bdd3ba6b1baa2d48f2f46839bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he216f20b4cf07c1d0173ed56a32747f3937716628b3d1b0684c711744aa20052dfb868efcb9229cff735796f32165ef042a64ff0a80a4b7683d919eb7ab59cda4e9a1e6c216441c7588b0d446beb526be7c8b4737;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcd45da9a7febb2783c971ebcb77393ab9289fb7a7edac2e2a8b3df3ebe3e19e4dfb66d2b065375e3a067203c193a27bfa141beb955c54c40e472694e8b1716c243d1d74c10d0588573ff6dfd84f4b28d8ccf1b4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7afac23c78e2b07c7819127670e9ae9385fd105bd336e976b22376085b76a63e7ec7705d6e2cb1085ae899792ebe9e36b790d3b080888fcd3ffb57e97b436988974a42a937accfd01f692f6a63eef6d49b240bf1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba205bf57624190d14f286565a9feab9f637aeb5f27a052d534542060c544b11fa0da3ccf85411a752629ee8d9b7a982a6f3cedd131e94b5d37e5b7a48a72df8b8a4f587a0836757077b4a73429f0eff8eed84dac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbd1696e0025c0b0f8ca361db663473b04c99215684f44d3a416e58cd9e859b166c3a7e819bcbb0eac3ef31a41b0a1de378915823f26c80db8f3093f583ff8214ddd36b06ecd69692c4122086a8022a45ef557259;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e52bd4ea642c44c3feebb70eac9c1f69a2cedead5a83bb4955b0347f17bc8c0b6e79e453bf4052c394a0a0ab74af11fd8dd400b13d32e9bd2c1f039786158a5a7634a8da051be256907d6b5382f8c6343c0ea304;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d728946599c668285b0d1184c9cd533a5e3add909eadfdc94e5c423b84dfcd863c89e83dbb5f587bbe7dc08c9b1b01744525bacea459cea879c8446529fe63460e8071e577f23b1c877900082e59bcf17111f07b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea9c53e5ca35a5b220f53392c1a793febb8f44de4f8b4799b455d4dd4a87090acbbf76d0b6b963754eb846063f702fa5c85058e523b3046f27f4feee99ab34999ef82403a68f35e5a035094361a1880b6ecdc6e15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha97374a493e8f1a3ebb2c22d1d5c37f9af0b2f3f517358e628932f48f88130748a73585e52bbfb81c481eef7eddd0bec6b9289c2e14156536a215acba83058176f94b81230701dcc3687eaac015aef4e1a2f8412c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h909c33717c2c6f7182760aa06221edffa46dd40fbbe687933b6aead587faca9f298dce4f674e9cd233cafe94ab3e4a599e06de2b7934b489b854bfd931a90a19091e086659d7a2ea7a7372eb47c12dc9cbdff0951;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd932c6188568c3f7a82bd739684797e84c34bac452b538cef290fb7687b5fe28b4740b6f9877a308fd87f320e7a902f56f80fd52e366766e0c3c94b324e132af28e946840fef15f1097d880ac86fe5df5af9b1073;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafd4853271253ab1463c026f5a2d9752a1a5a560f40fe7a5c657ef159f3e1cf610df3024dab18f335a58f29483d84894417dceaa54f54d4390f40cf308497c73554696f5cfd2df895344e0e7d24392c969ff229ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ac8948d59c6ba5b066458eb03837ab05089d20e4a9010c4b9b8a6aa91ec447d6b011bec6281994ed696b7ece343c4623399fb1a5bd1b436771d95d44a8cbdd7fa96e9cda229d1d1935e08609b34d1cdf667c6839;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82eaa069486bac30e03859c0e02fc66fe761f607879e29f2d2514bfa511d322bcbcfbd624e2290c6a5e6cafa8be8f35eb47f6f5bc3153918b7a37a53b0c9795a7cb6f918f0e44733b20451cea1eff37fbe6431e02;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h748f5ae914ad6f98dc4ef459527a59813457027da13a7d00e4b0c7954c87cbda754adba6976763db4327724520521203e3ee6b037fb3074f4fdea9887c4a65180770d9e62e697a0a720e2ca129f8c744ac5340546;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3478c2bcd2dba8b5b7070d2a00ad04f4ee11030c70b6190dfe08a4ade90ed45da0ccc583d5d8fb7f2120960bd3326ce694c53f945791c6391c8185a6aed3f9d25077c74dcb841f3df42cc12f750562a010d681aec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fc6d3d6430c898485db64383e5ae8f7a05aa925c0b221ddf0a289b35b8ef2ba3bb849f41049a7d70aea1a2a6fffa9feaa97bc3bedf6f2392fe515394851fd54bd355676ab2b96fc55c2859bdb7dae6f463e76402;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6d0166d5733e20aba46838f1937b424bd294cc62da44e9b1a3162bdcb760cca26211baafc9967ec6d8ac961d56cd6864a9794997b6882bc7a9c76ca965d7b5db48d40930a965a9e58ccc66f1781acba7f05094fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef20425d7c2c050fdb7f8f1a0e54a8cc21350d9260367991061c455f54137df29f9fd0fb84e47f6a7ed71f4fd8082d5efc33d35112eb152e01a79ecaf57a4eabad7a7b0a6716ec097b550aefe782122bb430bec35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd939fe7fac0d581fdea378e54a48502a495ed2e7d32a233075887ac553896a1fd6a6106afb8568eb4f71a8b25f6bafdd4fa7c61785fb5f507413da642b24cbdadfa96029a1d770629366d057e1f5acee8c5ac8401;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h148fe16a065a95d4c34d0896500096fb300861fc7849a139beb423cb257283c23dc5604acf00f8fddd683a8b653642e3b1ddad06857ed54b5eefd1a5ee8aede9138d692af4ff9cbdd2f122b81dd331fd5e954ab1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba41ed6872632fb2a0394eee56766d6d7f614b7818d358be7f606b797bb6d9f59c0f949a77c8391b40bf06ae77be1b524168f6cd20308a7e691e9274e1ea9f10c12c2ec030935931ffb0b47f7a482a7c949c6ec7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae5028a422a5dfaaeb07ee386e2cb2481dc617bf4e4d35d9b378712a25ce3607af4f1dd86a395c447162e26be217af2e5f55394b00015d283eeccfd5eeb820c6c93a601121fe7bbbe3404e2504d727c5649126cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h309193e6602527aef975ad7b2351ac524def2bb287b1d3b7c57f32c1103e1dc4e8748062f5478803d240fcccb63c8c4aca6b8efb3a3f4e253f85ab5038bdc39b937ebdf72c744ef67845256d56ff23cabc68ef2c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45e6cacbea241e33386f49d287bb528b5b17d690f20ae95719eddc0786ee2d6a53e90e0134ff649416406802fde44eaedc0158154b414f5f11df3007b238e3c22d665f0a8fe7eed5fda2eb7fa1c8f73e95d095ec6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf3eb3927c78089be81064cac467ab944516ac890e3de760f6a0dab441a0a4eaf13298b6e2d534325fd6c669333fd2eaf7c4006abbd05d5f5d5ea56c0bfd148db819c395f33f087c656c520645f2e202889553be5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc65ed3ffc17881f415ee0538e9d7a4e27b38d029733408d2f4306d3b9dacbcf8c1f7c96512a92d6b23a524f463a1194c0ffe755466cce758f915ed6ca2322297b78168e2a17f800f53abadf27121277c5931f54d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d9bb16e281e62def9e004aaf1d66d878286133408a2762053a5fb25bcb672e54b7d0014f2911350e07e9c764101e521cae7c8ab6c9e48f3ce47010cf9562862786f1abb25744895b6c05554bad6b17f9598c38df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47c7559b698383fbc9eda536055068814510982862cbebdc1d8003c003cf363ef05e477f754780d3a1bb7630ff30913f7d3655b4ece380724c0d53e971ae323a6c605b320045bb671fe5afd2989cc701a233fcea6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd135d375f4c33aed32a55687dfcd623bc78990e614a2a48d5a30d0c627e14c375cb6d3e0e58e35a9955489edaf7300061b17139024f54b5ddd8fe8acfa10a5c3644f81307b8125312109aa6a19461c33ed3538124;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32ead4b118edc02389501d63b1484d379d6891b33043165122c1b89eab57fb6321c96a7668880beb6993d435b6526f5d70f120717963278df8a48ce9c99aab5caa94d89a7a6a31d82cac5c479db458fe20a466c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed598b69d84f022079ab925aedfb86bd6221f0af9e533e8b4488c470834cee7ec8d3ea06cc18551a57b0b4fad383933d17ddb9459a383360ed591fc381388bdc0f81f05add9a39c3b818622ba775ac50783900457;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7dede54009942e388ded50a1ae03fc214159262d5f5fabc0b4120e7c23d613cab8cc05abe5a6c7f20355cc0c4429f0a27615ab4dda89c8d75424a90203b575ccb225827d5a8f5cdeee0311356dddd6f85d1d45dec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef1abd8fc4bde296ecaa97ad5399f6aed551ba251045a7a044a1c294d86e6a42d5b49ee8ae714f8b44afca9c62953bacd9d1b93eb81d07680e0d5f54184c52975960bed5a992be70032ed0681660b8f1c3a50a8fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed9cfb1242b28f035aa6b8c7f0a8b91eecd22928b27b376a48986f7d3d43319950eb19a236fb26f5b663409b46e8d8f78a4b521c1b45eb79cb2506b443669a174e58735914f8b0562455ff0bea018d66ee41ee52f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4f1b9a30a57c7aae7e5d83b86885507beee49be4b89909b15b105f4b57053345f0ba3f5e2b978f73779f2b965e0df69ac56d5f4fa09c01f88bfd43c56930345868aa4972045cfc1f03eb0bf8a82aa145026d365;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde03d16b6f925ebdfc3ab31a8f652b189eab9d523b618e42075700ee129e9b653a296b82ab98ecc9241591ee60a93c225215b8302016ab9e9313b0e1e351784c91e97695968cfeb28e1be58c125dd7b9def66a2c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9173668367fa57b4cc90af866585a54942049b7b21af8dca486fd80209b29ff79e74f1078c9f7903cf0978abda12f18525fce9243a0debfdc8447a4b590d70690822d19e58595dfe80bc0539ab6ddb133ec299e47;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d6ae9dce4649297405662631b6cbfa4dfdf281b62391e44de90617723c096aa0304935cd3dd8fd7af8f5dc8c9c84d689708d6b8a7b242904d5f8849b1844b730282be5ade1392c9426882623ef8408b93e28b35d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5af84abb48e052516e756ffb3caac2ae47bf9294968c4c04ba45d986d52f9677d1f94285f32df74c63ce71e06006a05ada36f598652b9f78dcb7239fe69d3eb54a5906cf6075adcffd67729313857c0873e2ced4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb33b4ffa8865666d1358f3454a190ee9f91e870db0b2b001813444de5d9b4d39108ff2fc915998ce827a55f8d3cf8bce451aaae342bcb5be943f0935bc4ba96e1f6a6d284bd22d24c047fcc6d836a21ce47b8b4e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h856f16215d7b109e5ae54c77d00828c6988d24ade6e9a8c7a1965903041159331ffaf5ed4298d961e90b582df144d1ae2956779d2b051b2567648f0e6444287fd32a29168562d1b99bf9dc9c5f8b360f1482e5e60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f712ad5de6c9de0cbdb8a3bf4ac8bcae0ddc99486ca80dbb3497b1a3c62910c0f61680a5709a72f700f3f8369cbb32f9e43f9633e4d21a445b13c7f5700e1de935e5f1423d7aed633a36ec32cc05616d0f77ba1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb096f6be7001540f944351544f485aaca117a7ea2deece8f42dbad60e912066b9c1419eee6d7e5ad0dd9de7c1ad08dafb0f82cc1282fc334290bef2fd3ef051a65a422b398950dc447b120fbf499799c8ff1676ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba5277d9780ad42f3dd217e48cf921b0a5f2919e7e94defaee70528fffbf6b3e433ea55dcd31d965675bbeecf49e7734a7a04146f8a3161323eaec8b251a6fbc66070f02210d4d98fa06f6251d8a4d790adeb0fa5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb73701f782774cfbff70ee37b17f8383c05252cb3130f78dcd754fc48de177e3ddd91c1b5d4ac78cb21a22d8eca0140e0ed2edcc4413f976c8e35f5c2f8f446979ccb9abec6989bacbc921136350c43dd4b1830c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe8b88daae56e87876e5a3c08958c838a41d42170cec08388eadeede1958611f704aa81df83cee282a6637ade12f3994d39b420a3888d21d40b6229e2f81bd3dc783d1df926d8e57d4ad0d58a1cc2e32d9fe4b7ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf395da00f16660e5cbb14e6bfc267fb15f953e50606e966c355de8a6b844538fc7907695f83ae971604894bc70f7d0a21e943e829901bda909dc529eb5f9c35be56437152f3c4035fc2ffab0bff9d16957b6ea18;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdf9ace06fbf9c2dd2634b1109da4b7976b6bc9c27376dc9ded0a8cd3b6c18e2c36743c7863f465d8d33cb3c9878d0c0a3828c3fabaceb4611e668812c5706ef5b7eb07538fc425e0294414478aa21817639ffbbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31363565983dd0647bb3e175d3765ff76d8fd6ac635e5940e73d60821f74f87d85d19309ac6a3be29d0e1b84897d320ebc180fe7da8ca13b52653fccea5a211918e4d16259dc9b3ba53466587e364207e6d97df9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6df189d15dc708616e72c52eb5b6c11cf2a5562e3af08f23ad0f461f922f3741fcbc7487c27fb31ace7b154736e5fd84046e3cb8727ba47c617cb71c3399bca7e6516469db40dd6e3f509e0b7886a4ee7c9a9c6f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h504ebb7c0225d72716adab478ad5f7252c81bcb6fa55186557bf86b2b2d4c2828a72dd56319c27783b1f40d165e72c4c1e9c63da873142180cc3196b5eba86cb6ceec08efe632e973272266aa65c67c5e04b6add9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf234ce1bc24625efed23f0903aac415dc104f4a0e7300832bde4f46316e21eff2f6fb3f0a7a065292d6dc608f848443c15f28ee60328b8257193d6d949c1db84f52a8a1adac5b41385a814c7b189dc22f6a56145a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10f2c1069994584369501a614a4232974e62fe3323f0d463d81010cf0ee4e1a294ff26d16a752d0b1cdfe485c2051a572cc14be424946b8f35cdeb0008b4d0ee64fafe8b98a62396d6a19cbc0fc297122ef3603de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5950bbe71be46119e5f89c60df5007ea22ce2ba4a2a52f04fd77f80a7fe2766805e2f0638d1ce91d34f5e3edf1deb051f33feb6fb9c2a7b4e48402faf0d12ae06c4a000aba8e88dc518f193c71122270fdeafafa6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac8156c8640121ef22769b39d7d4dedec712630d67396b568347a86eed9c5f3b0dee17c5baf80afd2f1b7ebda7a861784ff7740bf6b6d19286b847af174ce76b129bb7498b029829b0db49d4e94b55c8bbd85e433;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd86e371263a0cdba3b2f7f2ba80eacbdf172f5c038e10f83deab807e531cad33dffee175edab6140b51a3b73e1ed5e44bb1d73817f4c42a0d74aa05c5747e898d253985d7ac980d46018bf3eaa9df43c3963bce93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h769fedcd2f6650badb24db2b8e97f479668515863f00bfdb54bee30aa7842b58831680bbd4908fa3e575268e3e2ba75a401687443987371f6583a77dd6a511dd84f345bfbea03d57f98f6ac52663d020fffe04f0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29b0cdf0ffb3afc54e555ede13b3f9d96675ae7e6796384674535e045311774a67a3c4af4ca141707bd8f15574bebc7a12a61ff74368c475990653a7cc10147d958bd8a7b882fa5f2d58aac55224e48fe35862fcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e7865121897628ff63f7a790f14553d96284a9f9426147b7b1c17d24c52671288d2a3b7df463b6ff399c32895c3fb64552e4bfd6138314da39fc10d1d4875e70f670e09158ca49a734cb2b8aa848242206a7ce08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h726ba6ff75c5d707e690f02bc80e3f5b91101efb54bb32645592a12290e979a04255e6a358200cd99a66b1b72530cb0c4db4e26e803264f1bf5ffef19cf93fc5605a0e8ca6c88bd93a63f6086385399b5c14f441f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23e7b96b23719dfac16aa566b85ddf0faad5bf61850d9e1e5a458eda3adfa4750737a1ca0efab0dfdfdf0c4dd8d3fca2beb31a9bd7fd70adbaaa3157f0218b254b1d402e3eb011e0d6ef4ccd79724932e6c67c0d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd2bcfecf6220fffbc4bf0bbee941672a6254eda2b6bfc9793387e0e422f3aafe166738caa0e59042dd50f53f875785553bf16ec55c4acc6c50d1fb3bb0ef9fc726fbccb26c45f3f0c4312fc01ec049fce22c65b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba85786dd505a6758bf4ed4ad7dbfc8a95ebdaa6ddaec7d4fa1636780a9db1993b914ad7893ad74c14d32c4e287e57672939a37435460d2795ae3f25edc2adf2260d4a276603f58ec0e2fc7bc2fd561663af03514;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcc4319f8aa572a397a8ccbc5de0ce4b947826ffd4734b82f803c1d52f61a7de48e76a7b2b5aa1cc398d4c54e5277e478698a9b2ed793205bbe2f08001649801d7210e75d5e0ae1d100aec23e8de5ddd52a013ef5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b022c1755347406a1232ae95df13a1dde67a98498807ce0f366ed35a80a47f68b9d54ba8e2c1e2dff863c298a46ab323088ca4cdb42120df33fffaac413c9936b185b5e6ce3248dbeec831dca5129ad57116251b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9914533f6c00dd9d0b96700762c8b8354f8a079a0fc575a7dc93b3d6151b6237662dbdc1f2e11f4009078dbd2befcc8abf8f85314329c8f18056e925fa3eeeaecc30e7012160099881540349590b9d8f122863095;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35c2183fa8863b4570e83bdf92daa043527dbc8de271e8d914bd281afe12073c79c31fb741d94d3b42561c324ad4bc7d4bfef0ae54a4e5afc53e83a350dc1d3f15a80dab69c27a43ec4c3c328ebfd350180fe0ff9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe94d46a8f3b9ff24d94d4bfcca13e5b6ae0b0ccdb6986d18c66c723d9b43f4c74e1fbe1132ea569953b203d807de72762c0f71a1e7738765ac421b25e1d8385a8612585f661608fbcee4a310d50252811c80732e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a0c891ce041dc8800d04dbe70d864c341b9f40e78d5a91ed487c10bbe088fa151887c5b58e3f540290cce3f3b1614ad23b6c5f4e49d63d8c68a153be16f8321facda44d4f1413a6d34bcaf75d791774097ba5842;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab4c91617944e025b29dc6faaffbb5eaacc43de42a9fb0a3ec520233e4c1b75b4df92fc40eb4075d7963e8b6e990f642a734d6cb4f82805391253fc193e703adff99f38af069e547885f504dbd14dc283375a23a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84fa80d546b63af2e3ee3e1d8dfeea218414a4886839c7e8c3647e4ccb37635e8b4ead909caa77841033e0d29dd8dcd684a0f4c1836d91e3f926e3dd3c9aa5f0579fbcd56053f16ca74efb49be54bb81c86888405;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5c3843a2559e3528c2b2902eedf705d147e9e1d0e1b81096721e4b47d932f3cca88fb8bc062e27219a8d7e7dd75ef43bda64259c124dc7794687174430d8e59ea23b3b45b0c3ad996fa46aee5c9523aae309260b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcd009c4a527b479c15b06dcadb987a88945b7adc305f37457f9f84fd9f096d243b77d9b3d3d204303766f19829dc51d16cd9f90853accb5eb40cb308e38dae45760c8f891eee1ed28d8a02469dec4b5bfef49a83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha70426cf5fcdf5bcdfc5dc4f9b79c6e97d96f9ca9ffa8f5547d3ba9089b39864ce35c5c48f5e96ba2e936713656d045d10bb4d9288e4254c88ab987dd7a7db13042e87d2b6e3344831391231952ac42a7b8ec424;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3854d1638d6724240d46668d2c2b33f39816fc4b80a3e563557557d8fddc2ea07bc7f910594053f98eed63172a568c8381773a5d569f34a612896f05e97a998763ccb3e2db3db87ef3299417ecef979124d2363a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccc8fac89d46bc55b31ff1788b906d8908931c2539fdb5e123f5c9dd4b2240a9a6fad1a6a2361ea408e5ff2d9fa39b52780149fbc1aa791cefde7d8b8a48e04b0dc003f98c4bbff71b667f7505e4ee1262e5ad84e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf422fa8be02c7898119f3ce9cdea9cace9ae4ed031fb4f67c644e0f8d69ccda38d8124ba800ae178ec01e1c855e96e5d29d610b503b3ea854af7c8c53877fd4e61c32804477a66fa755356f4549e61db634ffbf35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23344ec0eb065bb33d14092b0d7019a5f4955ab3841bd298ba969fd5d0c4338b56a9d5854204539d9d947fc16af8db8073662aabeff124294c1ec2d5648c26279bc8e917ec17e57c384f1277347fbb7c78c53cfaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4496747250f8e8360237c18f737bed47dd103200e545438e58a7818fa8365f8c10978110fc2d5bde36896de8b0388fdae35b34d379a1593aee5a4237df602baed04668c7e7f5bbc308f8a73edcd701bbe1793d864;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb9b1951b149d417bcabbea4dd0055164d1e7481e32bb35dcbde5beb894deb8ba3074157146c6ce7fab7702185d5608fb2065325974a48b6190feb9a86994a2f875f3e8e4749ad2e9bfd4dd16fdb32ac1c912cccc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb25041067215db2dbaf60cddf2923faa104561250f7f5bfd6f4891fc5b5e186e51e91d3bdabcc8afd7f6dcb9655790b1e8fb1a8bc708b46997ce2ab471627af09a0f56e361c23381b1b5b52927ceb860c34372b77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1fe1f4f3d9af4eb69b3fc4e7b5d5f6ac17914b2102a47cf7d4ca842f44165d578252e228d2fd087560ac78130c886bacb11cd3bc539d5ab7941b0381121124b568bd1893ad911d31618e1b04a6805bcea8124143;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd1d0498e7cf365a98f3a7f8b46f6620abcf9422fe354aadb0cc341c1fb43e3f9174ceb595d721e41ee07fd7fdab0c7e9c94340fd9a70533aa0ef4c30b3d3601f67fe0d5d9bd4741b1f263c41bf76a97711b31c9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dc50a049051c27b3a0b7b49d14d02c4489c0ab531db1ba9308dc5dee5270f5fa4ae10262dca0897255c2a23de725cb457e58c61536416d627daab102093bfb74d99092443c2aa98f9e274b732d69267f453e2a3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee08034a083caee15e08eff1e8b4a48cada56682b058cb8ba86095405e7c0ab26d80d1f65c1520a78ae600ce90cd8ec6307d76d9a61e691f44406d966825c9c8d4bab184cf208cc19430c947d41fb8dbcc5b11f23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70891f66108a20219f645f607a66a92a511c26468a83a1e4514c0c93304e8e6a6d102929c69ce8d9ab42698ee63a93f67021d68b09d5bef99fac66949a7ff33772eccc6af4a2e2d7c495c482a14a7f9bdb9020747;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddfdb767cdc2175daa97b5d8edbf0e1b2c2505e1da1afd0f39f58d941769bc6f96dc11ac49976310252ee1903d5b820cc5a06637832e586efc7f6ef56f768e98b4a00bbc45133203095bcd054f1ed502a282f654e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha42a8c7b7bc363ab368ba56ea8a75902133c65f625a82ad1321e6ef684744714000fcd2c3e913a9f15d20a7a8d2573d254211ca414179e56f67764b05038ba1291144f498a1bd7d948bfaa9860f5cb49921a2a54c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dea324c8f08de5aed9e57c51d96ca5533f5268d3f1e0e4bb2a6f6753a5d3ddea70d822143aab3ab8a6da9371be42cd26a2bc89da6b27c91dc28e8d4e6fc54d500ec303eb1cce53fbd331cf0da356b32f64f5aae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h449cd18d355c637747802f981ac2e741a0996ead6d3682eb56f16f716dc0dc93a69229f3e4b0bdf459eaa2899ed2a8cc8cb552ff88682733d6547adaeadce971d1776a807c24ff8c2797463018eb7c16ed66a9b35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h849e420e1badc92aa175f52b09cf56dc16034c6fcd843d791d8fa75799d826df6af1bcb4affe84f9b642fbeb2f58b15e178452cb3545e8bf7ea7ab760ec2d6e1ab66e3727610c99205fd0d47a4190936bf3584800;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1067fd28de26c2702ec680fb3b6cf4ed9d74def7274fca1184b82e64cc05c06571d7d18f3149bfb4edf6b2617857f669b4bc8561327a4cf46faaf94ee6b9865bf527adab7d78c42e682e03c9644b274be26b8c7ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88023960f52cd9f2a44a3912bae1a9c867ba4a493bfe9ce1cca1739e987994560863bdaabd9016ae6fca17830a58023a12786c2f6643d393e90957b71b65619fda6a272f83d733dbd2214adfadc365b6621e6605e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bc0ae5f5f4363cd29f68d1323be4e8b46c5564f2de4a5d785b627dd8190245c096bab9bdbb743bc35d5ff08fb94bac8bae477d69ebb74d0bd2beeb54f450cac9304230db1cdecb883096279c4f4b9dde079ebaa0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c95c2768ef0948db54e41078288f0cb1622b485934cad15d4c365dcf83bf947be59b9ae7778af9b7d4369a0e1808a44d16abb23bdf41773f69fed5a9a06dd3e1640bb39f15eeebc38ede0e5d0b3d366835ae2b8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha95f5bf7b6624e84cee442f3dbe17b98d5d3767ab58437e43a2d5d7052034ba1dad205fb7370b8fcf77c83369ea846cfb9f865ca7d2ca2d8c0556560b7d550f3aead3c6286a7e98a5e1e47acc877c6489ecc86502;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha717f25eb22729bf20cd961ebb154c548a1a420ed416981e75de36cb55452e78a8033a953d062def2d80c5f1f8ad8512a4369cdd3f88669e5e0a4c3404e2950c2c54e07c537b96b8427c68aafeaff98fc997673af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3e961fb83cc911ad19cda7eadc06db6f58ad485929c839d51eee230e8c096e3c334b45ba844d3f09495dce1f00b756509228c15390f12f0395b8b8d708422c4d74f19bd457fd3642c9307f750275f9069162cbae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1aa72a626d070de65e254599b2016fd140cd8efbc905729a1ffcdc54d0c47226391f00e0eb66a5974e623024a88d4b3b683a2399219ce9dbb247ebd1adc1b6ac593f09d29c57ed8d55dfd506065b0610a471ee6e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fcce9d69e01028a2d37a16767fe4b3c9d2f544740de22d32cb3f8787aa39b2a44cb790da925aad85ba81576a99e0cea5cde9dc9744fc429bd0689d6943f99862b1be807c808074a2ed6c33a56b48eb74d2b06260;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb239ac03494df7243445f9ffeca2ea40e1170ac44117218571c0e2dbed8bc0d01946fb6006d45ea42765c66e11531ad7a965e619f0dafd02ece6bc2d325a2027c9553af5ce316688679d2fdf01fc1b666df981425;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23f2191aaaf377d9e78847271e5d68e64f06d846ebc06f847120523b09f41a89f894e4bb9660b684ec4e317a4d49513b244f60907b69c9cc6fa79740f908ad09b26b0066d24ec819cff06b2fd9ded0d2c822f4569;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5122c9e5fcefda19998a6d1e5290b5b35bfe90814de23b9160e246e827401e101aad57daacac2c6abaec3fde13c236f2ee7a76de1dbc64bbe6efc8e6a4dd41330fb32d31495c804efc9f98812e2ff829e0b8ea37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5bb2f14fb4d295733f3edcd4afce932cb690d8854234711988a5538e7a5c8fa9f8d533bce3238afb9177cb65b2e328de7d3a53c9bd13137c85c505cd8b93e57a08c99efd6883623b65a3db512b246e0a9736ae5e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c3950d2692e8e44b39539b36bc05092526208e241babd42293fa2bd4d048026d3b3a32fedfa61c73a6ba35a2e49525bff0d05c056f86c34ba66c0b893efb73b24568d3108c5638c68d94a1440f6424b499d489ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb236ac4eca9380078c188b75ea2fdd40adbfd0d347eb5ea4024b974099524aa936d606d319bb8b426b5cfcdbc7afb25d47b50d8752444a19a53cd3d8f12fb7ee2cb3ef30e06242be7db8abde9388a05a11a15470f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedcd4a8435c5eb6a3a7cfb3590bc00a1e94c14941c76b7148b574840086a1ecb17b7285322c4f5ceb70dd872a64db63d221d5282843e0680a95b76e91c32b1beaa0d1b9d18c2dd34672656f422375a946174431e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96699338abb54bf9c0ef3cc6d56c29666360d2081d2da618ba87a9cec609fdf517089908f30e0c365cf260d8c42cca4af08f7297e8aa6514a4b745f72862eaff8e9b79652e5aabbf62b28aa3c423d270ee66eb01c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12914d09560355be6090c98d830caecaf2e07ee1da0464b1c838b7bd8b4fd857e717c1583736fbb86ed3ff92d7b1ae501425ff21dbf325ded54f03b7fa2d5dd498171d2c71eecefd489eaf86b28b40c1d1cf17a70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd92aa08db94d92e6805b2c9c46d0f8034a8dcb8d715e7d41b7441996b74253bbf5d3e65871f221d5a758c801f7f5ec0de90d04ded869bd213406973a58d37ebe592f1e94d31c509e28082bbdbd84bdebd2415baf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ef3b3606ab7c2233762170890044e68cb6bb24b844b735c33b7ec757ba961d249ec9792e6c9f29b1c63f12c0d142c759b5d6ee4febfbd2459106781eb989311a95b7b5b487ff248fa8afed4af9f27db6c91ea351;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafda118cb60a4b82219ead8e01d98d70f3a7a732aa637e70abed1b7cc07b1decee187706a1549b5d1b0e1e863ceca5d254081261ec13250b8314263695d7aebedaaed53ecf8db4071b65340f4f3b8ec21ba46b674;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd5208657f3901074f7fdad528492bf76600fbde7ab39d5059ed5ead8d5a3c9af3f16c4653f18be4361964d06beac78dba0694452c80025bc19b28c2f51ebd0edc5aa5e1548ea138d41539cf98e5fa830562a3578;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cef9f4def15651946de0821e30e19757a02d6fdb5ba5c6f66e56671ab0c0cbcc54669c2267d8692927f6c31ccca81ce608bca9c31b32fe9edebba363c09c778883d1a274ce3a41048f43d396af90b0dff8b5ef1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfe0622c4fa097c921dc926744a9c453ec2da77cd1cb0392cda884820dc040c32190218d6cdc2b9464121398288b3dd44ddbad046cc21430fe87e4f6197b69b4e34e883a584cbb198af997a8c9875a8a47e1e5abf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20268a96e83470dda38803d6e0b553cb5b4f19681ad3ac7c681419e6dbcdb379a74f15b644ade2958848bfe99e84d2de334bf74105b4ec1d74af0c546ddaec87c4664762dfae4fe4ff9ee38e47b369c2de4ec11e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f465326d78c790bed4b3a53fd1ec4bbc33e52c940770c5286fa23c497f9dcf80c5e19ecde6ca9f421454e39febb94f9be35acab8398442c4b5dc305fbaeecf7fd98db6887d69fdb3b6e1f135caa46d2090caa0d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea75b4c38420c23cea543acb9de86093871cc09ef7baa25bde8f5bb0be9ae97f7ba87350cddf837e8883db73d3412cf396a1d7e7cede7754a3b0dafec3ea0131ad7a12d49ce0e351dcdb8aaa8a38d92ce12974aa1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8105862ffa516e8052c2ba7cb197dad2dcf8d37c067e51bd0e19d0b2a0b1e6b2d5f6c3e59690133f76f1cbe1425d16f6199d847c7fdf123fd76ace3ca9310e7aaa6ff98f9adb58e0de0b0af2d2aa8dc69ac3eacaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7df93dce7bb24b637aa1e78b0a5f1e2b2c454ce35f021d1a7a1199aacf044c672578aa8989d77a72f49f7275aa22ccda590de6a7578cfe6d86e0fbea8c6432a05a26e18d5ace93ea20a7e8b44144da783a38ced12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83da5f8274f787ef56a7bac6d1c2cb578729a1e104bde097d62f855785061eb3566a132911ed6554c3e5dad55b6e247deadb0ac873b0856daa2c4101fccf72ff8b3b66589f0676d2fd9fb6d94d623231c9531ac0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ca51d19e3251a055cc9139f9e2fdeadba4069941367541aa66e40199ef3def59350444abd38a84a987a71afeb9d6d7bddf9cf826c337a12be8dba818cf32f069a1d24f87c0553828094829ca41fb3956e6e7ff3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54697daef7c9c06fa947d0383a690e53284e53d7def31a44bc1410ca26bba4d6d252c9520411508cf5c6b9a3c37b21836811b8dce8be708aec03f615bf2e0712ab895fe56f118503bdfcd30e0933d24c75a5e6ae8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfacd879c41620d7edfb938e1b669a8b074561f878738ae6a901d2a5cb3fa3d3754dab8080a0274df453d4e51d8ad3a8e01e3bb3077ee94cdf2f3af987c31f82ace54e58984349de211e966c2c4345ad768c839e49;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf37b9df7b2947745b9f32f56da50dedd433edb8ae1f5c2fee457b154ad085eb13eccd13d05f21995350e81bb204f86a985ef325e317dd9b286f2fd546af769c99318c188d3040f5bdf8b2af7487d365d56c59af40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a795640d3d80607a435428e2de2844af37823f3b4032ad3b81ead5a636d5ccd8a5d130b4320239fb05f245e15f5fd97f6b278872b8dc0b30ae3906d8adf326ff46bc2558021c904522734bfac118c0162091aeb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43fffa23b94d59c14972908ac033e154204a7f98049569d483c2710e64547516eaa991a15bb750d99c6fc1f99b60ab63eca7944250110d3b12cb07777b34c89607085635c5be62556fc0492a9c3402e3568199d07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h902f553f89285e69bd1401ae3b7760ccc7f7468639ebe8ccd664e9c6585e17cde3bc09019f06e9b0bebb09b31871c3cb057120588dcf782a7bb57cde2f9481342bb3059a1b1a998df21e0f5558bc894af0c473313;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb24c9e12b463d9de8fe119c6253c50161e06a068ea65e054a0f70e14129a1569149f0b52547170d2f29f4a3911eadac7d355a8bd4775a380cee4911ceb0d14e52fa956ec6433838af0a57f8e8392042f434b6eaf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf00a88db298f5dbb88d360766a6a2276dc79fd341b6fcae7cde6b160205f7f829b13322cac9a0ab9647b2ca1d28d00019b2625ceb45c64a7a361e09419a6171573e0866f9b29f4a16b1cc367f8793d07f1d00494e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72c503cf6d896de6cd5fb19f96c794c45a0077b9703204a5d39aed8f9119e74331a46cf23d9f6cf61b14116fea9dcf9cbd7405be4dc0a4f6122f7dc198416929092b37b16bc54044be4f8c322eb8377a3e5d02d17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf821328ae9f5ebbaa02330521ec6cd61ef720b0b6b9776c96fe00dc69d3ebc9f61ea2386861ff437181f6e636c54e519478734893718c34f8c415e064ebce0b1b39563dbe49c6b36494e97613e4be58ffdcdece4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3b6510e0e48e5e161f2640ac37c64dcd5fbe262bbe8a24dba9fa62a159d915df1590b756e2efe72d54d091d34d68ee4b4efbdee0d16a45b18adc69c8e2fed7f794ab119d8f0ada90834b03273d5826c20d6b3b55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50af3f8b40641d5c5304fe3b407ebafd4fca518b47b9959fff5f2ae3239995b4e16b729f592f85314b1a73d00f71da742f36324768ea4d3391bd1fd892a56f3f727e440df9e261bca028b91036e5b95ba24341a63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cde1c7a617f4a5f86d3f9d65d9b99b3001c0717681e648625a8df0d13ffb3846e0d1d37b123cb3e6b91fc7566a0fe8a5bedeea41b774e68c638a7f8c29df37727abdb7ba4bb91bbdefb168d5137fd1c5926853a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53af51f41e2e8d180ccd1106798dc2997fbb88c92bca18fe6f16694b971b9c1f4a987d619f5db55aabdb907d95c160b6edc19603907c9acdd345fc71cc08be6efe84908f48d195c1fa5e4555b8fadcc22cb8fb6bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9045e98a9d9e8172d909a1c4a62f00fb758dc5d45bad414ab578dafef8c8926d4cf001a71b7b4ec95d3313d6cde8eec9cf0cf63fd9218da7d8f2778033a9413835ff913de6e22bebbecaa0717160b0809c3d29d1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73cefaaac46784e5e36b937a0c5fd59efb6920382d51aca2a266d17e034e3ec03975ce2758d5dd9059e668e31d52010b7b3a251e6df3642aef32e2f6bac23fe3c95afc050c5adda250be513ade5e0e6026303128c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5352619959ee01842cfe8b4b151c1d21e05edfaff911165e9c10969d6593c9f5801b6833400dc521411e05b5765a7f46aa4e06fb4e053f4d5101ce78bf22925f1445b45ea4e2fce6e3b0b8502e6f0b5fb02b82167;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90e021c0319979dd9040c5b1000c7b57f98ee186fa8fcace7abd225e0f2725dc455874fecd55191e193016431b77aa3116336a8fa6ce5593ed8c70390d7efc571174948197e7e9b224e2bc061a1bd2c9df6dde374;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd163fe3f910592f716ece6a37bee544e86dbdf6213c8c4938daaebd34902c59174ec0bdc87a42db3a234830afee3f085ce2fc3919733745f46fa86fe1243edcb63b76fa9903b93c1ef21137ca0e390933e7f87424;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd38f89953ae9f2b04a9120b2b2fd8914a16690f7864d515ae17d1903e5dd8da04078addea3a29871409018c7f604ae1766f409ece5929899aad9460992c12b90fbda6d850f09db43c3782ace34b93b9873980f846;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7528578451a7455a65f79f867255bbe6d3eba0a8f7575028775a35cb17538040320561671deea107ffe28519a8ef50c3d4963db100fa07f2dd90822736723a926be361adb4721400e4af9cddffbe8c27171327a0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hceecb5ccaa195842db15d69a48d485ff57ed14b0e888e3bb23320431010b3bc3cfd90a1b51258da763231371f66f69552df9c689170b2beb2076897491f5dcbe903d6d2922a26965b31e6bedfc43a9cd5403b89db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h281011cc73e21a8ca2f62bab5a34f2c579512fb73e91073cc272b34fcddc06a3baf2d1cf13959185d82b060fc52ee39be7fb02b5f045a4afa8bfb5c50fa4803dd2ff62fc3f6d0883bf4a24b0d887f11d1a25d6a27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb7e62e98dba50063b0ef2e70d0c5aa04ed424b844432aac8ef07e742f5abc8f1fb8cedd90c11329eedc47684e5a60d6c23aec520d487c799aefa7cbd551cc1cb69f6ede97d1d02bff64f21c2a2de345bb4c5624;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7a5aaac8f943b4a556f6930f13d4d58d20a15ea128619f5043cf85e61caa4d1089e2f39788f969e5d626b646852abbd0ff9d02e6ac010aabb68761bba067ad1ee9b0556f8bd0c4f32795bdd9a2ccdcff80bc9377;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e9d1ceeea95f43e86235c282ab0adc8619538136ae03642afa281317c6e3814f7539934aaba4e2862f405bcada564cc62686a7c54aa49dcdac11a8d2c01d75f7868b4d04ddf340df2d4dff42da25593fa8bdd150;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafc34664b26dbe1272ede5a26d3a1439fe01fd11f6e76b074539953f523a54c3b76f21fa75d733919ca8fcd65c3632f4515ef5a575aee5e3c6de89e204268fc00b3c1c7803e7b7bcb2cdd5678af0ff9bdc08a3fd9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haadf4b6167b815a027327176c347e9d1090f25723f921e9baba85e77eb69e71b296c74ea377fc01dfb2ab326541a6eef26955e0d7c6a0b2e22115c5ae5c979234d117cb4bf413d6807e48c3b448a7572c680501e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c1f02f2e652fce6ae6f6fc42690d628a1c3205cc643f05fc8a26ce33e97b199e57c147b5aaf18df339f90f45c2f0c3534725f9bc7069336c4fce64d45619b1a6511302478b5f0e8c4f24216f0cec4d0f446e3228;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9757631f74fdf96a2ef741a1bb57694dac1a30504bf132bee2a6812c65ca1206720b9ea44482f35b9b2c92a7fef2dc73906a35d23ef2881dac7a44e1393cefec1f6ba7646bb6a48105255f95198459e7ffcfb8467;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h695a032d2aa9516d6967d4eb25e9ba0369c30f654e502002e549096bea2567ccb44d0d0e56423e2bf38410060a2bd83d20b367267066e27fb5b6ca6f3a0fc9ee70dd6e0638fb5b02c2b45b994b74e616bc8aa8e7f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea10f015c99a0f4fa55f0abbc51526f90f9a39316c4721cbfce3cb570770e108ebb9e47f1dddae34f5a77290e51d44df05d694029fc981ef1fb9396fd88abafebc7f69fd945c4a9020fd8f22267ca948da36d604c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4760a6f43b96bbf1aea4d8fb4225b069d175d6146a745ea8e0d5b4a7725791e86133c311256d7bc6eb678a8907e110c67dbb27f8f520fcd74aa9423e7fe5ffba74f455a51e426fa525ecd53460c53fef978eb25ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35f64301cf549fee78642162a5255bea439ae376de29c09c93ae18f4888a3925d48c8cb08faf6f31a4880538bc40d44d24451e993110c43029ba676bf513fd88f08e5549740c997f74f85d7e2d1494cb442b498e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aa33c09905bc4848d39a10f631a307998790f35045e8270554f39d67fde375ae34e3c73e575c40cc6a99cc8bc7096de304ab8e03718f94bc184de0518b0d7db175a0db7a69387badb3214229b072e7066fe50079;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb21843614ec70d6bdc2655a4ff0dd2af80f46ac8ad4954992441df46e4f4af8510b479297e917723f525bdf24d57a87597161fed4321ff92e72c1385bde17945da4a1e920badeb4ed9e2f2951c4f9bbcbd2481e9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f2bfac84eb5e54590253e78b3bcc16c115335c9a45f1106df5017c8b8c3b0d95c2f34a5e0127a3f51aba4c9c68bf9d7409d2759dc221e55418ad339bb6df078fd26a4a7d47769e9f360c04c129a5f4597cf53785;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd81d3a593fcd105e2454e713fa548dbdf2094edaba1eb5b755d5ab5dac949b28092242e426621052f7a0cb9ec4e7764f6e3709fdc8a8615008ca65a10c21ead975708c322bb5e1b8bbbe747c3034f530ee95e3e3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h896874738cd285025c4a874f75cf217a88100b591cc69118f95bb30482d2d98402152035668d6a52b61b79973d777cf82d74647762e1e89d3c7ca310f9ea89f4bd0771d5d38c67f99f368a2e8dae6a3e8a6ecce2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30d4b6d2846a35da271c2f06bccfd864e65fbaf4b4a840c98f822c2d3329942312060464a3198598875b7f47f34ca012b6abc1505b8001b830c8f04d7b787853870a3624774408b4909bfceceec50b8f4177e0b2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11dd51d3e4c5b208f266875f7860a16c1f72e2857b86d14a65881db6c46a74829e9a766d0337db1a55aea23c33193a756440a16cf75d730ac0970d0d1f750f2a482ba8ff396f5e442eac84f3f23b6d159199593d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1c80272446caa1114fb0439cf0e4e3940fbd581248549a8790d3726be7c7ab424684c297a705315c2272b647cf5220adbd5100c8048142b6f49fb35ff6cc4078070bc2eaab1849eb69a4ef95627bb02101d58db2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27edfa04b9308c7bcc755076212d6e4b539a7bbfb984cfadf88ab99ca8c1219408b07de4844ff9a2b35033bf9d8590d87de0ea1e99f025f094b0f41b5104b7a31b27105674f7afe281c6269eea86eea100bc57a97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ce4c4a7ec7b9db0dcb8fe8afa0913202a1167ae420a2bf13023e5ca28ecba6120ccad4bf03f6c8ffc41cd90fd1fb02aee870705841069cbad4f493c54a057cfae683b49c578514eed130dbc2e1c41e493daaf6f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cd2ff6dbfe8272d8a9a886a3668867491a5c1d2beecf8b187e9142307a86b43b5797ced20f62d6238eec22340659681bbba0dcbe0d977527604d9c6cd1bce4e29e3ce61918024a4237b467f8b22485f460bcaac4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb2788a5521407927bd823a10c20e03fb6f357bf16115e380e904a0f0aef515ef554c974efa5853de49d38fca00437ffd50c4b41444b4804d6dd933167d4e03bfeff31c05272996f4cb5d2583fadd45fc178c4d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55af7bb888df0de4c1cdb8867838371ed5bd9eb8f21ba764b853a0ce37667d259eaf28af56c19e83466aa034bbf48fc5eca25376b756addc4fda6aa7bd63ec5c1b45fd0e7eaf97cc6eb04e99db0efe6d57bf5b090;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd432dbe31635a33431da922f61e167d3af54c8b03e5f1424e4ab377102ebb3d2a157534d28e56fde398dd4cb2913866a172f2656e44a8bee9eb303c2ae795e1db9c12cdd023d70ade4baaf09971da998cd447d40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19186a95cdf3a90bfd951d4ba7af18d97cedeea0e83cbb95a0afd3ede7dd577bc6d2dda8a0713d6da3b2077808347e218e0fe95e281bab42ff49d53961c5699fab9c32409a9a445a95ab6ed873e24fddaef64d84e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd96bc950e2c1fd0605034b1fb2460bd00e7b777fe09c99870f29902c95063ed1ce905249fe1eb554255044de307d15d9748b7ec2f4ec5feac29e57ba386e166195438185c0ed3596f1bf9b7b854ab260ca373a9c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e6434b6f4ae03a69d8c78961133315c7bbd1663ac9adc9f02c31b73d83feb684606bdd60a2febfeb2d446ab422ef844b1c51765b9c04c99acbd7ba7098917db34a93c6d746459e7f6a014f48abdc8e72fa00ef69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he36cf8375766b30ed6cd9f0302bb6370fb3b5878b089b9371eca58c352e8051c9303b5ecafcaab48fedc71ec6a12ba2554c9319f2a66bb2bbbdce142615fd6a484ff554582225e339a5b56f1024ca1f52c2f97b20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he30a891b50a05ccf146c8b06786fec0e5f556fc6c8ea5b95f0fd373309c82e21bf62c345ebea48858e1ce75f72157b03502dbfe63c23fc573681f0e540d6c190839f62e69f36f51b44a71bdbf4c64e15018b46da8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1eb2a4ea33b73c2b19dcf8d68535d9bb23434269f525eb607de7a0def2116947f80a4cb80cd415476b4fa999648e2fe157e6a0c359300319f9d260bdd1a2bac2bc8b3705dfad7d9be61f700bdf3d4cf27ef7438;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc34a83b66d1768975be44a2d5b4e531a2999b3dcb626123be8c347723e7bab85a97aacf33a64e17c996f4144ad861903688d53b940f72b3ba1c9bc78d84406e6cf7270a4e49a8a8a24a2d6ca1a148736bf8f716f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h941b71c7b77f4eda46473b344ceccadea582d01d013c0fc69bc43a1b2a0f53efcb0c9075abec4aa7d5c7741351418c1a53bb9e1d0f378e7679d6e395ece7403abb541ba9b62516c7ba429a9d5357029074b9a7d9d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14d973f8c44fd51a644ec6fdee9192a405059a1d7207699901b5a69747d2179c27cbe4e1826b4e3e0797468f553e0b2d30e7fed70f553a40a8181e503a5b9581d9457992d8c7cc7614282bd3d46b7efd22909a051;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81c8dba301d8f6822c9b525995947f38713f6bdcbda1984403ef2a43fb8261f90ad08506433888fceea1c28bed4aa3c6706405df74db71b01ca5413619935b6c01b510df9fa0295cbf54ff358877ba9f6acd2c803;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h866364e1a71fac751684b4874e45cdb4e2eb0e32665b5900d25625e6867611b4a381cb505990e5c404632208c04393639a126590e1dd61e886742c622a57c9c4777992ba86a9f340dc5a8e8527e317aa06a66e4fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed3f5e7c7560a6469df874d6955d43aa99d78d7b3607dd9d662a6949802066988d3bcc9a4e3742f93ad0f19c07272172dedae707effc42ed9d3f496e811927208fcbf8991e6ecc6b16a2faf746783fc6d37792720;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha37f839cd934a7caa4a75679769f4f5ee02dbf10bf87ea17c1a2ad56bdf8fd1641ab1e858c84338a7dced2312323d47d71ece83329d7c1431271f6ceaa1726c95a7d467e813a3f2e230d6df78447329d7cf690fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha50b471ce8938bb37fcf7bbff1c54e48656858c99853c2fee8dade94d419cd123fb4c34ab7248dc4df8a69eca2ba7472733368cb5bd8ef3bbfa9854b1f224f05a2192605f84c9f2b6a9f7f4498663125cf494bd04;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9450b43b977f781599824598aa16228c688d8e2d7b4064b6d909409168df9b070a702e217d15549a785a3f0f3a3ca501d0b31acf8d88ab5dc0978bb34f2dda2c3ce01b9f363be1f48d9b79835ba4dff8f6ac4f014;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9569975d711ac5d22d3213de79c02cc8af5495afc208193fa085bcec03023f72d1e33679ea9299549ee6c78ebf540341abd8d203ab15a4ecb133c572e6be121e721f807646e2117d883854e26ee7f4f6322c666ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd30ede63f934c247ce753ad1ba16c30d75d20fc729165ae4beb4e78007f05b2b04b0d864b6dc076868ab17f7f42f5e198b0e681068a7c4be1a4e7542048549afc2b49a5677db8d43d93b61065210bd6232ba0a73c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86a94cd062cfe3412936f2d773ac990cb3325aef8e3d82eae4cd03c0633f84a56825bdab023bb89dd447a7e40dc5ef42627448b0c13916ae41fc4f47a14fd3f3cb01168b8e35bd3623c703d0908fed9abab81091e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33fb73ceb1a77825257618a1c2c6f3e9bf248820926575399bec877003def18918f432ea9331bdd1c92c1fb12cd16b63b20f31b36302af95ddfb8fe61adc6cc8896a1851e7ee6c7476313cc19646a51feef4f5143;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcc49404c2a43b5406deca0fdf6b3f9a4738ccef626d7862f4b68c968a5de63f53338a92056a44c08c87f36c888cbca56e27d44b04a575ce637a0cdf02573dff55be9a6b98868883d6f2eb6f0e6d08352e664f82e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cbe18f3d787f94eeb2fba103591feb8671f5d73d2758e22dae9812a427aed268ac0791bb0da578387c96d55b8b9e1c0cedf6d49b204f6b7dc8c4fe2c517594f24fc54f1eda27d8340fa66acd5ba75352d89516ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba6265f8e6eb295f63af908ff14f2335d9d40481bfab515b1858126be2d9c710e0df94921fe621bbf8169d73e5fbd324c0aabd7427d72edb38fe6d427d3a045b9540544923fd5ac212bd1df097ca033d48f77a24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d8dc3aa0efa08bdb38a54fca24fa45b1e44db42821c2e50cc1d9bd4ff807e1f6dadc084e85b1cbc0f90cc410f58871f83ea1396049949567bb117a07992130c1da9a0b00b946a0b2d14e8b88a671cbe7d63e7811;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97235e87e86d65d1f2f7d413f48a498141f1ee0501c073a7ecf0c206ed4e35eebc6173a4ef722f8705f2ca38b7cb3606f61360f298156347245f133b8adf855d9698661ff9df242aa248de91aaf2e8e6693ac129b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h124e29bc226b3a049188a83870260bd9b85b92da5d10186dcd6ac86e1b90943de0ee2c94be2b1d17fc43beeacceb57996b10623cf3b6047f55b9fa5a674d0926db0528f202458dc6b0fc5563199f3c5521546e3a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha486d631d2d89e1b4bd68eba20d1843005ae338aaeaaebbd9972c0ae06e41f1dfa37ad9b01e894f611ef95fec2150c10f77464790bc661cd944ee6071a14c9d6f95a60593cfc161772dc628237cb052001b1bcaa7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74adf5633205783a35b559adb5f9179c672dec49fcea2dee86bb1ef4933fe3b5dce9c3ce7addd0a1e9cbd32c753d4af409daefa193ceb90f6f286bd45ccfe51bd46941aa6d6042ab1601448bbd1266e786f815771;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9c37478a48c1ed683e9cb30f9dcef11cb5385fd5c606a7822b1b7ca80edccd3f4543077fce341204ad470314e6a0e5db274171fe4d861c27ff521ae78a1704c5891cc24c05a3c4ac5ba4c05b7daecf988e7db1ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8bbc65d1a5caa2b8ca08db13d9090bcd2179956f47ddf832baa158eaa686280b13e18a2124a2fd9e7760d5fe1d243c58193fa624f639c3298282f444222fdf6991a5fb5c39e67c06b36980d27527d2cf8878d504;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5abef36e7bbff6d67d0d57fd8d19ccc52182e6062626db534e7d75c8d5546a83bc38bf71142c57b57fac880ce775993ffea560007db7686a5430f05fcc5e83655e904f596bfbdc53b1f32f003b07461610486ca37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d4e5227d5c28c77ce10a6aad9126a6aa3f69b45ea8b4de2ac8e5fa557ad85876d3de6344cfcb7e4cddc740a6b9ff9f443a4638c9819a8d17e935ccf763688545ea2c334f78bfa3e8dfd46a8a6cedae6d4ed3d7b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfb3625cd2ac2c4ab8a883d57cc3b856cbeebb197b6817e273df3f20bb8e92f39523395098f6781b36d34899ea7ac7800033711089aa1785acd87127aca9ecc03db380520869a6ec0ff9a04490e23983a0b54aa9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf034e746b7670cdcec979c5dfc1532987e1d7626dab8b31f6ef5eab45cc7cfe05d1f43e3565384e8183ffbb914615b85423b585327ee3162c85201d44dea620dad8f3d26d856726ea1f3bffe730621d20a5631cfb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bb5becae278dcb04ff818761379485a4f246f21ccc7995d3f9a9618dbe00220e7b0dea4c58f933c3fa8a780d4098b31e1c9fadfc7caacb152be01fb4180867652d75fdbc1b998f89ea0c5fa46b8b10800b174d57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heee909b5041293ebc3076feeb837c818621e234210aa4f3fecedd818445fb9cc85a1ab77539d21c4a637f4ac9e3574ee8e86d14ae597fa4dddae86b1281a1d85bad48197813b17b43cfbbd5719bcd620fd7114d27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56166f873b245ad78afe55206038ad811ee37a5079e2d64fc0fdb7ed72f468aa8c319f8f1c6145a247e8617ac496f20e1613598690386af96eb3e37da0f57c3e23433739e5aaed94a8cc1a60784999742f8f17e59;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8e78d8208b6cc5ed9304db48cf33407a47098fb80d05342db2966136570ef5b6852617756dfb154e9c157a9a2584e011941ce8dee17554636947c7b4cdee69da59561bf5742a38671ae44f7983cd87d5558d3788;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha32a8060ac79fa74155f2efcb18bd0dfa8f700583dabc027bd36931f9da84cb66e9963f8c3fe939fd31d520c0ea5991771e29e50e90cc0024ddad484584478ad5c86ec3bab894c8428fd91c96654e7d596979c95c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd0bfdbe7eee2372a5304f9db78b6996cfbf79ea5226e0effbfbd28e29a4643a769b6c2bb0b3a1b756a0f01d31c5cddd31b93d1357d34e14046e328df5cb31b1bf6f7a1c8c4bca2ea43a2d3267c35f078ab30f333;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf7f4c31aedc918685f2ced01298e7fc8a4b24f8b20d3c1f11506dc6ce2ad89b87c36f6ff2a585dfda42ac074834b16db25d84cd25d7018fe7f286c34f97b164a27bf56cacac6f6f112def3b8ae58e0b343f52fd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h185bd321b746977fa19263d6c862959ac255969153ac63b02371921db6c43685ccbd471e2d442ce0e4e699ad058c001977392de3926b3bc30823227db9c5604a38f4a70368cbf165e4d79d8df1b375e8026d00b0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4c8cde47198f7afab19ed93cca175ce0a484c8d8407510af1e9f2efa8fe77f0bcead0bd2e7b3534983867f3cbe1efb3448d124aa12279d57ce8bf8b1394d92fa709899bd27c433ac56bd23cdec6e25dc1a32413c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ef5d4da910cf3793345f6e912776b6dde99ad98c6b478e85348e4f5d6a0f0009ac2c18ccd7082be0f8c2477e5892a6a0f77f9667ffbfba3b0363b4a824eba2cf84466e8f0a98682b78ec3d20abf2f7c1b6f70fe8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff9c0d0d7cf12847d94740d0c105c13c00a5a1d2a291932a7b3b72202d9ec4bc117b4a5268343a493ca978ea8f5eb842c9aca18da0ab912eeab8e6ef836a6343d7a41212f680c4afa8ca6098c5e2f58089b80f5f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91ba640ed124bd02d66eea165ccb27518267064901b981755f83da565e76e5364dae2477cc13595b7c7244deec3218708357a55c70f6e78b340e7c8fed944331a35feee626e8ed1a38fee719f07484e066f10a19a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a60fb4011aecd65c94dc648dc8c3a21b6b192aa4dca82186bfa90aef49f6f7b7a92da536f29fc9a406682f9ddc9306c0df60c097f08f1a55acb6595174bf77cec64ca940327438b9211ae9fd1dbcc7dcf8981c6b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc25e59a670dceffa535bd20231e3e7ac6ecd858de71d21fb63f2134e9c9248bf8c76bbbfe096a9b171306dad103e923a1fb72642c873319bf1805397d6b903767172f2909202aa5cbec03879bd04e0a56fd550908;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0e736fa307f681a54658df45c33bba1ee3a2bbd41bbe16a145ddcb8a9697a00fa7c1c8930adf8d044c0db0aaf30d3da886353d63ef7913c39a63455194113fee0a00b8b991abbd9b0542e2c9eb0416e4d055a381;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0c150efd2b35808e74f3a231bb9878568c41894c106448645a49ff6c5489430adf9eae9648cbc7560b3975b9f936e23381d8275a887d5b08778bf5f1d6ea0d6cb93e4b95cbe0c74fce15bdbecffeb2788d4b88d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h475657f61bcdad2586180ed1c8ae5c8b495439e5e07ee26740b6d87c217555c50caf474e4a59319f176751edc78903acb8649fdac7b512ec199c17e9eb32042b908d42e393cb3bebb5b4224840ec008bac43237d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha811b78e91b197ae854b6fcf2492f312e559fc3522e5cae26f1d3c91723c86cbf61938434385304090a7ce4446c3a4194a84df401e22b4e317cb347e6a4a2f3ccd2cc07c8ff026e2de5430e8a63970d9f56eccec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8c36c202d58c44d867d3061f44e079f97cb3924d878d14ac5db8374f3a5c735776ae649324921e857f50196d15d947f9e7bad9d31cd840cb93c3f646283ecdb3f23519b781860460a4c966da16d55f1a1e1b0788;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfea0d7aa95b56a2ca0ccae4b3da9d6c6e03294a47f56221c4772b4c488bf00c29933a3bd1b62a464baad988d81b13d841cbe2046716e3d79946b95e4b295662e7de3e485e634389537f9c56437de53795a4ea2f72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8942a38932fd7fc882fac0f409de7ba966b66e643dfb2cce7929cb7255253c0ef245436effe8e3e03f0b01b620a8d6093a91c4938aaf3349df0368e0761ba13b0313e2373394d5d498b8469606d90dd2a2a582362;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h934090f927db4f8a5f1212c24571550970f8f0ba227b626c478934504b035272a432bef7f184f7647fb127e4f3ef11e639103634b5796e0a0780c43becf9f9ace17a26ee29e5f0389b0d0a7f676df987f7935ccb5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h799d2cb06318254c760933e8274f8f0e3bb1c1b8b87f36a1735f10693118770b6e3bea92fc697b2b8b0d4fbb30e26090d0938ec1bc315d1d295820accc70c6667745e0b053150f0c6839dee41860c55e0a78280bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1289f7e62ccc068f39e97dae0ada14ad9af628506c499d212d77022eb3a58c534f78b77aac781efb99bc8418bfd232ce2aa18a641759d67d478875acd0825c3d9dbdc3eb082deeeec140ad48f199800c08a35f08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8955af5f7343bdad8e205e1ae13d4b68bfc7de986a11a65e2910df63cb713e1f59e242faf26a8d219dc6abcc5a2eef054dfffaf5090918153c424a20867e52c4c4405388303d36bcde2303097685f17978b9594fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h741bc66ddd81f1d39fcaff33ed62c0187aa4114afc1e9d44838976189d14c3fc1877e0e029d3e69f44ffc293678c4ec8acf862b1be24864e68fcca16e3e67afffdf6a81a2563d83d7e03e5fae9ab3f20875d5b237;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ae8422cd150981d33b97e0bfe44ad4f12bf7ad8680138fe23dc87879932b2f8641568c458779bcd82af201929c5e0ccef09945fa2a9b25a5ba7687ccc5c2454fd57e531f1afdf885cdd143935ccf726bff1408e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he76046e9cd2dfea0f35ef0076efd73364d6ed59da7fcc77e59c0c5d0d353958c8291909e2ec51f16fae77176d1904ed6a62c04855e8e12642079a80944a81b8a206739282feab5e91b04774eeddba7077bc50d846;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f41f8e2a2bac8abcc10960e8c26c22d0c9afc7b8059e2e3f01a5c1190232a760719f9c27cb336a124c1f3dcfe59ad1b8d7ce0721c2aa287f1432982ad4911b33b40b25d6c9f8033a0ea5a7a8ae9403baa8d7e268;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha18c70ad16ea399c7893d2e514035e0c52499fe7016a95112b84d6c7c73354749c574d1edfa131fb023d5a2e0f3e4175ee22643dce3e4b4119dc770c12433973b97fb734d987f8c992bdf49e12809d005200c5c00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51f8f3ec3bdc6a6399a5bfd389baa7a53b58f17918ae478b93fc8a397d23e30f57a910d719a3779817224772db934ebcc914a30df3b32d3bbd9effd9d99795a68118d0b3b7e6b03fa37bed8d0c1d0f28856287848;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b4d5489c44319049968a39ce5cb4efd87b973b8f7f8937caa24e603a89a8bfe8d10463e34414d9f6908f8b108ee02e82890bb9737311175c048a03e345935d96881d195b5a509d8abbaff94717424d1a9b667b77;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d9e86c88be7b3b22e881da8c2b56ea70287b36e3578ba52b646ca431cf0c772901af80ca235d6ba73ea01897a8b50fc0ae234014096e1d0184c71fe1f4192926c4391aab87c9fcd8dda15ce278746a98bfc835e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1acddcd27ec0803b3d352e765c9def95e13e5fdf548d5e95083f5c1c3e5d0fb5772f9b7a0820b81fc34a1067be78d872129999bc732ee40de3522999cc45833d0dedddf3496846827140057b3f2487ac5cd06bc15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a0f7592c3e5439e17b5bfb91510678ae3fc05a368b9a8902b8de44fba2c9ec11dcbb6956b984a962099d0b6715c211b8c12d6af3605b6cf8accfa61481142e88f1d6ed9e13a99f531a6483fb54510985dc1d466f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dab15bc485c3b8e52d74178f8554a840f10564e15bd6cf0f5f49de30a76f041629817506f3cd7ea79a336e8331183ac125a1128e34b992424fa0f9eeac6057f90ee6577b7cac820354e313d929cc4945eae811d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha049e330e67dca3fc3b7db7abfba49b9959403f2898b0ff7793696f40b4f851293fa3d4811b69e74665211dd63e2216f7bd9bb014ae515657a6eeb20d21b8e97c6982adb6c2a5c3f8a2291c2eef27182a53231aec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebca95f0738cd8d3de3ee8f002cdfb2b9608f5e57ea53ac3895913c7f6df8c8c7530f3eb8d6ece5684b01e7ec2973af9b8b73e4c6402a04783f9307daaf4df83dabcb2bf70d8e0b6ca49c32f044f739ea2367476d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h796acc0a28b7489465c07b0f1e1e44692220d9fed2637aeaffbe65f3bda41935320dc792ae481a01d07fa1ceef9ac033579afa799ef6d587a52d1063967d86c82437a95b46b8f8d1fe0311015b74ba7d614b623de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha02eeb28eee8e25c315cf5b72edd907247694c6a683b435ad95252643ab05ee008a1cd994dc317bd336439236046f11f961e0f85aa3390c2b3e4d3d50bc81bc06656c229c15e45dfd5e45d050bf9360afd75a05f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h356f82829d225a70a5fd4406b746d2d3807a23b4600be13f244db46971c6ce2aeb0ab368af234719e7119e09005e687181cea854c6ce53103d821457178c3d127b58fb6b090f6fb62e6c18b7313468dbfd9967d6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h402bfc8b819bb9fa9ec97246d87fd2845a28b910981a68fe612624a611b920c1513fdf9172d0c2ee0e7971598bb8661d51c6032e09dabae6fbc37eb1f6e75066852808e4dc4089e94bd374e891a9ea17b01575497;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h592aa5b2ca166df776781487a326021de04eb75d495ee49d469c62803417b50994f9a44663daa359b30080300a66534465deaab4135993b01d694bbc013b3f455de8380fdd58d4f5d58bba85828a044c68ca7d1a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47079ce48630278b3603b47dea8bb9315c6f2d5d711100bb0bab5cd9eee81c63f0261c4a97c7be8724d8ee8f1a89a450bf49b2614b1e4315f3592c59c582266a9c18fdc1c2bb140c3b4a958e8af368c861d6b355b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ffbfc4e7b5c6eb7b76236b546620b98cb86c8afa2f7157e54a932be5768227e37d2863c6aed0b6823449447d33646c0caeabfeba95e028124e7c6c6b07aa8e0cf251dd22643b2bd9496bac5613f9ffb236551e08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1532d06e9a92480798422a011fac5c63010ce227c0de8bae9f2db329637b7e9dcfd17605b2ba0ca911daab4329560742bca0fdb3ace695a956c9d1e976352bd322a8a6912c7ec69f859311fa73096c022f5fe7248;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6136a3edbb7e92e012ecd8b6c4b5939837aa7470de6441661e59bdd9be9550f75f5858e2228d91b2f92f66396541ad1314a0981705c1d5c7be6a2c51d637af288c80e6e950d3decd6bc2ffe2c8042243dbb78d0ea;
        #1
        $finish();
    end
endmodule
