module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    compressor_CLA162_16 compressor_CLA162_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA162_16(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [0:0] dst22);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [32:0] stage1_0;
   wire [47:0] stage1_1;
   wire [63:0] stage1_2;
   wire [91:0] stage1_3;
   wire [74:0] stage1_4;
   wire [70:0] stage1_5;
   wire [59:0] stage1_6;
   wire [53:0] stage1_7;
   wire [89:0] stage1_8;
   wire [82:0] stage1_9;
   wire [60:0] stage1_10;
   wire [57:0] stage1_11;
   wire [72:0] stage1_12;
   wire [77:0] stage1_13;
   wire [77:0] stage1_14;
   wire [53:0] stage1_15;
   wire [48:0] stage1_16;
   wire [27:0] stage1_17;
   wire [10:0] stage2_0;
   wire [29:0] stage2_1;
   wire [15:0] stage2_2;
   wire [36:0] stage2_3;
   wire [29:0] stage2_4;
   wire [29:0] stage2_5;
   wire [29:0] stage2_6;
   wire [38:0] stage2_7;
   wire [29:0] stage2_8;
   wire [51:0] stage2_9;
   wire [25:0] stage2_10;
   wire [28:0] stage2_11;
   wire [33:0] stage2_12;
   wire [26:0] stage2_13;
   wire [29:0] stage2_14;
   wire [50:0] stage2_15;
   wire [17:0] stage2_16;
   wire [34:0] stage2_17;
   wire [8:0] stage2_18;
   wire [0:0] stage2_19;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [18:0] stage3_2;
   wire [13:0] stage3_3;
   wire [14:0] stage3_4;
   wire [11:0] stage3_5;
   wire [10:0] stage3_6;
   wire [13:0] stage3_7;
   wire [16:0] stage3_8;
   wire [19:0] stage3_9;
   wire [14:0] stage3_10;
   wire [12:0] stage3_11;
   wire [15:0] stage3_12;
   wire [15:0] stage3_13;
   wire [9:0] stage3_14;
   wire [17:0] stage3_15;
   wire [14:0] stage3_16;
   wire [10:0] stage3_17;
   wire [10:0] stage3_18;
   wire [7:0] stage3_19;
   wire [0:0] stage3_20;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [10:0] stage4_2;
   wire [5:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [6:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [6:0] stage4_9;
   wire [9:0] stage4_10;
   wire [11:0] stage4_11;
   wire [6:0] stage4_12;
   wire [5:0] stage4_13;
   wire [7:0] stage4_14;
   wire [5:0] stage4_15;
   wire [5:0] stage4_16;
   wire [9:0] stage4_17;
   wire [3:0] stage4_18;
   wire [4:0] stage4_19;
   wire [3:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [4:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [2:0] stage5_8;
   wire [4:0] stage5_9;
   wire [3:0] stage5_10;
   wire [3:0] stage5_11;
   wire [5:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [2:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [5:0] stage5_18;
   wire [5:0] stage5_19;
   wire [3:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[8]},
      {stage0_3[16]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[9]},
      {stage0_3[17]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[10]},
      {stage0_3[18]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[11]},
      {stage0_3[19]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[12]},
      {stage0_3[20]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[13]},
      {stage0_3[21]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27]},
      {stage1_5[0],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[1],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[2],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[3],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[4],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[5],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[6],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[7],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[8],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[9],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[10],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[11],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[12],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[13],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[14],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[15],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[16],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[17],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc606_5 gpc49 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[18],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc606_5 gpc50 (
      {stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[19],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc606_5 gpc51 (
      {stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[20],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc606_5 gpc52 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[21],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc606_5 gpc53 (
      {stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[22],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[6],stage1_5[23],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[7],stage1_5[24],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[8],stage1_5[25],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[9],stage1_5[26],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[10],stage1_5[27],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[11],stage1_5[28],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[12],stage1_5[29],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[13],stage1_5[30],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[14],stage1_5[31],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[15],stage1_5[32],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[16],stage1_5[33],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[17],stage1_5[34],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[18],stage1_5[35],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[19],stage1_5[36],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[20],stage1_5[37],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[21],stage1_5[38],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[22],stage1_5[39],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[23],stage1_5[40],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[24],stage1_5[41],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[25],stage1_5[42],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[20],stage1_6[26],stage1_5[43],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[21],stage1_7[21],stage1_6[27],stage1_5[44]}
   );
   gpc606_5 gpc76 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[22],stage1_7[22],stage1_6[28],stage1_5[45]}
   );
   gpc606_5 gpc77 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[23],stage1_7[23],stage1_6[29],stage1_5[46]}
   );
   gpc606_5 gpc78 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[24],stage1_7[24],stage1_6[30],stage1_5[47]}
   );
   gpc606_5 gpc79 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[25],stage1_7[25],stage1_6[31],stage1_5[48]}
   );
   gpc606_5 gpc80 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[26],stage1_7[26],stage1_6[32],stage1_5[49]}
   );
   gpc606_5 gpc81 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[27],stage1_7[27],stage1_6[33],stage1_5[50]}
   );
   gpc606_5 gpc82 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[28],stage1_7[28],stage1_6[34],stage1_5[51]}
   );
   gpc606_5 gpc83 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[29],stage1_7[29],stage1_6[35],stage1_5[52]}
   );
   gpc606_5 gpc84 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[30],stage1_7[30],stage1_6[36],stage1_5[53]}
   );
   gpc606_5 gpc85 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[31],stage1_7[31],stage1_6[37],stage1_5[54]}
   );
   gpc606_5 gpc86 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[32],stage1_7[32],stage1_6[38],stage1_5[55]}
   );
   gpc606_5 gpc87 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[33],stage1_7[33],stage1_6[39],stage1_5[56]}
   );
   gpc606_5 gpc88 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[34],stage1_7[34],stage1_6[40],stage1_5[57]}
   );
   gpc606_5 gpc89 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[35],stage1_7[35],stage1_6[41],stage1_5[58]}
   );
   gpc606_5 gpc90 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[36],stage1_7[36],stage1_6[42],stage1_5[59]}
   );
   gpc606_5 gpc91 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[37],stage1_7[37],stage1_6[43],stage1_5[60]}
   );
   gpc606_5 gpc92 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[38],stage1_7[38],stage1_6[44],stage1_5[61]}
   );
   gpc606_5 gpc93 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[39],stage1_7[39],stage1_6[45],stage1_5[62]}
   );
   gpc606_5 gpc94 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[40],stage1_7[40],stage1_6[46],stage1_5[63]}
   );
   gpc606_5 gpc95 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[41],stage1_7[41],stage1_6[47],stage1_5[64]}
   );
   gpc606_5 gpc96 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[42],stage1_7[42],stage1_6[48],stage1_5[65]}
   );
   gpc606_5 gpc97 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[43],stage1_7[43],stage1_6[49],stage1_5[66]}
   );
   gpc606_5 gpc98 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[44],stage1_7[44],stage1_6[50],stage1_5[67]}
   );
   gpc606_5 gpc99 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[45],stage1_7[45],stage1_6[51],stage1_5[68]}
   );
   gpc606_5 gpc100 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[46],stage1_7[46],stage1_6[52],stage1_5[69]}
   );
   gpc606_5 gpc101 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[47],stage1_7[47],stage1_6[53],stage1_5[70]}
   );
   gpc606_5 gpc102 (
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[48],stage1_7[48],stage1_6[54]}
   );
   gpc606_5 gpc103 (
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[49],stage1_7[49],stage1_6[55]}
   );
   gpc606_5 gpc104 (
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[50],stage1_7[50],stage1_6[56]}
   );
   gpc606_5 gpc105 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[51],stage1_7[51],stage1_6[57]}
   );
   gpc606_5 gpc106 (
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[52],stage1_7[52],stage1_6[58]}
   );
   gpc606_5 gpc107 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[53],stage1_7[53],stage1_6[59]}
   );
   gpc606_5 gpc108 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[6],stage1_9[33],stage1_8[54]}
   );
   gpc606_5 gpc109 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[7],stage1_9[34],stage1_8[55]}
   );
   gpc606_5 gpc110 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[8],stage1_9[35],stage1_8[56]}
   );
   gpc606_5 gpc111 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[9],stage1_9[36],stage1_8[57]}
   );
   gpc606_5 gpc112 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[10],stage1_9[37],stage1_8[58]}
   );
   gpc606_5 gpc113 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[11],stage1_9[38],stage1_8[59]}
   );
   gpc615_5 gpc114 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_9[0]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[12],stage1_9[39],stage1_8[60]}
   );
   gpc615_5 gpc115 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_9[1]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[13],stage1_9[40],stage1_8[61]}
   );
   gpc615_5 gpc116 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86]},
      {stage0_9[2]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[14],stage1_9[41],stage1_8[62]}
   );
   gpc615_5 gpc117 (
      {stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_9[3]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[15],stage1_9[42],stage1_8[63]}
   );
   gpc615_5 gpc118 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_9[4]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[16],stage1_9[43],stage1_8[64]}
   );
   gpc615_5 gpc119 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_9[5]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[17],stage1_9[44],stage1_8[65]}
   );
   gpc615_5 gpc120 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_9[6]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[18],stage1_9[45],stage1_8[66]}
   );
   gpc615_5 gpc121 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_9[7]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[19],stage1_9[46],stage1_8[67]}
   );
   gpc615_5 gpc122 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_9[8]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[20],stage1_9[47],stage1_8[68]}
   );
   gpc615_5 gpc123 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_9[9]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[21],stage1_9[48],stage1_8[69]}
   );
   gpc615_5 gpc124 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_9[10]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[22],stage1_9[49],stage1_8[70]}
   );
   gpc615_5 gpc125 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_9[11]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[23],stage1_9[50],stage1_8[71]}
   );
   gpc615_5 gpc126 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_9[12]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[24],stage1_9[51],stage1_8[72]}
   );
   gpc615_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_9[13]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[25],stage1_9[52],stage1_8[73]}
   );
   gpc615_5 gpc128 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_9[14]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[26],stage1_9[53],stage1_8[74]}
   );
   gpc606_5 gpc129 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[27],stage1_9[54]}
   );
   gpc606_5 gpc130 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[28],stage1_9[55]}
   );
   gpc606_5 gpc131 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[29],stage1_9[56]}
   );
   gpc606_5 gpc132 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[30],stage1_9[57]}
   );
   gpc606_5 gpc133 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[31],stage1_9[58]}
   );
   gpc606_5 gpc134 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[32],stage1_9[59]}
   );
   gpc606_5 gpc135 (
      {stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[33],stage1_9[60]}
   );
   gpc606_5 gpc136 (
      {stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[34],stage1_9[61]}
   );
   gpc606_5 gpc137 (
      {stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[35],stage1_9[62]}
   );
   gpc606_5 gpc138 (
      {stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[36],stage1_9[63]}
   );
   gpc606_5 gpc139 (
      {stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[37],stage1_9[64]}
   );
   gpc606_5 gpc140 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[38],stage1_9[65]}
   );
   gpc606_5 gpc141 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[39],stage1_9[66]}
   );
   gpc606_5 gpc142 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[40],stage1_9[67]}
   );
   gpc606_5 gpc143 (
      {stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[41],stage1_9[68]}
   );
   gpc606_5 gpc144 (
      {stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[42],stage1_9[69]}
   );
   gpc606_5 gpc145 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[43],stage1_9[70]}
   );
   gpc606_5 gpc146 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[44],stage1_9[71]}
   );
   gpc606_5 gpc147 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[45],stage1_9[72]}
   );
   gpc606_5 gpc148 (
      {stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[46],stage1_9[73]}
   );
   gpc606_5 gpc149 (
      {stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[47],stage1_9[74]}
   );
   gpc606_5 gpc150 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[42],stage1_11[42],stage1_10[48],stage1_9[75]}
   );
   gpc615_5 gpc151 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[126]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[43],stage1_11[43],stage1_10[49],stage1_9[76]}
   );
   gpc615_5 gpc152 (
      {stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_10[127]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[44],stage1_11[44],stage1_10[50],stage1_9[77]}
   );
   gpc615_5 gpc153 (
      {stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131], stage0_10[132]},
      {stage0_11[144]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[24],stage1_12[45],stage1_11[45],stage1_10[51]}
   );
   gpc615_5 gpc154 (
      {stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage0_11[145]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[25],stage1_12[46],stage1_11[46],stage1_10[52]}
   );
   gpc615_5 gpc155 (
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142]},
      {stage0_11[146]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[26],stage1_12[47],stage1_11[47],stage1_10[53]}
   );
   gpc615_5 gpc156 (
      {stage0_10[143], stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147]},
      {stage0_11[147]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[27],stage1_12[48],stage1_11[48],stage1_10[54]}
   );
   gpc615_5 gpc157 (
      {stage0_10[148], stage0_10[149], stage0_10[150], stage0_10[151], stage0_10[152]},
      {stage0_11[148]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[28],stage1_12[49],stage1_11[49],stage1_10[55]}
   );
   gpc615_5 gpc158 (
      {stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_11[149]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[29],stage1_12[50],stage1_11[50],stage1_10[56]}
   );
   gpc606_5 gpc159 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[30],stage1_12[51],stage1_11[51]}
   );
   gpc606_5 gpc160 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[7],stage1_13[31],stage1_12[52]}
   );
   gpc606_5 gpc161 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[8],stage1_13[32],stage1_12[53]}
   );
   gpc606_5 gpc162 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[9],stage1_13[33],stage1_12[54]}
   );
   gpc606_5 gpc163 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[10],stage1_13[34],stage1_12[55]}
   );
   gpc606_5 gpc164 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[11],stage1_13[35],stage1_12[56]}
   );
   gpc606_5 gpc165 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[12],stage1_13[36],stage1_12[57]}
   );
   gpc606_5 gpc166 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[13],stage1_13[37],stage1_12[58]}
   );
   gpc606_5 gpc167 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[14],stage1_13[38],stage1_12[59]}
   );
   gpc606_5 gpc168 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[15],stage1_13[39],stage1_12[60]}
   );
   gpc606_5 gpc169 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[10],stage1_14[16],stage1_13[40],stage1_12[61]}
   );
   gpc606_5 gpc170 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[11],stage1_14[17],stage1_13[41],stage1_12[62]}
   );
   gpc606_5 gpc171 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[12],stage1_14[18],stage1_13[42],stage1_12[63]}
   );
   gpc606_5 gpc172 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[13],stage1_14[19],stage1_13[43],stage1_12[64]}
   );
   gpc606_5 gpc173 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[14],stage1_14[20],stage1_13[44],stage1_12[65]}
   );
   gpc606_5 gpc174 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[15],stage1_14[21],stage1_13[45],stage1_12[66]}
   );
   gpc606_5 gpc175 (
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[16],stage1_14[22],stage1_13[46],stage1_12[67]}
   );
   gpc606_5 gpc176 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[17],stage1_14[23],stage1_13[47],stage1_12[68]}
   );
   gpc606_5 gpc177 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[18],stage1_14[24],stage1_13[48],stage1_12[69]}
   );
   gpc606_5 gpc178 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[19],stage1_14[25],stage1_13[49],stage1_12[70]}
   );
   gpc606_5 gpc179 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[20],stage1_14[26],stage1_13[50],stage1_12[71]}
   );
   gpc606_5 gpc180 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[21],stage1_14[27],stage1_13[51],stage1_12[72]}
   );
   gpc606_5 gpc181 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[21],stage1_15[22],stage1_14[28],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[22],stage1_15[23],stage1_14[29],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[23],stage1_15[24],stage1_14[30],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[24],stage1_15[25],stage1_14[31],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[25],stage1_15[26],stage1_14[32],stage1_13[56]}
   );
   gpc606_5 gpc186 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[26],stage1_15[27],stage1_14[33],stage1_13[57]}
   );
   gpc606_5 gpc187 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[27],stage1_15[28],stage1_14[34],stage1_13[58]}
   );
   gpc606_5 gpc188 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[28],stage1_15[29],stage1_14[35],stage1_13[59]}
   );
   gpc606_5 gpc189 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[29],stage1_15[30],stage1_14[36],stage1_13[60]}
   );
   gpc606_5 gpc190 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[30],stage1_15[31],stage1_14[37],stage1_13[61]}
   );
   gpc606_5 gpc191 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[31],stage1_15[32],stage1_14[38],stage1_13[62]}
   );
   gpc606_5 gpc192 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[32],stage1_15[33],stage1_14[39],stage1_13[63]}
   );
   gpc606_5 gpc193 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[33],stage1_15[34],stage1_14[40],stage1_13[64]}
   );
   gpc606_5 gpc194 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[34],stage1_15[35],stage1_14[41],stage1_13[65]}
   );
   gpc606_5 gpc195 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[35],stage1_15[36],stage1_14[42],stage1_13[66]}
   );
   gpc606_5 gpc196 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[36],stage1_15[37],stage1_14[43],stage1_13[67]}
   );
   gpc606_5 gpc197 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[37],stage1_15[38],stage1_14[44],stage1_13[68]}
   );
   gpc606_5 gpc198 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[38],stage1_15[39],stage1_14[45],stage1_13[69]}
   );
   gpc606_5 gpc199 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[39],stage1_15[40],stage1_14[46],stage1_13[70]}
   );
   gpc606_5 gpc200 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[40],stage1_15[41],stage1_14[47],stage1_13[71]}
   );
   gpc606_5 gpc201 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[41],stage1_15[42],stage1_14[48],stage1_13[72]}
   );
   gpc606_5 gpc202 (
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[42],stage1_15[43],stage1_14[49],stage1_13[73]}
   );
   gpc606_5 gpc203 (
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[43],stage1_15[44],stage1_14[50],stage1_13[74]}
   );
   gpc606_5 gpc204 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[44],stage1_15[45],stage1_14[51],stage1_13[75]}
   );
   gpc606_5 gpc205 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[45],stage1_15[46],stage1_14[52],stage1_13[76]}
   );
   gpc606_5 gpc206 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[46],stage1_15[47],stage1_14[53],stage1_13[77]}
   );
   gpc117_4 gpc207 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[156]},
      {1'b0},
      {stage1_17[26],stage1_16[47],stage1_15[48],stage1_14[54]}
   );
   gpc117_4 gpc208 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage0_15[157]},
      {1'b0},
      {stage1_17[27],stage1_16[48],stage1_15[49],stage1_14[55]}
   );
   gpc1_1 gpc209 (
      {stage0_0[160]},
      {stage1_0[31]}
   );
   gpc1_1 gpc210 (
      {stage0_0[161]},
      {stage1_0[32]}
   );
   gpc1_1 gpc211 (
      {stage0_2[152]},
      {stage1_2[54]}
   );
   gpc1_1 gpc212 (
      {stage0_2[153]},
      {stage1_2[55]}
   );
   gpc1_1 gpc213 (
      {stage0_2[154]},
      {stage1_2[56]}
   );
   gpc1_1 gpc214 (
      {stage0_2[155]},
      {stage1_2[57]}
   );
   gpc1_1 gpc215 (
      {stage0_2[156]},
      {stage1_2[58]}
   );
   gpc1_1 gpc216 (
      {stage0_2[157]},
      {stage1_2[59]}
   );
   gpc1_1 gpc217 (
      {stage0_2[158]},
      {stage1_2[60]}
   );
   gpc1_1 gpc218 (
      {stage0_2[159]},
      {stage1_2[61]}
   );
   gpc1_1 gpc219 (
      {stage0_2[160]},
      {stage1_2[62]}
   );
   gpc1_1 gpc220 (
      {stage0_2[161]},
      {stage1_2[63]}
   );
   gpc1_1 gpc221 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc222 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc223 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc224 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc225 (
      {stage0_3[128]},
      {stage1_3[58]}
   );
   gpc1_1 gpc226 (
      {stage0_3[129]},
      {stage1_3[59]}
   );
   gpc1_1 gpc227 (
      {stage0_3[130]},
      {stage1_3[60]}
   );
   gpc1_1 gpc228 (
      {stage0_3[131]},
      {stage1_3[61]}
   );
   gpc1_1 gpc229 (
      {stage0_3[132]},
      {stage1_3[62]}
   );
   gpc1_1 gpc230 (
      {stage0_3[133]},
      {stage1_3[63]}
   );
   gpc1_1 gpc231 (
      {stage0_3[134]},
      {stage1_3[64]}
   );
   gpc1_1 gpc232 (
      {stage0_3[135]},
      {stage1_3[65]}
   );
   gpc1_1 gpc233 (
      {stage0_3[136]},
      {stage1_3[66]}
   );
   gpc1_1 gpc234 (
      {stage0_3[137]},
      {stage1_3[67]}
   );
   gpc1_1 gpc235 (
      {stage0_3[138]},
      {stage1_3[68]}
   );
   gpc1_1 gpc236 (
      {stage0_3[139]},
      {stage1_3[69]}
   );
   gpc1_1 gpc237 (
      {stage0_3[140]},
      {stage1_3[70]}
   );
   gpc1_1 gpc238 (
      {stage0_3[141]},
      {stage1_3[71]}
   );
   gpc1_1 gpc239 (
      {stage0_3[142]},
      {stage1_3[72]}
   );
   gpc1_1 gpc240 (
      {stage0_3[143]},
      {stage1_3[73]}
   );
   gpc1_1 gpc241 (
      {stage0_3[144]},
      {stage1_3[74]}
   );
   gpc1_1 gpc242 (
      {stage0_3[145]},
      {stage1_3[75]}
   );
   gpc1_1 gpc243 (
      {stage0_3[146]},
      {stage1_3[76]}
   );
   gpc1_1 gpc244 (
      {stage0_3[147]},
      {stage1_3[77]}
   );
   gpc1_1 gpc245 (
      {stage0_3[148]},
      {stage1_3[78]}
   );
   gpc1_1 gpc246 (
      {stage0_3[149]},
      {stage1_3[79]}
   );
   gpc1_1 gpc247 (
      {stage0_3[150]},
      {stage1_3[80]}
   );
   gpc1_1 gpc248 (
      {stage0_3[151]},
      {stage1_3[81]}
   );
   gpc1_1 gpc249 (
      {stage0_3[152]},
      {stage1_3[82]}
   );
   gpc1_1 gpc250 (
      {stage0_3[153]},
      {stage1_3[83]}
   );
   gpc1_1 gpc251 (
      {stage0_3[154]},
      {stage1_3[84]}
   );
   gpc1_1 gpc252 (
      {stage0_3[155]},
      {stage1_3[85]}
   );
   gpc1_1 gpc253 (
      {stage0_3[156]},
      {stage1_3[86]}
   );
   gpc1_1 gpc254 (
      {stage0_3[157]},
      {stage1_3[87]}
   );
   gpc1_1 gpc255 (
      {stage0_3[158]},
      {stage1_3[88]}
   );
   gpc1_1 gpc256 (
      {stage0_3[159]},
      {stage1_3[89]}
   );
   gpc1_1 gpc257 (
      {stage0_3[160]},
      {stage1_3[90]}
   );
   gpc1_1 gpc258 (
      {stage0_3[161]},
      {stage1_3[91]}
   );
   gpc1_1 gpc259 (
      {stage0_8[147]},
      {stage1_8[75]}
   );
   gpc1_1 gpc260 (
      {stage0_8[148]},
      {stage1_8[76]}
   );
   gpc1_1 gpc261 (
      {stage0_8[149]},
      {stage1_8[77]}
   );
   gpc1_1 gpc262 (
      {stage0_8[150]},
      {stage1_8[78]}
   );
   gpc1_1 gpc263 (
      {stage0_8[151]},
      {stage1_8[79]}
   );
   gpc1_1 gpc264 (
      {stage0_8[152]},
      {stage1_8[80]}
   );
   gpc1_1 gpc265 (
      {stage0_8[153]},
      {stage1_8[81]}
   );
   gpc1_1 gpc266 (
      {stage0_8[154]},
      {stage1_8[82]}
   );
   gpc1_1 gpc267 (
      {stage0_8[155]},
      {stage1_8[83]}
   );
   gpc1_1 gpc268 (
      {stage0_8[156]},
      {stage1_8[84]}
   );
   gpc1_1 gpc269 (
      {stage0_8[157]},
      {stage1_8[85]}
   );
   gpc1_1 gpc270 (
      {stage0_8[158]},
      {stage1_8[86]}
   );
   gpc1_1 gpc271 (
      {stage0_8[159]},
      {stage1_8[87]}
   );
   gpc1_1 gpc272 (
      {stage0_8[160]},
      {stage1_8[88]}
   );
   gpc1_1 gpc273 (
      {stage0_8[161]},
      {stage1_8[89]}
   );
   gpc1_1 gpc274 (
      {stage0_9[157]},
      {stage1_9[78]}
   );
   gpc1_1 gpc275 (
      {stage0_9[158]},
      {stage1_9[79]}
   );
   gpc1_1 gpc276 (
      {stage0_9[159]},
      {stage1_9[80]}
   );
   gpc1_1 gpc277 (
      {stage0_9[160]},
      {stage1_9[81]}
   );
   gpc1_1 gpc278 (
      {stage0_9[161]},
      {stage1_9[82]}
   );
   gpc1_1 gpc279 (
      {stage0_10[158]},
      {stage1_10[57]}
   );
   gpc1_1 gpc280 (
      {stage0_10[159]},
      {stage1_10[58]}
   );
   gpc1_1 gpc281 (
      {stage0_10[160]},
      {stage1_10[59]}
   );
   gpc1_1 gpc282 (
      {stage0_10[161]},
      {stage1_10[60]}
   );
   gpc1_1 gpc283 (
      {stage0_11[156]},
      {stage1_11[52]}
   );
   gpc1_1 gpc284 (
      {stage0_11[157]},
      {stage1_11[53]}
   );
   gpc1_1 gpc285 (
      {stage0_11[158]},
      {stage1_11[54]}
   );
   gpc1_1 gpc286 (
      {stage0_11[159]},
      {stage1_11[55]}
   );
   gpc1_1 gpc287 (
      {stage0_11[160]},
      {stage1_11[56]}
   );
   gpc1_1 gpc288 (
      {stage0_11[161]},
      {stage1_11[57]}
   );
   gpc1_1 gpc289 (
      {stage0_14[140]},
      {stage1_14[56]}
   );
   gpc1_1 gpc290 (
      {stage0_14[141]},
      {stage1_14[57]}
   );
   gpc1_1 gpc291 (
      {stage0_14[142]},
      {stage1_14[58]}
   );
   gpc1_1 gpc292 (
      {stage0_14[143]},
      {stage1_14[59]}
   );
   gpc1_1 gpc293 (
      {stage0_14[144]},
      {stage1_14[60]}
   );
   gpc1_1 gpc294 (
      {stage0_14[145]},
      {stage1_14[61]}
   );
   gpc1_1 gpc295 (
      {stage0_14[146]},
      {stage1_14[62]}
   );
   gpc1_1 gpc296 (
      {stage0_14[147]},
      {stage1_14[63]}
   );
   gpc1_1 gpc297 (
      {stage0_14[148]},
      {stage1_14[64]}
   );
   gpc1_1 gpc298 (
      {stage0_14[149]},
      {stage1_14[65]}
   );
   gpc1_1 gpc299 (
      {stage0_14[150]},
      {stage1_14[66]}
   );
   gpc1_1 gpc300 (
      {stage0_14[151]},
      {stage1_14[67]}
   );
   gpc1_1 gpc301 (
      {stage0_14[152]},
      {stage1_14[68]}
   );
   gpc1_1 gpc302 (
      {stage0_14[153]},
      {stage1_14[69]}
   );
   gpc1_1 gpc303 (
      {stage0_14[154]},
      {stage1_14[70]}
   );
   gpc1_1 gpc304 (
      {stage0_14[155]},
      {stage1_14[71]}
   );
   gpc1_1 gpc305 (
      {stage0_14[156]},
      {stage1_14[72]}
   );
   gpc1_1 gpc306 (
      {stage0_14[157]},
      {stage1_14[73]}
   );
   gpc1_1 gpc307 (
      {stage0_14[158]},
      {stage1_14[74]}
   );
   gpc1_1 gpc308 (
      {stage0_14[159]},
      {stage1_14[75]}
   );
   gpc1_1 gpc309 (
      {stage0_14[160]},
      {stage1_14[76]}
   );
   gpc1_1 gpc310 (
      {stage0_14[161]},
      {stage1_14[77]}
   );
   gpc1_1 gpc311 (
      {stage0_15[158]},
      {stage1_15[50]}
   );
   gpc1_1 gpc312 (
      {stage0_15[159]},
      {stage1_15[51]}
   );
   gpc1_1 gpc313 (
      {stage0_15[160]},
      {stage1_15[52]}
   );
   gpc1_1 gpc314 (
      {stage0_15[161]},
      {stage1_15[53]}
   );
   gpc606_5 gpc315 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc316 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc317 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[0]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc318 (
      {stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21]},
      {stage1_1[1]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc319 (
      {stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[2]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc320 (
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc321 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc322 (
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc323 (
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc615_5 gpc324 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34]},
      {stage1_3[24]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc325 (
      {stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage1_3[25]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc326 (
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage1_3[26]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc327 (
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_3[27]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc328 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage1_3[28]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc329 (
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_3[29]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc330 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], 1'b0},
      {stage1_3[30]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc331 (
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc332 (
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc333 (
      {stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc334 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc335 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc336 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[16],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc337 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[17],stage2_4[22],stage2_3[22]}
   );
   gpc615_5 gpc338 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[49]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[14],stage2_5[18],stage2_4[23],stage2_3[23]}
   );
   gpc615_5 gpc339 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[50]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[15],stage2_5[19],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc340 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[51]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[16],stage2_5[20],stage2_4[25],stage2_3[25]}
   );
   gpc606_5 gpc341 (
      {stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[10],stage2_6[17],stage2_5[21],stage2_4[26]}
   );
   gpc606_5 gpc342 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[11],stage2_6[18],stage2_5[22],stage2_4[27]}
   );
   gpc606_5 gpc343 (
      {stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[12],stage2_6[19],stage2_5[23],stage2_4[28]}
   );
   gpc615_5 gpc344 (
      {stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_5[60]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[13],stage2_6[20],stage2_5[24],stage2_4[29]}
   );
   gpc606_5 gpc345 (
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[14],stage2_6[21],stage2_5[25]}
   );
   gpc606_5 gpc346 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[5],stage2_7[15],stage2_6[22]}
   );
   gpc606_5 gpc347 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[6],stage2_7[16],stage2_6[23]}
   );
   gpc606_5 gpc348 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[7],stage2_7[17],stage2_6[24]}
   );
   gpc606_5 gpc349 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[4],stage2_8[8],stage2_7[18],stage2_6[25]}
   );
   gpc615_5 gpc350 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52]},
      {stage1_7[6]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[5],stage2_8[9],stage2_7[19],stage2_6[26]}
   );
   gpc615_5 gpc351 (
      {stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57]},
      {stage1_7[7]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[6],stage2_8[10],stage2_7[20],stage2_6[27]}
   );
   gpc615_5 gpc352 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[7],stage2_8[11],stage2_7[21]}
   );
   gpc615_5 gpc353 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[8],stage2_8[12],stage2_7[22]}
   );
   gpc615_5 gpc354 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[9],stage2_8[13],stage2_7[23]}
   );
   gpc615_5 gpc355 (
      {stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[10],stage2_8[14],stage2_7[24]}
   );
   gpc615_5 gpc356 (
      {stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32]},
      {stage1_8[40]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[10],stage2_9[11],stage2_8[15],stage2_7[25]}
   );
   gpc615_5 gpc357 (
      {stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage1_8[41]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[11],stage2_9[12],stage2_8[16],stage2_7[26]}
   );
   gpc615_5 gpc358 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage1_8[42]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[12],stage2_9[13],stage2_8[17],stage2_7[27]}
   );
   gpc606_5 gpc359 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[7],stage2_10[13],stage2_9[14],stage2_8[18]}
   );
   gpc606_5 gpc360 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[8],stage2_10[14],stage2_9[15],stage2_8[19]}
   );
   gpc606_5 gpc361 (
      {stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[9],stage2_10[15],stage2_9[16],stage2_8[20]}
   );
   gpc606_5 gpc362 (
      {stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[10],stage2_10[16],stage2_9[17],stage2_8[21]}
   );
   gpc606_5 gpc363 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[11],stage2_10[17],stage2_9[18],stage2_8[22]}
   );
   gpc606_5 gpc364 (
      {stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[12],stage2_10[18],stage2_9[19],stage2_8[23]}
   );
   gpc606_5 gpc365 (
      {stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[13],stage2_10[19],stage2_9[20],stage2_8[24]}
   );
   gpc606_5 gpc366 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[7],stage2_11[14],stage2_10[20],stage2_9[21]}
   );
   gpc606_5 gpc367 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[8],stage2_11[15],stage2_10[21],stage2_9[22]}
   );
   gpc615_5 gpc368 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46]},
      {stage1_11[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[9],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc369 (
      {stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51]},
      {stage1_11[13]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[10],stage2_11[17],stage2_10[23]}
   );
   gpc615_5 gpc370 (
      {stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_11[14]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[11],stage2_11[18],stage2_10[24]}
   );
   gpc615_5 gpc371 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], 1'b0},
      {stage1_11[15]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[5],stage2_12[12],stage2_11[19],stage2_10[25]}
   );
   gpc1343_5 gpc372 (
      {stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27]},
      {stage1_13[0], stage1_13[1], stage1_13[2]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[4],stage2_13[6],stage2_12[13],stage2_11[20]}
   );
   gpc615_5 gpc373 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage1_12[28]},
      {stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage2_15[1],stage2_14[5],stage2_13[7],stage2_12[14],stage2_11[21]}
   );
   gpc615_5 gpc374 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[29]},
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage2_15[2],stage2_14[6],stage2_13[8],stage2_12[15],stage2_11[22]}
   );
   gpc615_5 gpc375 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[30]},
      {stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20]},
      {stage2_15[3],stage2_14[7],stage2_13[9],stage2_12[16],stage2_11[23]}
   );
   gpc615_5 gpc376 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[31]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[4],stage2_14[8],stage2_13[10],stage2_12[17],stage2_11[24]}
   );
   gpc615_5 gpc377 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[32]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[5],stage2_14[9],stage2_13[11],stage2_12[18],stage2_11[25]}
   );
   gpc615_5 gpc378 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[33]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[6],stage2_14[10],stage2_13[12],stage2_12[19],stage2_11[26]}
   );
   gpc615_5 gpc379 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[34]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[7],stage2_14[11],stage2_13[13],stage2_12[20],stage2_11[27]}
   );
   gpc615_5 gpc380 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], 1'b0},
      {stage1_12[35]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[8],stage2_14[12],stage2_13[14],stage2_12[21],stage2_11[28]}
   );
   gpc606_5 gpc381 (
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[9],stage2_14[13],stage2_13[15],stage2_12[22]}
   );
   gpc606_5 gpc382 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[10],stage2_14[14],stage2_13[16],stage2_12[23]}
   );
   gpc606_5 gpc383 (
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[11],stage2_14[15],stage2_13[17],stage2_12[24]}
   );
   gpc606_5 gpc384 (
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[12],stage2_14[16],stage2_13[18],stage2_12[25]}
   );
   gpc606_5 gpc385 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[13],stage2_14[17],stage2_13[19],stage2_12[26]}
   );
   gpc606_5 gpc386 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[18],stage2_13[20]}
   );
   gpc606_5 gpc387 (
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[19],stage2_13[21]}
   );
   gpc606_5 gpc388 (
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[20],stage2_13[22]}
   );
   gpc606_5 gpc389 (
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[21],stage2_13[23]}
   );
   gpc606_5 gpc390 (
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[22]}
   );
   gpc606_5 gpc391 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[23]}
   );
   gpc606_5 gpc392 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[24]}
   );
   gpc606_5 gpc393 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[25]}
   );
   gpc606_5 gpc394 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[26]}
   );
   gpc606_5 gpc395 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23],stage2_14[27]}
   );
   gpc606_5 gpc396 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24],stage2_14[28]}
   );
   gpc615_5 gpc397 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[24]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[11],stage2_16[16],stage2_15[25],stage2_14[29]}
   );
   gpc615_5 gpc398 (
      {stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[48]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[8],stage2_17[12],stage2_16[17],stage2_15[26]}
   );
   gpc1_1 gpc399 (
      {stage1_0[27]},
      {stage2_0[5]}
   );
   gpc1_1 gpc400 (
      {stage1_0[28]},
      {stage2_0[6]}
   );
   gpc1_1 gpc401 (
      {stage1_0[29]},
      {stage2_0[7]}
   );
   gpc1_1 gpc402 (
      {stage1_0[30]},
      {stage2_0[8]}
   );
   gpc1_1 gpc403 (
      {stage1_0[31]},
      {stage2_0[9]}
   );
   gpc1_1 gpc404 (
      {stage1_0[32]},
      {stage2_0[10]}
   );
   gpc1_1 gpc405 (
      {stage1_1[27]},
      {stage2_1[9]}
   );
   gpc1_1 gpc406 (
      {stage1_1[28]},
      {stage2_1[10]}
   );
   gpc1_1 gpc407 (
      {stage1_1[29]},
      {stage2_1[11]}
   );
   gpc1_1 gpc408 (
      {stage1_1[30]},
      {stage2_1[12]}
   );
   gpc1_1 gpc409 (
      {stage1_1[31]},
      {stage2_1[13]}
   );
   gpc1_1 gpc410 (
      {stage1_1[32]},
      {stage2_1[14]}
   );
   gpc1_1 gpc411 (
      {stage1_1[33]},
      {stage2_1[15]}
   );
   gpc1_1 gpc412 (
      {stage1_1[34]},
      {stage2_1[16]}
   );
   gpc1_1 gpc413 (
      {stage1_1[35]},
      {stage2_1[17]}
   );
   gpc1_1 gpc414 (
      {stage1_1[36]},
      {stage2_1[18]}
   );
   gpc1_1 gpc415 (
      {stage1_1[37]},
      {stage2_1[19]}
   );
   gpc1_1 gpc416 (
      {stage1_1[38]},
      {stage2_1[20]}
   );
   gpc1_1 gpc417 (
      {stage1_1[39]},
      {stage2_1[21]}
   );
   gpc1_1 gpc418 (
      {stage1_1[40]},
      {stage2_1[22]}
   );
   gpc1_1 gpc419 (
      {stage1_1[41]},
      {stage2_1[23]}
   );
   gpc1_1 gpc420 (
      {stage1_1[42]},
      {stage2_1[24]}
   );
   gpc1_1 gpc421 (
      {stage1_1[43]},
      {stage2_1[25]}
   );
   gpc1_1 gpc422 (
      {stage1_1[44]},
      {stage2_1[26]}
   );
   gpc1_1 gpc423 (
      {stage1_1[45]},
      {stage2_1[27]}
   );
   gpc1_1 gpc424 (
      {stage1_1[46]},
      {stage2_1[28]}
   );
   gpc1_1 gpc425 (
      {stage1_1[47]},
      {stage2_1[29]}
   );
   gpc1_1 gpc426 (
      {stage1_3[81]},
      {stage2_3[26]}
   );
   gpc1_1 gpc427 (
      {stage1_3[82]},
      {stage2_3[27]}
   );
   gpc1_1 gpc428 (
      {stage1_3[83]},
      {stage2_3[28]}
   );
   gpc1_1 gpc429 (
      {stage1_3[84]},
      {stage2_3[29]}
   );
   gpc1_1 gpc430 (
      {stage1_3[85]},
      {stage2_3[30]}
   );
   gpc1_1 gpc431 (
      {stage1_3[86]},
      {stage2_3[31]}
   );
   gpc1_1 gpc432 (
      {stage1_3[87]},
      {stage2_3[32]}
   );
   gpc1_1 gpc433 (
      {stage1_3[88]},
      {stage2_3[33]}
   );
   gpc1_1 gpc434 (
      {stage1_3[89]},
      {stage2_3[34]}
   );
   gpc1_1 gpc435 (
      {stage1_3[90]},
      {stage2_3[35]}
   );
   gpc1_1 gpc436 (
      {stage1_3[91]},
      {stage2_3[36]}
   );
   gpc1_1 gpc437 (
      {stage1_5[67]},
      {stage2_5[26]}
   );
   gpc1_1 gpc438 (
      {stage1_5[68]},
      {stage2_5[27]}
   );
   gpc1_1 gpc439 (
      {stage1_5[69]},
      {stage2_5[28]}
   );
   gpc1_1 gpc440 (
      {stage1_5[70]},
      {stage2_5[29]}
   );
   gpc1_1 gpc441 (
      {stage1_6[58]},
      {stage2_6[28]}
   );
   gpc1_1 gpc442 (
      {stage1_6[59]},
      {stage2_6[29]}
   );
   gpc1_1 gpc443 (
      {stage1_7[43]},
      {stage2_7[28]}
   );
   gpc1_1 gpc444 (
      {stage1_7[44]},
      {stage2_7[29]}
   );
   gpc1_1 gpc445 (
      {stage1_7[45]},
      {stage2_7[30]}
   );
   gpc1_1 gpc446 (
      {stage1_7[46]},
      {stage2_7[31]}
   );
   gpc1_1 gpc447 (
      {stage1_7[47]},
      {stage2_7[32]}
   );
   gpc1_1 gpc448 (
      {stage1_7[48]},
      {stage2_7[33]}
   );
   gpc1_1 gpc449 (
      {stage1_7[49]},
      {stage2_7[34]}
   );
   gpc1_1 gpc450 (
      {stage1_7[50]},
      {stage2_7[35]}
   );
   gpc1_1 gpc451 (
      {stage1_7[51]},
      {stage2_7[36]}
   );
   gpc1_1 gpc452 (
      {stage1_7[52]},
      {stage2_7[37]}
   );
   gpc1_1 gpc453 (
      {stage1_7[53]},
      {stage2_7[38]}
   );
   gpc1_1 gpc454 (
      {stage1_8[85]},
      {stage2_8[25]}
   );
   gpc1_1 gpc455 (
      {stage1_8[86]},
      {stage2_8[26]}
   );
   gpc1_1 gpc456 (
      {stage1_8[87]},
      {stage2_8[27]}
   );
   gpc1_1 gpc457 (
      {stage1_8[88]},
      {stage2_8[28]}
   );
   gpc1_1 gpc458 (
      {stage1_8[89]},
      {stage2_8[29]}
   );
   gpc1_1 gpc459 (
      {stage1_9[54]},
      {stage2_9[23]}
   );
   gpc1_1 gpc460 (
      {stage1_9[55]},
      {stage2_9[24]}
   );
   gpc1_1 gpc461 (
      {stage1_9[56]},
      {stage2_9[25]}
   );
   gpc1_1 gpc462 (
      {stage1_9[57]},
      {stage2_9[26]}
   );
   gpc1_1 gpc463 (
      {stage1_9[58]},
      {stage2_9[27]}
   );
   gpc1_1 gpc464 (
      {stage1_9[59]},
      {stage2_9[28]}
   );
   gpc1_1 gpc465 (
      {stage1_9[60]},
      {stage2_9[29]}
   );
   gpc1_1 gpc466 (
      {stage1_9[61]},
      {stage2_9[30]}
   );
   gpc1_1 gpc467 (
      {stage1_9[62]},
      {stage2_9[31]}
   );
   gpc1_1 gpc468 (
      {stage1_9[63]},
      {stage2_9[32]}
   );
   gpc1_1 gpc469 (
      {stage1_9[64]},
      {stage2_9[33]}
   );
   gpc1_1 gpc470 (
      {stage1_9[65]},
      {stage2_9[34]}
   );
   gpc1_1 gpc471 (
      {stage1_9[66]},
      {stage2_9[35]}
   );
   gpc1_1 gpc472 (
      {stage1_9[67]},
      {stage2_9[36]}
   );
   gpc1_1 gpc473 (
      {stage1_9[68]},
      {stage2_9[37]}
   );
   gpc1_1 gpc474 (
      {stage1_9[69]},
      {stage2_9[38]}
   );
   gpc1_1 gpc475 (
      {stage1_9[70]},
      {stage2_9[39]}
   );
   gpc1_1 gpc476 (
      {stage1_9[71]},
      {stage2_9[40]}
   );
   gpc1_1 gpc477 (
      {stage1_9[72]},
      {stage2_9[41]}
   );
   gpc1_1 gpc478 (
      {stage1_9[73]},
      {stage2_9[42]}
   );
   gpc1_1 gpc479 (
      {stage1_9[74]},
      {stage2_9[43]}
   );
   gpc1_1 gpc480 (
      {stage1_9[75]},
      {stage2_9[44]}
   );
   gpc1_1 gpc481 (
      {stage1_9[76]},
      {stage2_9[45]}
   );
   gpc1_1 gpc482 (
      {stage1_9[77]},
      {stage2_9[46]}
   );
   gpc1_1 gpc483 (
      {stage1_9[78]},
      {stage2_9[47]}
   );
   gpc1_1 gpc484 (
      {stage1_9[79]},
      {stage2_9[48]}
   );
   gpc1_1 gpc485 (
      {stage1_9[80]},
      {stage2_9[49]}
   );
   gpc1_1 gpc486 (
      {stage1_9[81]},
      {stage2_9[50]}
   );
   gpc1_1 gpc487 (
      {stage1_9[82]},
      {stage2_9[51]}
   );
   gpc1_1 gpc488 (
      {stage1_12[66]},
      {stage2_12[27]}
   );
   gpc1_1 gpc489 (
      {stage1_12[67]},
      {stage2_12[28]}
   );
   gpc1_1 gpc490 (
      {stage1_12[68]},
      {stage2_12[29]}
   );
   gpc1_1 gpc491 (
      {stage1_12[69]},
      {stage2_12[30]}
   );
   gpc1_1 gpc492 (
      {stage1_12[70]},
      {stage2_12[31]}
   );
   gpc1_1 gpc493 (
      {stage1_12[71]},
      {stage2_12[32]}
   );
   gpc1_1 gpc494 (
      {stage1_12[72]},
      {stage2_12[33]}
   );
   gpc1_1 gpc495 (
      {stage1_13[75]},
      {stage2_13[24]}
   );
   gpc1_1 gpc496 (
      {stage1_13[76]},
      {stage2_13[25]}
   );
   gpc1_1 gpc497 (
      {stage1_13[77]},
      {stage2_13[26]}
   );
   gpc1_1 gpc498 (
      {stage1_15[30]},
      {stage2_15[27]}
   );
   gpc1_1 gpc499 (
      {stage1_15[31]},
      {stage2_15[28]}
   );
   gpc1_1 gpc500 (
      {stage1_15[32]},
      {stage2_15[29]}
   );
   gpc1_1 gpc501 (
      {stage1_15[33]},
      {stage2_15[30]}
   );
   gpc1_1 gpc502 (
      {stage1_15[34]},
      {stage2_15[31]}
   );
   gpc1_1 gpc503 (
      {stage1_15[35]},
      {stage2_15[32]}
   );
   gpc1_1 gpc504 (
      {stage1_15[36]},
      {stage2_15[33]}
   );
   gpc1_1 gpc505 (
      {stage1_15[37]},
      {stage2_15[34]}
   );
   gpc1_1 gpc506 (
      {stage1_15[38]},
      {stage2_15[35]}
   );
   gpc1_1 gpc507 (
      {stage1_15[39]},
      {stage2_15[36]}
   );
   gpc1_1 gpc508 (
      {stage1_15[40]},
      {stage2_15[37]}
   );
   gpc1_1 gpc509 (
      {stage1_15[41]},
      {stage2_15[38]}
   );
   gpc1_1 gpc510 (
      {stage1_15[42]},
      {stage2_15[39]}
   );
   gpc1_1 gpc511 (
      {stage1_15[43]},
      {stage2_15[40]}
   );
   gpc1_1 gpc512 (
      {stage1_15[44]},
      {stage2_15[41]}
   );
   gpc1_1 gpc513 (
      {stage1_15[45]},
      {stage2_15[42]}
   );
   gpc1_1 gpc514 (
      {stage1_15[46]},
      {stage2_15[43]}
   );
   gpc1_1 gpc515 (
      {stage1_15[47]},
      {stage2_15[44]}
   );
   gpc1_1 gpc516 (
      {stage1_15[48]},
      {stage2_15[45]}
   );
   gpc1_1 gpc517 (
      {stage1_15[49]},
      {stage2_15[46]}
   );
   gpc1_1 gpc518 (
      {stage1_15[50]},
      {stage2_15[47]}
   );
   gpc1_1 gpc519 (
      {stage1_15[51]},
      {stage2_15[48]}
   );
   gpc1_1 gpc520 (
      {stage1_15[52]},
      {stage2_15[49]}
   );
   gpc1_1 gpc521 (
      {stage1_15[53]},
      {stage2_15[50]}
   );
   gpc1_1 gpc522 (
      {stage1_17[6]},
      {stage2_17[13]}
   );
   gpc1_1 gpc523 (
      {stage1_17[7]},
      {stage2_17[14]}
   );
   gpc1_1 gpc524 (
      {stage1_17[8]},
      {stage2_17[15]}
   );
   gpc1_1 gpc525 (
      {stage1_17[9]},
      {stage2_17[16]}
   );
   gpc1_1 gpc526 (
      {stage1_17[10]},
      {stage2_17[17]}
   );
   gpc1_1 gpc527 (
      {stage1_17[11]},
      {stage2_17[18]}
   );
   gpc1_1 gpc528 (
      {stage1_17[12]},
      {stage2_17[19]}
   );
   gpc1_1 gpc529 (
      {stage1_17[13]},
      {stage2_17[20]}
   );
   gpc1_1 gpc530 (
      {stage1_17[14]},
      {stage2_17[21]}
   );
   gpc1_1 gpc531 (
      {stage1_17[15]},
      {stage2_17[22]}
   );
   gpc1_1 gpc532 (
      {stage1_17[16]},
      {stage2_17[23]}
   );
   gpc1_1 gpc533 (
      {stage1_17[17]},
      {stage2_17[24]}
   );
   gpc1_1 gpc534 (
      {stage1_17[18]},
      {stage2_17[25]}
   );
   gpc1_1 gpc535 (
      {stage1_17[19]},
      {stage2_17[26]}
   );
   gpc1_1 gpc536 (
      {stage1_17[20]},
      {stage2_17[27]}
   );
   gpc1_1 gpc537 (
      {stage1_17[21]},
      {stage2_17[28]}
   );
   gpc1_1 gpc538 (
      {stage1_17[22]},
      {stage2_17[29]}
   );
   gpc1_1 gpc539 (
      {stage1_17[23]},
      {stage2_17[30]}
   );
   gpc1_1 gpc540 (
      {stage1_17[24]},
      {stage2_17[31]}
   );
   gpc1_1 gpc541 (
      {stage1_17[25]},
      {stage2_17[32]}
   );
   gpc1_1 gpc542 (
      {stage1_17[26]},
      {stage2_17[33]}
   );
   gpc1_1 gpc543 (
      {stage1_17[27]},
      {stage2_17[34]}
   );
   gpc1163_5 gpc544 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc545 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc546 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc547 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc548 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc615_5 gpc549 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc550 (
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage2_4[1]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc606_5 gpc551 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc552 (
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc553 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[4],stage3_6[4],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc554 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[5],stage3_6[5],stage3_5[8],stage3_4[10]}
   );
   gpc606_5 gpc555 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[4],stage3_7[6],stage3_6[6],stage3_5[9]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[5],stage3_7[7],stage3_6[7],stage3_5[10]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[6],stage3_7[8],stage3_6[8],stage3_5[11]}
   );
   gpc615_5 gpc558 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28]},
      {stage2_7[18]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[7],stage3_7[9],stage3_6[9]}
   );
   gpc615_5 gpc559 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[4],stage3_8[8],stage3_7[10]}
   );
   gpc615_5 gpc560 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[5],stage3_8[9],stage3_7[11]}
   );
   gpc615_5 gpc561 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[6],stage3_8[10],stage3_7[12]}
   );
   gpc615_5 gpc562 (
      {stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[7],stage3_8[11],stage3_7[13]}
   );
   gpc606_5 gpc563 (
      {stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[8],stage3_8[12]}
   );
   gpc606_5 gpc564 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[9],stage3_8[13]}
   );
   gpc606_5 gpc565 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[10],stage3_8[14]}
   );
   gpc606_5 gpc566 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[11]}
   );
   gpc606_5 gpc567 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[12]}
   );
   gpc606_5 gpc568 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[13]}
   );
   gpc615_5 gpc569 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46]},
      {stage2_10[18]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[6],stage3_11[10],stage3_10[11],stage3_9[14]}
   );
   gpc615_5 gpc570 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[7],stage3_11[11],stage3_10[12]}
   );
   gpc615_5 gpc571 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], 1'b0},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[5],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc572 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[6],stage3_12[9]}
   );
   gpc606_5 gpc573 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[2],stage3_14[3],stage3_13[7],stage3_12[10]}
   );
   gpc606_5 gpc574 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[3],stage3_14[4],stage3_13[8],stage3_12[11]}
   );
   gpc606_5 gpc575 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[4],stage3_14[5],stage3_13[9],stage3_12[12]}
   );
   gpc606_5 gpc576 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[5],stage3_14[6],stage3_13[10]}
   );
   gpc606_5 gpc577 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[5],stage3_15[6],stage3_14[7],stage3_13[11]}
   );
   gpc606_5 gpc578 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[6],stage3_15[7],stage3_14[8],stage3_13[12]}
   );
   gpc606_5 gpc579 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[7],stage3_15[8],stage3_14[9]}
   );
   gpc615_5 gpc580 (
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[8],stage3_15[9]}
   );
   gpc615_5 gpc581 (
      {stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[9],stage3_15[10]}
   );
   gpc615_5 gpc582 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[6],stage3_16[10],stage3_15[11]}
   );
   gpc615_5 gpc583 (
      {stage2_15[33], stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[7],stage3_16[11],stage3_15[12]}
   );
   gpc615_5 gpc584 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[8],stage3_16[12],stage3_15[13]}
   );
   gpc615_5 gpc585 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[11]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], 1'b0},
      {stage3_19[5],stage3_18[6],stage3_17[9],stage3_16[13],stage3_15[14]}
   );
   gpc606_5 gpc586 (
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[6],stage3_18[7],stage3_17[10],stage3_16[14]}
   );
   gpc1_1 gpc587 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc588 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc589 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc590 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc591 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc592 (
      {stage2_2[2]},
      {stage3_2[5]}
   );
   gpc1_1 gpc593 (
      {stage2_2[3]},
      {stage3_2[6]}
   );
   gpc1_1 gpc594 (
      {stage2_2[4]},
      {stage3_2[7]}
   );
   gpc1_1 gpc595 (
      {stage2_2[5]},
      {stage3_2[8]}
   );
   gpc1_1 gpc596 (
      {stage2_2[6]},
      {stage3_2[9]}
   );
   gpc1_1 gpc597 (
      {stage2_2[7]},
      {stage3_2[10]}
   );
   gpc1_1 gpc598 (
      {stage2_2[8]},
      {stage3_2[11]}
   );
   gpc1_1 gpc599 (
      {stage2_2[9]},
      {stage3_2[12]}
   );
   gpc1_1 gpc600 (
      {stage2_2[10]},
      {stage3_2[13]}
   );
   gpc1_1 gpc601 (
      {stage2_2[11]},
      {stage3_2[14]}
   );
   gpc1_1 gpc602 (
      {stage2_2[12]},
      {stage3_2[15]}
   );
   gpc1_1 gpc603 (
      {stage2_2[13]},
      {stage3_2[16]}
   );
   gpc1_1 gpc604 (
      {stage2_2[14]},
      {stage3_2[17]}
   );
   gpc1_1 gpc605 (
      {stage2_2[15]},
      {stage3_2[18]}
   );
   gpc1_1 gpc606 (
      {stage2_3[30]},
      {stage3_3[7]}
   );
   gpc1_1 gpc607 (
      {stage2_3[31]},
      {stage3_3[8]}
   );
   gpc1_1 gpc608 (
      {stage2_3[32]},
      {stage3_3[9]}
   );
   gpc1_1 gpc609 (
      {stage2_3[33]},
      {stage3_3[10]}
   );
   gpc1_1 gpc610 (
      {stage2_3[34]},
      {stage3_3[11]}
   );
   gpc1_1 gpc611 (
      {stage2_3[35]},
      {stage3_3[12]}
   );
   gpc1_1 gpc612 (
      {stage2_3[36]},
      {stage3_3[13]}
   );
   gpc1_1 gpc613 (
      {stage2_4[26]},
      {stage3_4[11]}
   );
   gpc1_1 gpc614 (
      {stage2_4[27]},
      {stage3_4[12]}
   );
   gpc1_1 gpc615 (
      {stage2_4[28]},
      {stage3_4[13]}
   );
   gpc1_1 gpc616 (
      {stage2_4[29]},
      {stage3_4[14]}
   );
   gpc1_1 gpc617 (
      {stage2_6[29]},
      {stage3_6[10]}
   );
   gpc1_1 gpc618 (
      {stage2_8[28]},
      {stage3_8[15]}
   );
   gpc1_1 gpc619 (
      {stage2_8[29]},
      {stage3_8[16]}
   );
   gpc1_1 gpc620 (
      {stage2_9[47]},
      {stage3_9[15]}
   );
   gpc1_1 gpc621 (
      {stage2_9[48]},
      {stage3_9[16]}
   );
   gpc1_1 gpc622 (
      {stage2_9[49]},
      {stage3_9[17]}
   );
   gpc1_1 gpc623 (
      {stage2_9[50]},
      {stage3_9[18]}
   );
   gpc1_1 gpc624 (
      {stage2_9[51]},
      {stage3_9[19]}
   );
   gpc1_1 gpc625 (
      {stage2_10[24]},
      {stage3_10[13]}
   );
   gpc1_1 gpc626 (
      {stage2_10[25]},
      {stage3_10[14]}
   );
   gpc1_1 gpc627 (
      {stage2_12[31]},
      {stage3_12[13]}
   );
   gpc1_1 gpc628 (
      {stage2_12[32]},
      {stage3_12[14]}
   );
   gpc1_1 gpc629 (
      {stage2_12[33]},
      {stage3_12[15]}
   );
   gpc1_1 gpc630 (
      {stage2_13[24]},
      {stage3_13[13]}
   );
   gpc1_1 gpc631 (
      {stage2_13[25]},
      {stage3_13[14]}
   );
   gpc1_1 gpc632 (
      {stage2_13[26]},
      {stage3_13[15]}
   );
   gpc1_1 gpc633 (
      {stage2_15[48]},
      {stage3_15[15]}
   );
   gpc1_1 gpc634 (
      {stage2_15[49]},
      {stage3_15[16]}
   );
   gpc1_1 gpc635 (
      {stage2_15[50]},
      {stage3_15[17]}
   );
   gpc1_1 gpc636 (
      {stage2_18[6]},
      {stage3_18[8]}
   );
   gpc1_1 gpc637 (
      {stage2_18[7]},
      {stage3_18[9]}
   );
   gpc1_1 gpc638 (
      {stage2_18[8]},
      {stage3_18[10]}
   );
   gpc1_1 gpc639 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc615_5 gpc640 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc641 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[1]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc615_5 gpc642 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[2],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc643 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[3],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc644 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[2],stage4_6[4]}
   );
   gpc615_5 gpc645 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[3],stage4_6[5]}
   );
   gpc615_5 gpc646 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage3_8[12]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[4]}
   );
   gpc615_5 gpc647 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[13]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc648 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc649 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3],stage4_10[5]}
   );
   gpc606_5 gpc650 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4],stage4_10[6]}
   );
   gpc1406_5 gpc651 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc615_5 gpc652 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[0]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[1],stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[4]}
   );
   gpc615_5 gpc653 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[1]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[2],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[5]}
   );
   gpc606_5 gpc654 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage4_18[0],stage4_17[3],stage4_16[3],stage4_15[3],stage4_14[5]}
   );
   gpc615_5 gpc655 (
      {stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[4],stage4_16[4]}
   );
   gpc623_5 gpc656 (
      {stage3_16[12], stage3_16[13], stage3_16[14]},
      {stage3_17[1], stage3_17[2]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], 1'b0},
      {stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[5],stage4_16[5]}
   );
   gpc615_5 gpc657 (
      {stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[2],stage4_18[3],stage4_17[6]}
   );
   gpc1_1 gpc658 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc659 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc660 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc661 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc662 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc663 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc664 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc665 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc666 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc667 (
      {stage3_1[2]},
      {stage4_1[2]}
   );
   gpc1_1 gpc668 (
      {stage3_1[3]},
      {stage4_1[3]}
   );
   gpc1_1 gpc669 (
      {stage3_1[4]},
      {stage4_1[4]}
   );
   gpc1_1 gpc670 (
      {stage3_2[10]},
      {stage4_2[2]}
   );
   gpc1_1 gpc671 (
      {stage3_2[11]},
      {stage4_2[3]}
   );
   gpc1_1 gpc672 (
      {stage3_2[12]},
      {stage4_2[4]}
   );
   gpc1_1 gpc673 (
      {stage3_2[13]},
      {stage4_2[5]}
   );
   gpc1_1 gpc674 (
      {stage3_2[14]},
      {stage4_2[6]}
   );
   gpc1_1 gpc675 (
      {stage3_2[15]},
      {stage4_2[7]}
   );
   gpc1_1 gpc676 (
      {stage3_2[16]},
      {stage4_2[8]}
   );
   gpc1_1 gpc677 (
      {stage3_2[17]},
      {stage4_2[9]}
   );
   gpc1_1 gpc678 (
      {stage3_2[18]},
      {stage4_2[10]}
   );
   gpc1_1 gpc679 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc680 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc681 (
      {stage3_4[14]},
      {stage4_4[4]}
   );
   gpc1_1 gpc682 (
      {stage3_6[10]},
      {stage4_6[6]}
   );
   gpc1_1 gpc683 (
      {stage3_7[12]},
      {stage4_7[6]}
   );
   gpc1_1 gpc684 (
      {stage3_7[13]},
      {stage4_7[7]}
   );
   gpc1_1 gpc685 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc686 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc687 (
      {stage3_8[16]},
      {stage4_8[6]}
   );
   gpc1_1 gpc688 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc689 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc690 (
      {stage3_10[12]},
      {stage4_10[7]}
   );
   gpc1_1 gpc691 (
      {stage3_10[13]},
      {stage4_10[8]}
   );
   gpc1_1 gpc692 (
      {stage3_10[14]},
      {stage4_10[9]}
   );
   gpc1_1 gpc693 (
      {stage3_11[6]},
      {stage4_11[5]}
   );
   gpc1_1 gpc694 (
      {stage3_11[7]},
      {stage4_11[6]}
   );
   gpc1_1 gpc695 (
      {stage3_11[8]},
      {stage4_11[7]}
   );
   gpc1_1 gpc696 (
      {stage3_11[9]},
      {stage4_11[8]}
   );
   gpc1_1 gpc697 (
      {stage3_11[10]},
      {stage4_11[9]}
   );
   gpc1_1 gpc698 (
      {stage3_11[11]},
      {stage4_11[10]}
   );
   gpc1_1 gpc699 (
      {stage3_11[12]},
      {stage4_11[11]}
   );
   gpc1_1 gpc700 (
      {stage3_12[12]},
      {stage4_12[3]}
   );
   gpc1_1 gpc701 (
      {stage3_12[13]},
      {stage4_12[4]}
   );
   gpc1_1 gpc702 (
      {stage3_12[14]},
      {stage4_12[5]}
   );
   gpc1_1 gpc703 (
      {stage3_12[15]},
      {stage4_12[6]}
   );
   gpc1_1 gpc704 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc705 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc706 (
      {stage3_15[16]},
      {stage4_15[4]}
   );
   gpc1_1 gpc707 (
      {stage3_15[17]},
      {stage4_15[5]}
   );
   gpc1_1 gpc708 (
      {stage3_17[8]},
      {stage4_17[7]}
   );
   gpc1_1 gpc709 (
      {stage3_17[9]},
      {stage4_17[8]}
   );
   gpc1_1 gpc710 (
      {stage3_17[10]},
      {stage4_17[9]}
   );
   gpc1_1 gpc711 (
      {stage3_19[6]},
      {stage4_19[3]}
   );
   gpc1_1 gpc712 (
      {stage3_19[7]},
      {stage4_19[4]}
   );
   gpc1_1 gpc713 (
      {stage3_20[0]},
      {stage4_20[3]}
   );
   gpc606_5 gpc714 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc615_5 gpc715 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1343_5 gpc716 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0], stage4_8[1], stage4_8[2]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0]}
   );
   gpc1343_5 gpc717 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc1343_5 gpc718 (
      {stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc7_3 gpc719 (
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], 1'b0},
      {stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc1343_5 gpc720 (
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc207_4 gpc721 (
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], 1'b0},
      {stage4_13[3], stage4_13[4]},
      {stage5_14[1],stage5_13[2],stage5_12[3],stage5_11[3]}
   );
   gpc615_5 gpc722 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc615_5 gpc723 (
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {1'b0},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1],stage5_15[2]}
   );
   gpc1_1 gpc724 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc725 (
      {stage4_2[7]},
      {stage5_2[2]}
   );
   gpc1_1 gpc726 (
      {stage4_2[8]},
      {stage5_2[3]}
   );
   gpc1_1 gpc727 (
      {stage4_2[9]},
      {stage5_2[4]}
   );
   gpc1_1 gpc728 (
      {stage4_2[10]},
      {stage5_2[5]}
   );
   gpc1_1 gpc729 (
      {stage4_4[0]},
      {stage5_4[2]}
   );
   gpc1_1 gpc730 (
      {stage4_4[1]},
      {stage5_4[3]}
   );
   gpc1_1 gpc731 (
      {stage4_4[2]},
      {stage5_4[4]}
   );
   gpc1_1 gpc732 (
      {stage4_4[3]},
      {stage5_4[5]}
   );
   gpc1_1 gpc733 (
      {stage4_4[4]},
      {stage5_4[6]}
   );
   gpc1_1 gpc734 (
      {stage4_5[0]},
      {stage5_5[1]}
   );
   gpc1_1 gpc735 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc736 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc737 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc738 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc739 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc740 (
      {stage4_9[5]},
      {stage5_9[3]}
   );
   gpc1_1 gpc741 (
      {stage4_9[6]},
      {stage5_9[4]}
   );
   gpc1_1 gpc742 (
      {stage4_12[5]},
      {stage5_12[4]}
   );
   gpc1_1 gpc743 (
      {stage4_12[6]},
      {stage5_12[5]}
   );
   gpc1_1 gpc744 (
      {stage4_13[5]},
      {stage5_13[3]}
   );
   gpc1_1 gpc745 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc746 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc747 (
      {stage4_17[6]},
      {stage5_17[2]}
   );
   gpc1_1 gpc748 (
      {stage4_17[7]},
      {stage5_17[3]}
   );
   gpc1_1 gpc749 (
      {stage4_17[8]},
      {stage5_17[4]}
   );
   gpc1_1 gpc750 (
      {stage4_17[9]},
      {stage5_17[5]}
   );
   gpc1_1 gpc751 (
      {stage4_18[0]},
      {stage5_18[2]}
   );
   gpc1_1 gpc752 (
      {stage4_18[1]},
      {stage5_18[3]}
   );
   gpc1_1 gpc753 (
      {stage4_18[2]},
      {stage5_18[4]}
   );
   gpc1_1 gpc754 (
      {stage4_18[3]},
      {stage5_18[5]}
   );
   gpc1_1 gpc755 (
      {stage4_19[0]},
      {stage5_19[1]}
   );
   gpc1_1 gpc756 (
      {stage4_19[1]},
      {stage5_19[2]}
   );
   gpc1_1 gpc757 (
      {stage4_19[2]},
      {stage5_19[3]}
   );
   gpc1_1 gpc758 (
      {stage4_19[3]},
      {stage5_19[4]}
   );
   gpc1_1 gpc759 (
      {stage4_19[4]},
      {stage5_19[5]}
   );
   gpc1_1 gpc760 (
      {stage4_20[0]},
      {stage5_20[0]}
   );
   gpc1_1 gpc761 (
      {stage4_20[1]},
      {stage5_20[1]}
   );
   gpc1_1 gpc762 (
      {stage4_20[2]},
      {stage5_20[2]}
   );
   gpc1_1 gpc763 (
      {stage4_20[3]},
      {stage5_20[3]}
   );
   gpc1_1 gpc764 (
      {stage4_21[0]},
      {stage5_21[0]}
   );
   gpc615_5 gpc765 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc766 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0]},
      {stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc767 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc1163_5 gpc768 (
      {stage5_11[1], stage5_11[2], stage5_11[3]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_13[0]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1343_5 gpc769 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc770 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1]}
   );
   gpc1406_5 gpc771 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[1]}
   );
   gpc1_1 gpc772 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc773 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc774 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc775 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc776 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc777 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc778 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc779 (
      {stage5_7[1]},
      {stage6_7[1]}
   );
   gpc1_1 gpc780 (
      {stage5_9[4]},
      {stage6_9[1]}
   );
   gpc1_1 gpc781 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc782 (
      {stage5_16[1]},
      {stage6_16[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor_CLA162_16 compressor_CLA162_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h653feda2e2d5f17a579ab0c7e08e3135b769bd50d7f78143b27056354d35dfd87b0de1b6cba33ef3d74e05139ec369f31fc17606bedc8a6921ea7f241d6654ed3fe7aecce121089835c8c5fe150abc4f5b57f8c22cea35482cf935188c11d2623a82ffafbd245d228a34987e762faeb725d3c2c87e375a7899928f42672d4d35f461f838517668612da0f775710567539a8d49546ab11f5ae18643c1396f4fb6b5f9b51751fc8f66271a5b070f5f40a9fe0b7be1259cf15316f3e6eb2bbcbba3805f604ee59e375ac688d69075e25fceb1b470015c1caa67c2035f47bccf98c6122abc08bd5742cf95384867b94a5f191db07332d33f93b84190bc95bbaec0647806fdddb4213aeed44de7e8bba1a949cff734c93679e18bd034c613eb086fce8050a0635f70a245a750e862d782663d35d0f927d9cde1a3b322d1c79c2a08210d2c2bd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfab23f13e9452b26ab1fa8b3b894edf482e401e3b93631dab200e3ddbfd1e7bf9f43c818b960b237c19ace945fc952e2d4cd3df2f3b167a3515895502f75326d59a6af4408d7ee5175f0db25c717dde5ebbfcc817909cdec379e9f702da876807d8ff658a6ecf1e7c6cd1ae914616570b306866394f48d0b6193577b072abf6244d1fd3c17200e747406abb8aef82fb98695418a6d05a78e91da07b04e88b50847a482f21b0751cbc6dc5a4dadaad80b7ca38eedc855649c22c70ec4cf0150659df1c70f0a3769a204aaf6050c60a23df8bdf19380fa18599fb03f49f4cb2e7ccba57237966b052544b20d2c936e1b3de3cfb59f9c2953d43152e7760c75b878968f30a3e0406b33e90cb74f7a8213f48f48ad656d4441fe0e4534c216f04fa220378d83f8145578dbb16436ce817ea2db99bf835334d36cae4479810432a21c8301d2cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8e9aa943d3db49b5b0b46fb397090af6dc121a74e984f772000abc00afd1232f1bf9edc31311fd025076470d227c59f7aafdc93cccb2fc29ecdccabe3b5a80dccc0d1984c3e02f0e2d3df93f8c8a587f4b0bc19c77f67122b33fffb84a780b375082694a119200cafebea701e9dca196830bed655f1ebcfa9b7be279d6ee32c803355b8c6a22918232c42cc62c10241f00df5058203cd55404ed5fb3f16a1e57161a31806d5226705c777c7a34ca3a60ac85d54fb4d9921d1a1e3b96f9ac300108427aa8556b5402e67a59e95bc52825c50a9f70fa557ab5f000346280de5431a4fb8c9da1da17a9036ba3ca08ea978c46944a0e2edb91a4b6242109342fddc7cc766e7014a21d8d40a4db02e425110f0e933ff9976d5406a3105df05e21d88fd13aa11cfc18fd8fc859676a460af963b2e47624b588e51fc27c749efc212d77ad032ef2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h306c219fcbef42400391f15b28139a68fa96badcc2b4eb8399df4ce1e0767675c53b639855730c107c8074979963116e7eb1e6f18c70ca89875fd48a7e9065262a46c44fb4659424428fa47881b4655890dc2c8ab2ed2cbdfc96dce01c477da0ec20736a2fc99a116b2a4626122006133172019802baf20f22c29d92d063ed20f35f54bfc84da3435483f719958a7eb3a237e1f97380d1280601c8d41e6465082b1a1500e3827693e38c3250ff7b918a6695dc2c9ed555f26e5a74f9b789ac638e1f0b85bb4c69169a85175fa2db67778c5ca04d6dcbb14c4888e05730c9a63a90538c7aad88344f0543c0711b53b1e6544589b3847f34a6ed77e20ac849d817b223937153892859821a3414137ab6894f043f4194a7df8db6c47c8f8630c7b2ba83039d6d103c2317ca078d9886147eb21d99bc16fb670b3c09c3b53f4d0e931bb810ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'haac768246972610d1be7070d25bdc489606a2e9afc9dbe9da901091cc265fab52a9d6c0eb795aa27ee1bed90f54a27a78413cb6ea0b7f0c44606da834d46d8c08fbb56461aaa4ef7b6eadcd73b29a0608fb4a62ec04bd24b6603bb7fce7a569bba094c26e7153fd787ee90e8d7e5987919064565ab67f5a96b1732ca65bebdb283d6ef60bebbab8b567a2a0f06c2effc733bd594f263676935ffea073fb06addbf03756bd2a9e22e61be189c92339d39eae85894f66db1555b3cb905528ccc441a1c75863aab81e16bb33a442832fa4cbeb88f337a50d67b0d822f96e359e72833eab72c32061c1422d0b34b932f0a754352603e4d54e572d66fc96e49b3ee043da15e5c408a8698c26ca56aa9055ba7a697a9c7911632479854b4ee648daabad482ff035b9071fcf9a72ebfac40aebb76ae64e019358e717d6cc8a5cbb35f68dc6ce5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1fa42329efeb62526f0b16a6f732876c3f93d12d54273bd924f9cfd73327aa1692d7221cfbe41347f932f6e5b8dd84fb49fe8741123dc435a12bb97e2bcaaf1255dd43352bbb3b1f352f552457f56d36db00b00c96d7ab5517124f507be50c011118faa389b962ee7b076c24f5e1920718924a8be30f57423196c3749abddbc623709476e230a91eeb2e60b1add410365858224310d60828d71463f32cdf891019a95af6711caf507d0f1501b6b3e6cec1bf51fce9da2038129710c124f8b264eec242d8d445952df9d699d459b8134beba72da94a4ea21708366277032e9a35a06ec2dd1cccc15db317602eccee7faafa0020fefe771637e7a0a608c2201bbd0ba8861a44929863f478dce4d032200da45798a6ecda2185ee3655351ac3d46636e0febaa29ab2ece7111340fc1fa1d6b0129e9887b10eabbef692586befdca4fd5cd97e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hcab22ee3dfa3ec7ed84b93b47524cc76220af9f652bf07e8593f8eb93f23e6ac0a21d573f0b89212f28be6909c66cd35e55ba8cf9841debc06f1ae65f2abbddc6fe8a98aa2414780b150886a10a4f1ece4f174b7298a3458881953b31d9836371aa631652f07b76776fcae7c436a1034c39481ab8161d5b24a4e1dbd10f8f718b16c5b685d9258b4381a0f9813cd830bcae00b2348bfab6ad4a4bc2bf91dacfe073576b473fe86a5696380baf71931f8a876cf8931eb28ec2c62d4a1ac5ebb2ce534464080d49270a5e3e91708284f49798fcee6d59dba35310a23065912ff19cbd898673467d3e821681fb46f1b34dfff3b686b8d6bc0de645f4b0ff0d7916091f1ff63ab4512c861cfc4cc0d07bba2944ebab351bfaa0d935b781ac31bcc49402e60c83d28a724938d892b161cbba7b13eb698b9569591898ef8bd073ad83f2943ff5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb8569454b681ad3f148bea84b41eac6d1bf32d387eae3d98dc2f78fbff1471961552f83295af901362f8681d9df354c4bd565f86d9907072a41b11d1fe80324caf277b251e49f830639180099141a9679fb3d08c10aa19b84ace36eee64b80b1b668240990b1bdaad73215b6c3c2f2258362e6226214e77d09ba6ecb721d74bf180b2709ce633eca313feced417d1730ffe181deba302187fe123b1f0a6e0a92122b05841ef63faa4da2ff9f770e875d23ecb70f398b344fba451ff5e29606057543f57bfa3db6070f6a946b06efb82592d2f1f7f35b3456a365fbeb913a3d77d8223e5507796124ba26f9487c037f0fa98ab5b522f630f4bcd4521bb3601e14fb64bad35057679849c3cbaae8464d09df302968f2d090281de25cdfbb279aafbb0c41d01d74567ab11ddee396e753f81e7d1b44763aa8e46730be36524ad80924af6a2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc9ddacc0d949f8cc1ed27a176114cc7c86d7bb9c82384d2eac89430ad8f08f408ad8073864696ec0744b8b10a1bd0817fb6d3f16dc59e22558287f05193d4605d06e1480c5ac44ce6d0078874e8bbeb79b263449aa1e6f1044602e0a95866f9686626df522e2ed09973d4aae077a1a33b27c41088d5ddff4a33cadf75e84b16a7be67f530d562cbd1a74c0b4fd183efd061aab501fd6db757d457f04e3c22f35cd6fd96415ac7a7ea5eeb47983ef98db90a60942da06ab3a96a08173327a19cce8b83a5ca17003a7bd02a09cc66a80957972bbc5795d8866eb3332118b8f4a25e4326827fcafd82abccc404baec26f0b4a83eef2851359a94d5d0257c30e67014cb9395264b0d58b6afda76a8cb4338bbe551a8e129f9c73780229583b8688448adf40fbf92cd82f143c6d24103a555280058540e8459c2b536528b2f75620f68d3453a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'haabfa0503df910f1a00250468a1bd3511d7204cac9373a4e7d872cc25165922993280d2115e27f3db7a0de33314e26f0bb4a6eeb0088e39744198346b201ed331e3cff615153763f848d9db5e525553d635cc007f386e54679121f43b7d9675b8b7295373d22f0a15e205d17a3616702dd8bb6b96c693d12821ccef2598e708a67f12c5e97c21096fde643a868442b89d623e525fa30ddfa47f669d0a1227b9e5f6dc625ac61d51a27801f845bb9786abe131e7f66ac6eeeea7f13b7775b44756240c030fce5c11d36b2e03512cacaf053a824530edce49535df818811c9a40428c73d90da1cd7b353b61f73e4957e61ad2416ed01166375726a2e1fb140535d95bf7f40229212523f687f6e13f10d6757fde962425e375f3e19f60e707aa3a3252e0cbbda9af34ddd4f2bb2d3d8f8cd3c0a004dec7e652525981eceb3c3a0d9c7a46ad1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hcf9e6c72a14dccf6d6e24784b0a64a5c640270e42a9a13008edfcb9c846987e8c706189aa231213c8be5e69519eca9a6fe6c47dbcec7a100a44af7f2b23abbd4b8e40679844c5d8190933e3cfb26c5d8450a9044aa36de7725b254ed146cc297d9969cbab294d717650a5970ae597ff7372c5ed019087153a0e18d6f0bd82971cd17598441d2efbea266f3efe9aab8005d34fc498632a2d50dc95288c4792d6d38530d57beeaf2522e75cac97b28bfa903cd552b216390f16bb1ce37c0eb31d1dedd211ac0bc06ee21dcea0424cee17ad6fd96513dd55ef9ced98bc27588819318edd018d13fb00808cb430205b81fa87570f96e513ed421443537e1d403d4fda107c20a28679541f689cfa34276630a0d3abbb4c1e3b18a1999e0e7a90dfab26fe77fd96de5a01e2c0f128e7fc4da6b6f996f58f899b0767ca4ff0949dc5fdeec290e04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h62130febcca7b0f19dc46be6423e89392fce4408566c7aed1c782138d2fb9c3e74df51b21ee3703f058937458463df6bebec6602362e7a819c350f947390564a85e0c054669ca1003295159b1ff76bd30de3df1ef14b0bdeb6d5d3422330ba44a258ddc89655eb59634323f53617a5e9e4ceb7427f43d13d3529c8c3802cbb83c1202c8abc5db131a6fd786874ff375fe3af381e02c4491b322e02f6eed50748e548ba6a31346d02bb9cca06c6f6c48d4708c55cb9b0935b76b71fd4c244d89c7828c859fe15d4553bfd6c8c3eb2fbf1f5d6be385072751ac6761a1fca3c9813ac1042f8cc45e03f1ba9442675555758a1bc284c95cb42aee645a378bec30113e47a22513ddd183049a9fe387a66fa1f3b579d06873b8178a3016fc8c5adb2697ecb6150e5c0bae3e2e3b97ceee02a7b669396dd31e79708c2ec68a74e497cf2a1095982;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1d9a5172d90ce2b28a466e25b00cb631583c2a3458e4224c5b79ad93d0b91ab80790289841db03f25451a87a7cc63923fa85ab7c5c6e589dde5c318e9d7c739ea561ac15db1e3331dc1bab39984548e04872c7adf42ce5a4636a7a8a2d4229d5d5c2e7477b0c8a55bf0a8b633dfd4aefaa1f488a082e6bd33278d0c7c48a310ee7e3f6260ca16778c11a7b3d09210f2a41de32a3e551e220c2192ca55e4577c4e0bd754617b4afb67e6daf2b77230a73fa130246c0eef0d0d792337c8391d006b86b7ad235731a79c76f2a4da633bcb918cbb1451ef17bcc2922f209a71bfa8727e55f4d6a60a8be8f446a8fbbc709bf4ee8e30db23121a27eace56c587defe66176a61f38bdc648c0906b98e64c8490cae0647b9f18a512bfc4e6056f30b72a252d4360a1a034493516bfb40e3e7256187ccbee6bf4a035e225b691d19f5e058b3af04c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2cabbbee8560adf4a679d8be6d3a83374fd649ae9b4934765c3c1038c68a6d4ad458df799c550682dda2d09d7b3693dcb2932d02b145fc69590c22a3bce1fc571e0bd73a5c4b4e3a849cca6c5ca03149560212dc9425068caf618930407d57d1dc0bc5a98cc7bbd475b062bc320676bf41ebeae509814968b044b5dca9076e1b310435818818104425c59ec9d870be444c929dd8ad5d0e9dd4f084759519bd68f1c8be0ac4dbdc97d675bda8cd6f5acf49894cc46ac195d57e94092d0de762e226d9b5fe4e11b4e88f823b5a4adcd867a8d3f981c776db95e16b11ae52c181a3d37dcceb216e090ca81fae6f8b6e8f3a16b512f4a348b2d54f5293130b5b6b7229197449d4975fec200ad85c941193af83bca49c852362bae1e9e04b50640c50d3d65f2c20043e4a5329dd7f31e6e85c6edbb4fba50c7af56992a3a49699f6a889d20a67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4297d9b2f65ce5f39199d9ba8f9bb37bcd135ff43d28cc3cbfa91b5dacd8731b12ba7764f7274984bbd13ba106b153767be2cae828961860fc375608388dcd710032134647c8e8bd83b622d4e97397461e93b0b13d40df2020b680818b88b568d879385e3b7c23a245aca069f34663ca763a2d970f3a083d090a1f4dd0d6153d062f2ea7fef5fb3f5f08548557f2e6a0872fb728305da035b07b1c3ffcbb83c26e7bc28fcd7f2248a812c7ec0190cc9b29d612df160aa5ccb3bdef26384839585ee0cec5283c1792896551e7311aa3bb4653c60e65a6ae1b7ddb751f9aa05f755df221fa713cca53093789c99f29a553baaad0479b24e572abdfcbdd89a11036fbecbdb590817aed1c174d5ab77932427893451c51b56f1081c52e4da5641b44ff2ecc50fae5cb6ed7c2bc7b01f858cb353d6b79a0cd0f189b9dd6fd16f4b3a7af5fad99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hba2d4c0f7a932d52bfc5d4152b2572e038da715bb1ff6936d87ef29c6ef7005d49952c868bb870e67bab16425b7a74bb45888cf0e067e86bae98d5aee8fb461bbb0c6661d429111082cc6c9c92b8dffbefbdc7588b66c3aecc27d71b735b6a20ef587b64ce94fe2279064ac277e93260db28293542e3b26cf79165c98c181635f82eb625d2860d65dd4f9e179ccbec2f06ade649f59f9faa3cf19ac00664f557edc71984192dc532bdebeae3431313cce52d07e740213fb4dededd05ec32979e008e602935c5d478294b2fdc0016a465cb2019b4fe3ab09c1aa3e90b52afd7e299d53e63c5b05dfee7dcfb5fd794969b1fd753037ccce15fc775fa51fb67e14723a4c60bc0eb497474d549991abf8cbfef8f64f425472103aee2fc05771bbff60c5d619fc62cc9c48eaf13006772b50f60b530675123140384916e4b9cade56e1423bece;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5efe68bcce520bbc955f443c4bbafbe0a4e1c57286b04b99099743f4eecd1f2be95c88b7fa66a02742e57b67a3590b4453693247ed4e13f12d0eb1cab4b91e35d5c6dbd74a1446789ef2e00ba41453de0a16ab50bb03f850798802ba7f4b2e857359c9ddf4b8649927152f8ae186046c6e1ea9bf8d26651384b508a6292892124d30cc54ec1eadb78a7e0d939a50b4fe469534dbc506b621dd3ce89101afddfab7ca8d9df5dcb8f85d9af7472f314e1f5ee463ac604a563c69e4d8e0bbbd4c8596da04241681d4e7d44d832e85d290003ef72fa6e7fb371b43aa91dbe4b44b5735a16e9a921a236fb65c99d59748b3be00e60474d542df490ce69f0148bb0740ed5861b01bd72bbc229fd62965331414e979accbae8a8412decbe28daf73a6874d8600b0786cdb034fc247282740da849916c5f7c8e615af17a906f79f15aa11fa273b00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1d29637018da59cf8921f505c0c0a72bf122e19a789a424b1ce4bdc96ab11f09f78916da00452962aca64f9482aa4b92c8dcd89f6818df2380ddf63b695c7ac37260cea1f21f03bf0a387e874f6cd9f7d03915657cc7249dba192d65cf90757bbf8871b63810f097517c201b9744a2464ea1937066717b31bd9d09711b19b0f4be77b3509110472d43d622b237f2ad738efd2d09f4079358dc3887787f63979b2617b56e89f0e9dfcfe0aa9883666068f786632e45d389c60df87bb605b72dda3862a1abff4b7f66433e7e04f012bf2a65a6f7c5020cb11259ecc6b103b601f2b85675c8f046456253d410e4c49b7ce6a499e59c14eb3eea8fe3dda280af6819ac8bc2e1a5ef3f395b56fd875ed46801477366f99d34cdfe6114793fec3ef1a4d1bbadf052f81a78bc2a93f26d314b4adc54ebf22fbf87de69f2659dea9546cb5820013a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h7f8104117df1f73a64475e3e0564eb07eb8b65a1b6f1ba6345ca309bdb9c79f0180d802725dcc5d5d5f15aeec24100a10643229747290749d5cf46076623d88aa3bbbc7726388fcae82847d5ff6a2b50a37ba0c4b2c80773e9b3bb0f8e74337f0c51be35420c40c1ab2609d26dbeabae1b8c37c3eeeba1288b904976eab9154349d416ffaaa056881a46640fb0d5b8b9a54bf66b1dd719800fd46dfc9af0c25d5fb33f1eba2ba1cecce544b96a40f48c013211720cf953d04c3d016288e6dd9e814c9762f6c7b75d430757ab6e80ab7a2492c2f5715514a705b2f0d0555497d4f056aad2e0a437c11916742b87c9671d7262e42d38c3dc7a9dde3d4feba24fc0e3ec86cf9eff73d918f84c87980bad8265a2136481a778a01966f80fc5aaf5d0f3dea5cadaef7dbb5d6b24407226cce6012b11bd9d273aa1fa4d022b7209821c6b945db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9825692ddd121180d2ffd3abb823c2a0949f8285537a722eb5e5731629b1046de7cce005279fd9a828c3d23208e200aa171cd2648a6327a97af6fabc9259651a7ec6fa64ae6a74ae8f3e0cebf3017dd94898dbf70e85284c9e7a1f9b1224a51e432599f272cf826a35ab848adf19cbcae72483881c7cce0f5c0a782ba3f56f0f8c4249ff9dd5218c38461b2577ce43edca7fe21c1d3057c896407ca42715e064e87b0fe0f2adfea15575903618d7378150caa67e591560645d6609ec0d358ca5d09d37f36f0cf0a4b2f19cda38383c85e5f7ca66d2c97228934b5d314b89bc438690a2318ff66afd54588195387611c6219334e9c1eb5edc2a12b7c503d54728e2da44c66b67b249bf6396b658acbc2af293c42a3294f090a733260a1e7bddba185aef3e8978c0f07308fff49dd4b279d342690a1c37fdc4c23051b4b62fa18fea51dc1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h7152ca1d766b8f55418fd40b5f59c61f909c871529d66c12bc195fb1365e114d986175929f8ad77afdeac54f7eb3495b4c6f8a4dc340eb6a1ac94ffd1d68f0710440fc85c70eac4b2bf39a27e5fce581d7f7b6d095321f8b06adf8615c438cf68a9e86505b0c3e550912e11a1d95e82707eaf672ab9d4ef96604d978f09f43219d51e0762f00f040bf9702a8536af9af610f24d668d2865b59bd192cec2e9faf4b31c76567ffb8894f1d1f42ff01b19a3170070cb114314f45921e296f5f9ab3cab8b9839071285477066286f8434eb1a79c309f6eb096204d03abe0b784f9e083d14f5789923a29822eef7ca0b98cd47b3b2c7128836ca0eddf0a087ffbe111729893ef2b49873ca5450bcb690245602b7536e1fea370a4cb2ae28fba9d2765a656f8de21b12b7c186d930c4d724f9a5d3971f167f103ce5df6e9299598bfd893215e12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'haad5e032ba20a014748fbda4023be7b6a6ae9f22862581e26b0556f282af57c33a09419662a4d7c9c49f0569e30a1129ca889b0f544da36474219a118938321e438fd20fe10cffe0d846b2b309a4c7015097577fa3b299e3512f01bf4385af25e2dc46b9b40004dcd6a3da192a1e399cda8f6f0083d3127804feb04490f7aec79c9d6a9b9432be4d8452c48e32d2c7bcdf120f53cf7f90ba75b09ac0cbfc8e8cbff2e83ec6b95ba6b390cf7c0a74ad4d1286c8864030bf6c9e1ab3a40b7f20c9546bc022704d0f42bf5a7f326c533bedeb000c0f31f614764bdeb4b89b0538d778d59dc3a1f43c6a9770de4d30b1b68f623b806215203548e091213eac23055038f57580e585622c9226348e2ac40edbc7fd868e5f176ccadabec4f2274ed5b4445c2d0206c699caabedde99f5045cdd2bfb889b5d4ebabdd2bf66926764cbf158caa66e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h142d4b6991af38653f04071d831e0c4799a0d140a3b31fa3b9b9f22262078e219a0f25c3bb53c9117b663b905bf269a8b21eacebc060d0d8ea0ea7d9e85dab223097eff2a4807ba6d86cb42e71dbe6f9e9a4217497598db2ef4f82bd56230276c1950965a64d3761f34745101768de0919642b86d721c56cf5d17fd12eed6201f357ea30ab3e7053e68a0b92fbe894807b766ea49a6113d515c7531eba6b537acdfcd300f12f089bd8cfaa9499cb9057b79b1feab6502c6925ab2bfd59ec9375f5f7e127e61613f089e3635fd55c41fcbb5844398b950aed9e8958232f1b0274b98d5868a80c9c5448dc55562f5be043e0d5297d17a6a1a7ca416e7b474935151cfda6874dd6d2e6c82a215f26a7229e07a36e418d6fecaf4185c1860b8eb4434e1574b7ef1551da7c2b9cba584a81372566b908daff49d263de32bccddad6d6e1481826;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha5fc16f0cab074aa05e828f1fab074fc813f87a200044a3d5ea7c0b272b8de0cbeacea33b2cde8b58d93fea809036e6e4656e8d20b472ca5b34a0d5c43edaabe35686a51c8cd5afa35946427955a1a0607581596196879c9f884970dc5c3f7023f8f2bdc2adb8c90f68b8332829742600886a5d6d868f70a1423514b41a1db0da7b70a99bbd63f673dbee6119e288ec0df5807361bebab51173a1664d19bcb20004b6562c064cd3991e3559e327a782a429c8222ddff9b4529019bf545728a417c3a71a09437cf20071838ba00cc59ea6c1752a963c502717433a64fa5cd65a7c483f56ca9a700ce06bd28a524e822000af2bdce684575d53a8244c14a1d0b8b5e9d31de9993a57d3b7b1d3a855ad49e52c810dc55856d8a109854d48adf75199dff6fd0b0fbeccf6e2744f305762b03c9d8c42a3278ee10445345c59aa44f113e7f2291;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd61e95e35327fda7c4f46747e465df4d3b75ffa99e6663ca0a099ca97d4fa72c393def787afe3180a154c4b6560a2921f6d8755144efe7c781c3f691772e42d1106a143127eafc642bdb48afc61d4810c0173a20a6223dc2c38c2ff269ee4c4907aafc544e2293ee66eeab9602ed8e144de134fb80a80a6bc209b1fc871cc8a643a8d432e8272d46fcf356675af3e6e9f6011d78d40d985b8713c21b17de142244e79d47f20a888ea6e34e99fc40096bee40670dff0a12222a8d270c354c50ab1cf9f4f3c6c4ed670ff88f7f47c48baaf7f67951615cf484bdc6556e8e9a84ba5cdf4b55eeae5b6e57d58004d0b039ff84f22efb06a50e71051c694acdfe6044edba6cf1e1d1cf3b47d05e837c2e142e7fd3ee01183e46d20bced53d365ea0282a7d497a5c55e69488de94126d24f3038613edeae93af8df913511e9fe34d33bd91c9c73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8e137ccc1e3c44eaa4a5c7e3ddc7e54b00268ce1458404a5de677d1d7a83cde4153fcc707e86c38c6988b0cebc2bd3602aa5a97934a8efa4ec72da6a61ce0fef3f8ec654724633923f04b3ab1276e6d549dd072b6f82c4087636b3cf25a09211ddf92595195eed57f0e42054917c6ee3c1dbcc1d159fa437ea2844ef6a36300f2b0a9c277ceb8ca0325274dd64a45c3b1dd5f12869b7f8aad0fcf9f45dbbcefe781a9b45c61b12fe3c63191ea9d269d5cb614135ca9fe74ffd9ca17feb8930b8bcd977614cf76ec9ecfddd3f3421fc9c3a6d783b1b9a8a6c8d8e0627f0c20025bd58fc337e09b99a51fbae0f57b32f4f09fd784be5707c1ed2bb7384712fd26b61ad733c4be7a659be76ac1c01d965e5d17a91d4f3bc5e67edb205f22172cf1026d96417a57dc093a6a4de28ac5718d75f2b27f6e2eb96739988423468a742d6c7390a81;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc62c810b50103579af27de9efaf096044f6e2914e7c913df1fe58028cd36f7e53139e7a308b1d38e08c5aecef92f3a626f2358c7726a63fbc87cf0f9575e32a99555e1991fff0676e2af3e0b5cab2450e67ae33f8757fb84035912e346b6f8bce0baa9f531423d303a8a7c771cd4589d9a4888340f10850dc8916e587b2edfc10fec4e40415dfd6d7789b5d3ee3f486771793794e6d315f5390c78ac293143d733e8bff036b2d68f5c574d89d0392531c8a797860e3892b2b3484ca5b9325b8ffeadd42c30607f85f1b6b796d62b7a89d83c30c54b369e77940dcca9de30ff7fe25a80c507ff4a7da53fe3b6a7a81964bf22b18b13430e91d2482261fccf3c7a9394d67c3a570f8d091515c849c8736cbafcd8e68188912b35ea4b2adbc113c6625b9d9c280e976361b45ef4cc1dd510cd78a641d08e3cbddbad7d2168ee17e6fb258ee5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h321d3f4fe0a1420d46f5fc68189f8f0174678106a264eff480ee1d717c8d9dc660ddf0b0907770345af0ffa8092a00bda8c701f3f1b211140cebfb963acd9a7be166bc40b764ea1c1c2692e237efeb8908f9ae1868b478ec7d5f6d0dbd87b509e9228254bfec2db7fec898c51a05027b5702824a6463cb62942e9313e3adde663187a51058ee0f6968aba0541b864ea9ce25d5a1f044ad3a944053fa5b0d55532008558f1967ea03f149a9c741d0cc0d3b9e47d115e125d38e67519e1163328f878a08f60cb3f9a70a9021220f05b9b362c3f88be01d9597043d01fedbeecba698e6b79127805bcd4f899ec9ac917a384799c8807bb3d7be1ac8b3f8344867dc2f84672b9424ed0bd8ed9e031fa30ed5652ec9bb1de2f255490cd4f00cc2f622998ef588ba042ed0c87560e063e750a1287f764a0fcb008df143fdad48dc37a68a4756f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h7850c726b55b920a90f6dd5f2778353265cc35c0989fb3d18aec1ef7869ace717dddb76a2afc7274071eb0821c890d59c96fd2573a374b72cc6083e7ff36b198d7998724f3a5b75b7d21476505fe4244e40b76097bd3e94668778824a2ff995b0dc9a9d65f3058d4a1fa1b77c3b0f295247e383ed1c4fbfeba7f77b3b0f98aafdd7836337376ba76cfc485bacdf0e360efbd184be830255118651d3c69d9ec546b3fe496fc9a9ef9d9079ae3016027a29b214e5ac5974e384f219d08e55edf9aeb39d19f25d2ec29d0f97697e188207b25c55b8b89985771ac4c1852e7d3170364cea2e83bcd128fe416654f84db87f399956a1d00c79b9fb74f006b95d823e8ca128edd3c39b1b36d7c41c1103dd16d5b523d33e70c3a35ae3a0fe9a4317d2bc7bce715d81b0d0617e6ce34e0f668e622104df37fc6dad89988ade3a11474b9d322001d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdde6586cab7232c325f7087e35f94d0a81851c06f1bd466d939eafe7f0a9e44ff9b84e022aeefc5ad039640a2b9d38073c7b6853fdb8578ddd5e8ab30bc5c88728e3c977ad8b108b024d02097506b1459d5a24f02c75690c763c1879ad4df5216540fea58c819febc0832eb69c6ef1008f0cdb516bcfce9d8c01838d42927e36259c19f8257a1e189f38a8a651ff0a16c0a21ac4116cc55d1918653a1fe5ecfaf8f15573e0630429e647e576abb9c154e601c84dc200fca560ca7b1b6803f3ebc3fcd4bb39abc8051eab6346ab884f651aa52f1ecc59ea96c2d932278f37d89a3f671a670299cc0dc5e1f74e318b4068a0877f37e4584ede3c31b320acc7c472a098f0647c683078863d804f3d2fa7175025aa39eb434276714eb78222550594fa183b019f87554202c48f59039f9712c5bde5de169b96d6ce75b6ff11e5855b945e85fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hcfa96dbb7291dec47102088d2c504835e6e28d523c8db61c4df458cadcef5bee892cdf58851a679eaa5ff656d54b6f9808c0dfd990591b39f19f6575e4d863ff111669673b90b9c28e468478e12e6bdfd182731c0637a29c5fe1e2832607e441160095c6db9f1b916748950a7690a845855169507e96e1f47294d9c82ce6e66b4db7e683568c5b270007950ac3c0373c38563565b3da7b1812065897ff5395ad2fdd74d3e74be526034aa8d00ec53bcbd9bdd59527f28e3855623e169eb94c900d2b0c28d9651482f5319418d29739b784b191fdc20880878533f29e5cf1ebc227379f65634257052d21a9021b7601cf26f1e0f841bcb0ddf48e139800ab231371037fb098095409ecbef88f269e668f0b6873f757b609b27c08f2ed79289e76f420da6f6d9657a3b59745e00159f637057ec3202806ed9d648896d4ae70b0b7046f15bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6db9ddadf52af349f342dbeda4e03f03e8068020ae5c7b637e029b426d505a5aaaadd7a2d78d6467aa837f8639d80f0dd2383e9092c87c3970da45ff86149205344ea5041ce5a98150838a6b70bc77ee4711daf49518ed403218c02aae73fbcd83087ae1ec950e64e8af2f321952dbeba04f9c6940e70c75e1b0b31ba0a0774e35c1831ad959d55d8c628a9750e25b262bab48a1ca6b8ad3c361ba1b2913f6a8ee9c7e3a64cb98a474dfc12d523068474daaea3df0aaeb24357b20111d73a7a0b4717c6e14ee6f85e26e174de11e315b4c4ca2ad968ec9ba8a3b0f6d33e8e840d1bc79e413001f96865c2cc1831b8c394fbd1f24d99a1fef6c397b5d90f46afb59039b1e9c1956ad15890f1bee167314a16733f2c00eeb2d3595883706d080308cc74e5ae7adff22cfe744af84f1c20a5b3172b58af35b41866d904a0632c195cc3f565;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hbcef99968c1990ab30dee9990e82a503a4e61a8301fe9e3e542c2b9e567cbe3dc51afbcac9dfa961083e7e273b79f1285cbdd29bc1be1b6affe83ecd14c29be198bba9cae0440d0b8e12d5e68eebcecb128a3861c0b75dd9283bc9d420fb74b7d2e16c4f0c56e6f2dd16c2070cc0070c8e3cddbe2a9d1a3743870fdce92b49c4dac1729b8f7cfd4edb299085b23da1ec15e6da2ccadf32ad7f3d2493407087a9a1405e33f02ce8461e775c24ae0d12c7e3f661b29afc6881b3a160f1f3f2864337030b2a4b0c47c93616f02ac8ed62185a33da432e53f6ccdafea43b46a280ea2d02af17ee249c6c91c695e49e6bf275ef90a8dd8e82d36bcf4c2d5702bc32538d55b758d5c913b38e5ac7c2d40af09d509f54c1c3dbb5d4c3cfc9ab7f20c3a7df0fc7cee39ffa1bc9c1a99f48c7732adcd8e1be793015a0ad556315bb1c9e5729f8d3b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc6209a5db2a54438a2132a59bfb38c4f638c80d3face9b3728a92b2105af9f4e81135e3f6bff0414b272554def1659c1ceb8e2acc9bc4cd66257e5181a8a6c2f3f7c2010688bda033ee5c478110359cf10151e0f7db745c38ed064318c3eef82cecd718143a935c3af3224dd23ae2629fddc4ebcb7d5a81b8f41ff99163c8e0b721eb84bd3c6c172092abc7ad0e83c24502b9ecfaa580761fe02d05ecc58bc1f5fa7146335c2fda62114a9ac17c97dbc6b2a70fce0926e6ce426062a6a80ee5fb6e0a50929a83dc26b34463556dc313620d2692afa30b20c74828de81763c8bcf568ac0c5602da33472ab28ae1f90f5d7392b8dfe5474bd80a1842b0cfe5833c5357662682458f32587a024fca75ccb2d488e01e1803b0e8a0f621918d2ce085ebecc757d99d31bfd3f946c4381903b2477cba9209294c1117ed69e01d6ef27df4f67e3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6a15494c39a407428acfc7f892c7151802e8f950c2363c063e856058945990600366175e73dfba4ef28df1e4a20ccd3a4a86600d3e1b20c12d04a7f0e5588f06a4bad02480fc2d8a08454486e01a1c2120b52f829e3b045194b7af5fec3c4acc8441725212e03b46ed4219fc0191489a5a9ed98b53686a1af4058fb96bf8a486636bba800a973553bc650e9cafb323277912d0b253ac40628f0bdb65fc909b4915cdc902cf46380b71149af1d43fa55b27c431716460f6a4e940fe183407e5da8e224c678beb00ad67412a6493fc34836563419393df0efe7a265ea7c7608866d8830e11ac05e3e154d62d0b606eaf1e892071f79f00d1145ca9decf7e64dd5e6831a72bc24c0b62d3bb9d0b1bddc6d6392a8f7489025ad97d6a41f4a629b5c2f89afc92cc279f97b96172389ed4328c2f363e4df0412afb4ade25bdfe68be16c1dadd3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf69b33acdf474f828677b8b5d921dfc533a90b49113c9c5c66d7ff810b60fb80fe5db08fe5bd3937ab791c321e4e43f38942b33733150c8ef0a998a2790960026cd111d15975803cce1a3fc3996dfc867d7fdd64d8f38554826a4a7651ebe37b6c25a1fd76eae5f077a21547d2648dfd636d6a6de18e2aa3e6a57e506242ae56846e32da51d623ac46285eea479af3cab4dc6952beec0bd9572b80b2b630623860f398c92a4f9aa85d8aa48409fcaf1d1a3871dc55300154897149bc6e10e9e879365da978cb07d29a598afd7c5763b2a73287b9693145773d8b6728318e44e8e42deb62ce6a929e0907b85ed4e05e6cc006396bb2af0f1d3fd2d4c81e38f1b154e5d8acd5c5a7079d62c9c112461472033a507f89ec5077b1f86e75c6289783025716a9c7db874a53ddab7a86c44d0178215655e0d3583e5b069326935a334e1094dfa7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3119d024c56a47fe9b8a8eea801e07167f22059bbe9d72aa2acaf1e40c7b0be6bcafeb311fbd414d08808a433b7effa8dc84ff56ec14933c49aa73288b12a4877a237bc8103dd1a1aff1d2316c241366c709113cafa100bc03cd48af6153945e4730ad0f46011976cac4d035665645ec3e807f6131ef821d3c085e8808ab78a0042647f95bf222d0ae1419b9b488dd22083856b37980184f8bdad8ab5c4b386bfc1d377f630cef36a459c31383174df19a950783e3326e61026d4dd41f7a1e6fd7e530ae90f978ea9b46396fe7b167b1c590efc3f19abaae6e4b92e28ec71966cf12fcb5f1de106bc3cb3fe2aeb44bab123c8eccfd7626f773c6696b6fc12a28de55588b589aa13930d59ca28e681b6c511a3319b53213f01c6ad2d15acf402f43ab1b66dc1defc5dfae1c68bbf70f27f6621e3a116f12d6410772fe990eb08341d7d5c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfe69fc39ca208e3f2fb2e190237ccfae5d1833bebdc0204c05d5a3a9b13d66d423bbc35ddaee9940da0d3aa39be4177825d24822123bb1e0b2793f40f9d6d46c10971b3a993438502b9e43c711cc2de2083bebcb107a85c66142bbf85ce41566c3ddb26c309cada8a599e681353a1722dc97495d277be63f72f6d084de967fdf4666b6cfb67c26d4eb37330a265a51df15e16fecc8cc5f4844312a5e8fafb13585112a6b048675fbe7bdec799381e65018c76ad6e06d956a383b73d996419a659b4c348f6b4c138e4c81aa4a82d3208b805b1ade588d722dcc725631bf81f5bfa1734052e9acaa141f1f268664624e2ea1edf479ed24de5f2bd852104aa0be6278ee045aec32a5de8ef7fbc9507cc78ef828cb8e6423382c4e749b00f144bdf335f7cf46b96b1cac15d89512ceaec96e693f5a640454befce2d46af1a413150a638fd9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd1829a473e1b12fa05afc0f140ace9093ded864f00489edd553afb4a2330c01d571481af42f37100e610a86962b8c5b75df06bf3db43922998b1d838974ee7a4db4140a880f1acd5d3cda5584a69c3e7b3cab713cd4b48c425bf2513bb7dad9f0759af14bb6863bc310d6267aa134117106204466bb01cc36353c865245c12cdd9123d70a32a9c6be2e1dbbaf08fcd4d312c40f4a48645bd3ada351b069204562bc5c7f75182dfc19b4e3d6c2bbfde84a81312f01de8cdff7121a6643430c24b08866d0884d5369816d96225e346cb814f171da75fc37d008fb0573b01f6e30b429ba4c69177a6d0ee103b600c1a68b6e429e91e5458427f32a4daea2d882169da3f44e09364dfb933d6fa0c24418a1628ca576916471b4455f2001ad85eeadf9b1352818bf79f81c4eb4606a990eda1be69ae21d31ed605c56d6a794cf5ee2f0f6b7dcf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc0c7d52a13200b244ba6e618de962b09e32922181b65d2d607b91001c73556daa25ae00b8cfb44b8725bf50ac74533e908749e7e35a96fdf18ac4515412532bd6b62b7271180b8299456f85ddc0d730e5eeefc91d0b0b3bc99927a9b0ef84c813ed3340fdff08e9be4ec98ea7908271001fbab1a289967989d9809c36ea34a69e82e387490154c9c741d1ff36686da3536c7618d4b10276a3f720289e060b07135d9db19bad183c4c832587cef186c8cbc13eb80d92c4faa2b8d492619d2f6c288683285a31f91482fb834f31da622def9242c676080a2ab589d5f8c8d7c05069beab80c16ac1a76fd6a4941214934b63ce7dd8b5c181d801b39e4cc9f0d71184fd4921e3d4d806a514d189e5430c4e24718acbf118e7d0ec1cb02758ac49dc7226e58e4e69024c7ad3296cd2d17bad60b281ee722b603b096eed75fa91968ebb99871d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he9344f756441dc477883ba35f9e50cd6c0a7d70f5eb5b1459d9622dfaa9d8e6f334712a19f4456f49d2f2b30eb237ebb492818f9dd0b044715e1b0c227829f81adae729bcb68970a2bcb1162a19c155327098760ba87770877766be0da22459244c96f74c85f914b087f96a8906962e281a9d62fe7a9591f2dd942f0922d99d219d80b79285691a3ef5441f8fc53414bd7f63c5faf86ebebc5dfb89311c668fc35c681f1cba4aa36afc3b6de82356a6a8fc78afdb4f20218cbad96b2a20d8e3bd0acb8c8e727a34f792764090d566d3f03fa5b24b2f2ae28abe9e270825aaecc15ff492ac256fc02f0cf99345e1483ebbd9bb964800f26125bec3c13731757578e93c05df05371ec3d250f983efbe4da3a6492eed1d036265590aec4a9b232cfbb6a34ebf4d9d0bacd9fddd838fd0a50c26650cb96d3e77f50d9d1d9401b7955b3d62e4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h51979a9795be7688bec36201d104ad1350fe926a30ea90074ade21f5f7827b8e680553076e8f6859073f4e77d7c5e84d346d1e9b594dd47362deca3cb07f93806788b5bf2c2ac8b3af537a7b3b51744004a6c5f7c14a2843d3aef38092c85345c485ab9e015b98ef4161ae466f6b3662fe964bb64128efa3c0339f9f0840662a64e70f4868808c62db9eb2d41456dda85c6c104a5d8c351a0fd1f106959b83efc89306b879d58ec56a0337020bf3004b7405bb26fe52f2d8af55157117a4938d9447e34ce050933202e5ebfe3833aea5951f830621320ad7361b663adf078f4d8fcd257c0f9211e82bb9df9849adcea98d967c8f76b3a8a2422984de0a3c368f7c45adf07e8571c92cea6bdd89abba97a55bcbd0380e535d8850b3e03a2fc87610d6b814607e9de012c9ac52766750c701d5e231d2cc48a76e34adf5a979be72aa146c0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h92e00767f1c2acd1900db28a3b3424d2497bd69226f6c490e39f9ccb6fb548298c82f092c77861c48dd5ff52b2e86950b34b3278f97852b28a5a6b472b75e91b44f1a0a09bf4d2019395ac2c5ae79c2c1ddcc9b273234d246b1b22e002a613cb04bb865f2723a0e6f366ae234a3d4076bbd163e5be3e169180f7016aef8ec1938ac762efaf78ea52058ed0b24653eb23f5a2fe7271c1948a2a4405157af322093a7386dc4384676568143d4e3784014ff9731f797b707ead87943b7520088c38401bfde21d50fbedefb1f5f2983720f798659368c0a8f1c9440665710142424701256cc73a8507f76ac7a1b8e1ef3e86274a643ab78ba7225df63b4d6bff917c292aae3228985940eb9667ee3bd95bcaa71c7f09dfc25af09e7b3f460151c0d089ac37feb4c91eaabd1570da866a70f180c5fcc37291269d9845d9f78c9b84b73ea8a7b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf9838f884f3ebffbbf3ff0de7ec94e9e541680fc1eb2ef031f9d9fe45d14364b75fffa2b174d04f58960fb45a4268e979696575abc7ab1148a78e286be3080b73dcd45e2af5ad2c61dcd08e81625a987aefa3daf82f7d5cf660182e98904b1eb6ef0f1f0d95acedd1ccddd54af8a45b2d84b2526dfc9383802707536f30198930791febc85e48d217d62a6307f04e298889900c7438ac8d7333628fe0f1f6452e5538424b444b8cf4a14b8acca8cb9aa022192fd75e29ce179d128b9116e5f0bc162934a5418c8e082329a8251de575a20910b98edf9aafdb78bf85d77ab44cc018d66f3f1b0fc362174d1e772994361f9b58a9dc368ddbe07edfcd2adafbc1d799d7f0f18cca544d8b9f25ab7d08fe1aeee21aaa79b3c77e1df8b9066d9eb612018a1ad838aec5deec37be5678d5f733e321a3c2c077f0dd0428cd087ba7f5b55c8b61f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8abf45ef7dbcc37e69e966a92a12dbabe43d0879de3d70cd42012e2de69c675c36a5aea60e3aa55857a275c7e730add2396e2d31d69e116829fcf10fbe987dfc328ba4867b1e22f215b31b002767dd5f754830f1170c5b0739664cafa3c6d98b9c4010244692fd3483456093249f7ef4886e5fc1b88b61ee993a4ddca8b211232924e839828e841af5dcb8622a243b60c8b9bf33161b2c3a04c92a1f4adeed7ac92132d80380ef595a29280ee2ee49b495906a8be9c0eb487a91dc34354229ee2a4c2b059f9114357c87ed59b4fec0a11cd59b2c0822fc1f83d1c4f088ea338ed234553d54ac4eb0bfcd66e5f7e7dc537206d11af81dcf20a61c17e1af7926c20b395ae4452a71d3a5c738d35e959e11e840a5fe2ce0f811219478c509f6d0171617c02a1d6c8bcb59283369da56fc886c9f8d6d8fe29c80b811ea440ae1aac4c9eb671a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf85024de5ae7cf65e27aca22e53544c01f3dc304f29969880a984b8acbfa0d38dc2abdf209a60a4616d27b7d89235265bc965ff12a42dc3ff19a013b17bb92b1c34dc2de13fd595074aa41b4ef07b279bb71e45c20e926a4f997ceb53ababa37fd45fb7130f1dd1349abea3e7df25ff41b753cf10bf13ebd0fdfbecc9d0a9fd1813e819300dc3f7a373879630c9a90b9d5f8845c483720d7993a92e6dd7c428ecae25479e836911324054bb145fa2cf230e1eea63e0341aaf2b643df1a75fdd19fd8b8d13e8e7e0cea26e611460b6d5d2d2e4c1403583ed6c43dfa65849cf463250cfcb4097ba37990e6496b451e8bd5d494ddddc27608fd0665a00de66308b71158cecb03b4a873e86b4b32c0251cf25d21b4575c2f600ddf0451be688ec7e955f8e39be4e8fe438340ee21662ff212cf73537090870aae0015586afc3761c04606b154;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb4a060cfaa1bb9a90f8ee20d554616c858b724b7590b17e3bffc79795559b42d535ad39096904932c788c967309884912703914990a4030615676b1a4a471211a0bd52189ac76e2fcfcdf98b835ee20a1802fa3fa532d62a888488ef27ab0464d61af1b80d4ad3d4d1c23e68745623a8901b6364c3e6b66c2a207ba66acf20c109134fb0e99f5c62e494c42ad79d51a4c8581e3c9c1ed3bd1692e171a7589d5ec110ca20f596821c71bda34acb92fc62fd621096949597c385f72de7f2148792759f72b94a251a422efe3bd5c6fcbc7ed4e7fd4f1b351dd157bf8a1f259d820bb1576487383dd92fc1cc0536a9a543668484c4e6b6dfb8304e12f97d6786bc11b7fce21b9096ad994daef69532c841a812ad39c93da1732081ece7ce58f8b2f92676f482ca99ed21812baed25ad3cbf59b732cca4b5e49d7148938dcaca517a3503f6b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h94e69694788532119737a511bfbfb6952757702a1d22b0e60f9598cfe73bff25db2ec0c0cf7e0bcfa9f6a07aaa3328a12d78275ae4bb8246a038fcfd5a5253144e81b43872e489d1c33e337fd45eec2a6bb74fd269943f9584655ffa9581c54a150ec05451db0b5c2c6968aabff449a070cbe6ea1958a6e7549c7bf0a9427238932f4bc4081ba7ef875ef898f2fed30becd857d64e8c637a4c9c7e3b5d95be0425b04dee6782e6e1540c7ea8024e9f3d54fc48ded3b0eba4dbe97aa1d5d0d800066fa6ebd5570adaf7a37af86cb2908fd55e15fc80a3e2ae083c75969a34366e74b284955e10ef5df68101610310efd192829ffc08b69103351a2cba8ea2b27cec5dbc1454ca6d814407d3ce362dc8564ef4299708e1f88ed14c596a9b1ee2e2567f71c94afebff8c533422bee425e0a2a9fb3aa4e3e9483e16c298ea6bb93f0f0de400a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hce29a46069ab777613a4ce7217b38dd388082735c0c068f5e461c9ac0b45014f3fb713edbdc5365dc20aa88418dd74317bfbf9e3f27d65821a5d3de7a3ff677608ba18601ba6f11ad7794328c99f11704f62c3290e44c4cc85ce30bd92550d9a66b91ec3b8f4a1ec1cb0892f76712e4b7c2f2a56e73028885aa57a9140c75bc8e104944a430768d6e3d5ee84609730a0f114977ebe9a45f0db9530c8123797e71eef9f17e88d599d09ae180621ce9dc944d3eeb4483e7a21b2534ba5e3d8264f4cec030510801b4e0c3df1c84acf7ecab969ea30b77ce5fb318a678732bc29940b25dc21ee19600fe13e12223a6b1b09bb9d181c31b1b912a27d054f6adbcf5bb3ce0ec767921bd01189c0ae321aae7cf288e81b78e702062993debc9414bcdb6f0b1b430031ec2a8c2f637aa189d49e14dc818da8e5bec791d749fe0efcd85bda3cc617;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3f1cef041cc0ca7fcfaf35be14c244d96a83c07deb076897339ecdf3e69773a7e35a45a038da0849baa7ea27ee7f0084dbf3575642b01c6bc4de476c7ddf6eacf836f59cd1ec6d9bae4295912c9370d0a12ffea65a8bd558d9f80b6d0ac646c777e22ed1d3d4f6bd5c7c36ef3c857c273c3bd36f51f2e12f2c66f9068d12fbf730d7f3f47019c8778fbf73a9714b4de5c04d251bb28cbb023e7437cc3b6ebe36ef437a1f8841d2655b2fb9ca4e478ed94c60aab9af4859ccc828ae69ceffa5926a96f3ba23b903b6340b729eb22ce56933631de5b4a27819d552881fa2edb59740197ba008af37c8dcb4d28514144381f0bc5e73ce434177b4f46e88239d5d9bc9408ed2bbd64b453a60b5c11004fe93c38a6da5350e7586216e3c30f0a37e6b7fed0839d4865f2d5781f62576744e7e4f86aa2f87ea37d8b5eaa700ff438eaac4dd490a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h11bc1f8d0c4a952568bd163c4a48209499eaab5148e265be9b8ee507cdb59ffa912101af99a5d90bb4dac2584d89b874ce9cbebe18c71c1cf3016798f9305f71d70448a862296db4efb368f50829688591d160a688d6f814cdd1622810da8c6148f5c626a98122373847f259ac55470e7d2aad82f915a66db8f66df42ff0530d05fe398f2cfd376074391429e231cb4ad5d28ad3c2f8c1ab5a432cbae47fd4ffd305aa1b74e61aa69289e95fc8d5d806b65476a08d1898d5459bc0e5ae91ba92c7e7fa6e7d13a9d553c7ab8e2b9d6e274a0e1fb6f17bf518506a9c28ab005f01885d0cc24f9141a1a08c0015ac4d53f2c8dbcd7304bdfe92ee33df0b107a3eebbc647d91157cb9a31a325057d6c2a1d6e4d70ab559a8942226c2fab73cc48887a7be5088476a902a7b57cb70990be7ea6ac148e675bcf561745488dca39025c862bf2727;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5de3308128ebd3421307c5c564b1f102abf4fdd0ce422e1a5cde8bd0a265b05c5351c9951c285324f9d453d400c43405d6516c3d511b99c6f94554aa67897d3f5971d8c490d2b4862e0143d941901541237b0dde1ba3bb75ee6548bd0e240e385bb500cbee216a4ddadeff2a3fa623f44e0e7857f71ef8c3231df139b32197c9b575c4af8514b2496d13a6e2499dff2c7bfba890b4d8bb23e1cf13cae422fdfe559bd68c0f443a340cdd5d192d48f7fb6c0ad51f60d887371a9b8d993daf86bf06febd066603afe6f60b86c8559aab63116ca6f48a9109df55e61fe3086b80d331c2d3be3ab8a813fcc9fd11ae644202d49f0be2c12e8201f6c6baf3681f0781aae4c5cda197735cf148b27f4894730480e24aea5dc5f1a936899451a84c713164ff430dc5021b267de0ae74d91b4385d28fc951a6c67b125cb5574f6c184e6bcf8f372e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc7c511019ce94f999a07e690d95fed100f1135cc867bae4faf6058980845277a0c3a722f4f19fafbba59389c9099ddd647aeda0ab27643eb1a464b9b2fcb8cad2a16ea926a357d55364a7f3901ed78e1c84813011568e6ab3ebfa329f97a1212030dfc06530f28869ab81a13c341c0f6778a9f147dc72b6df21659c5c3af2d55a403d7d15b9e1a205554574f2d6271045ffc6e92f2c7cefabecb17b5cb4ee289387c57cdc9a31a05a1cde05445c49f9d9581196fce8e6cf09f00175af32696a5555337d491141455592e8a734eac7ca23691bfaaaaa1367fe49ac28315e5ca707a3ea894c51d35411656d2cb9ab18287ea861a266ec07f3974d1b83fa2d189fcb90548fca363d522c4e321273c3864cfb074da30e7f7bbea619753824420ccb8af6a9194679d23622cd780ea3a86e5194a8392405fb59f4769379b086532f851b4e49c6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha2d852633e288489c619d85400a6a232f839162e2f89fb795b827bac61aa49f421638a6ab00425388cbd25bdd8ce3fc4bc7782874f772a5a4d091ea5d4c8a9cd71d978ed3a3f541432d54d4a27bd3eb1b41c7c27f01d1e61cc17e07ffe16a93f5ac2fe2677d1f6b85285e0e7e2a96c1f03e61cd9e67458d4cb9288b3a1569f1348a713442009492ff290d34e6f5ce069f127f361e5885ceaf48761e1daa9a1019c003c5a3036556492bf4c3d52c131129eefd38f7e2670a15dac8220d621c91a0b97e769122c14e4a87cc87cf045d3ab3e3b7137cfa650e75d8d4ef495cf6b176e0f462af1e4f1717b57eedc4c847a1088da174d2b8e16d001b1db1b797e8e7e52e495da99839fe0c796fba8a39b8d28fce6f3f50d97c7c155c07b91c62a880499dc1e184762d7998cc08de7f4d95c6e9295b92a3a9c8aa5fce4b9c36efc9325cade3a90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2cf701dbda09a1de53d43218300e5046d9de288735b7c050dc350c0efd685008a682d7ce1cd76b7dd43008f9c7ef8ba9a8a8272e2bee787ecf4d52033cd9455d15fd14891a769d093357d6433d2d3e616d7d78d971d15676b6ab47d09980a29e78d008b3168916b083b76df1fbd12c01ae034b3491b2bb053a31a1236ece737b016b32663047e29e6857c4d7526111d098b42b78bca153ef98896861ce571edd56dff3c5f446871b744897bc7fac317c0af5212f73e18b1b0ec989a93f2890ac158a637d0bd44527803fafce766758ba19c45ce7347b55140fdc3e1f69079fc769305e4367fbafc739a4a798c0c00923a74c95dab8dc32a884e3fd795eba5c1199bfd5e254bed93be3814f9782e4161ad99db21b9d816440fa22666ce06eaf273efe5e787852264d33d94b734631f34f8f7a56b2c31be108d97157e1481991a555b8a469;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha8c8aa722647604ccaf63c8200fd405cc308063585ad61de89c169538ad96bceb88f31d4b04aabaa3d7abad9da7c18dd462567d2f74c80b7f1e538e129e617ab32d09164d74f9fc952828f7e5620a128641a878b14ba3094df80f56a70eefc1396c4b4e9b9245667dd24825119458a019299f2c299fd77339e76b0ef27c38d6a0ec4e40064f620cc7fe5e9d0644afd4d0b7e2ac96b74e3d3c6c0bff305412b05c176c70b68920df0ad83c0659e92c3a4666fc415cb17b1aae8e1d753162b5e3bf6228b6eeb88a1df2b1ad370630d1acf6452717241e57833e01383a40e73e99158d5471500170fec51ec8bdc450400c460e4c0e63a7e8e02c0f0c729c64791ddbaa736d58418cec13299cc190063f21b95d96a615a781d74a2d922b0fc46b958ea3fc59a33b7b1a1546bd535db52e3da352584eafecc805f9bfad299ef14f64c630ad8a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h186779206bd3508966e12846514faea02c79eed237c738887ee24212d361df18e8f9f31fe15a13f0ce30340a3fdd9f153deb1450455f16421b575d239d15c064c28d82a8cb98dbae5015bd485ae56a61160a439848dd6682d6caafb2753d56c9d137a68fa0d7bb66aaeb8eeea74c8eaadf736243d15750705e252b9771178c757d9cfd8d885be521e4045ce1cf87f8ffd7c70d480f4dfcb3a64294ff3d5e21154392b6e9db9e34cc6680ffc8bd4556d909da84f327108b483b9c7107fe39161dbdf58f551656cc93e8770e25ad04a53cff8797ad686b0914d97fb4369c08c98017361a9a854c19e5d6c1a900b81fe9171ba2ade6b04e9c87fe02ac14e4fc1547da5b6116159a1a637beb89bb67d76d42c1482ab9ba83661183ee58a430cd84f3f405ddb548b40d4ae9d3a761efd22bff173a5b1e4276b88f375a06885b111e101b636352;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfaaf5d2d685996cbf2516aec16ea33bba97e710765867829c6b99a55a51c7c3587f08c7b4e64dbce60592b332a69c090d5eb6d5ba21a218848f692344ad87953aa87216c81302dbc14ff0363a4c62650f437b0af11bc8a851f737f3b99cc62882312faad8d96df025a2bdaa6acbca4e3e097ba7e66b46984e02f8e84d6914ceef53229307c0bdacdd9fc5df400c5608d76dd15ab8ec6ba27d295d565e9df36dae40429c90d94d29817f07c75e1c681ed522aef2429221c4664a95ccf77294ed18a1f750baa5bc7db0b40476c7e246672ca291e7665b7c453cec3de0a5b1eed5cb39e5ccd607e68bb8560274634a155d2e2889d29c8d60bc572ce6b080177be28b2393562f83ea49a481a1f573f672860414ec0605b0bc7b2970184061d3e83f450b7095fb8a64278c2f03ff1173184380da4df7c231f32996623b45301e3c8b6e0c881c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha5af6f359a07701f75e180ffa84f256b83ac17c051f00b2730afe8ef7ebd5a19d6cbc85841fecc8c364daae7380845fec33a0d3765219b8e95c7391924534b8752af287f612e47cfbf86a5adbcc626fa8fba22126b279f252ba5852a4d69f12113bb32f8f2d43d8941042409a8c8c5155b8f3f21003d88d19198600c06582dcb6359953bac863f19372b0f204adc58307c2cd8e5bd8eabe59eac6326ef37349c27aa7728e1499994aee7b30d0b740b07edca04da738d86b768d9a92a3f606a1cfb1d412ba30ac022482774bd9ad43f1b9f1051a8f21f8e3fb95b9b151c415f1607fc8bf76e3ead4d763cb5005419772233f49492bd871b7e94eb3e19a7f10d20a54a9dc95774078211b4551a0e08cbb158ede2d126aa335e33441291de672d4ef35d5ae91ed32c2446f2196d3affd2bb1d40b318df7ba0defa311e618b0e6ff45fcec4b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3ff9e6e23633568960c548f52e00db53a180a35c9b05454f60cebf494c4f645bb7775e3ac6fcf13c5b07d79036fba9fe4c309977fae0e984502a9302026515c401947ee8ddda9db447b48e86641759530abb7bdc6148fe53cbde75c4e4ec304762f6731d7875edf1f97306590b6d32470776c6e5b4eecbad306afdea107206e990ee9821910e9dc9c3f66523afd664e6e877b49576fbf3f4f4a7cc0dc0c624a39cc888064941067b48d388f04445a36a6b7819fc641bd29821a5aab5190ba7056451a35508029f915427b13c279474b5a33d90fc7f3560ba3fd28f5091e36e4701d2b4390ec4363d222a22995d740e401a226b97f72a6b81ab66011402209925120d106387efba4e185ca184901ee3d7b908a3d7b18097e7fd2d99d6b11a3ab9bcec9185a456842fa4a8974a3b56e5e7d0cd3994877d8bab05af5366a3429af9a8c54f23;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf20a38801108b18224f39b65244675d56fa0777e957e646553a72f12c4a91ab31f5917fcf9e05e55cb7850ccebdf4b891dda4b35111daec5d266b7f6927a400450c6aa6c45df2faad38c1dc32f937f6013882003f476efe67079597be2c6f923a56912fdad65497555d3be4851bfe0b02c8630c96b4d6a05866e185cc658e58c356f6d48eee9d209c8f1c777ffdbeb4401b412ffca31d2e10fb28753f0774cfe8a5ecf54e65ef28ed63dd75084ba45b4f8870bef93eb7a1d9a6d441c32154a368e051b1447a4521dc5aab5a3c6c1384e0cd516ef5023afc07d77da6081c9549a65cc2a53120b3a8844d7d09128df2c3884c6b1bf32cb3d2881a5ae010feeb30bb378ebfdc30e3471f2d9992a5a614bbc00f4ea9d69052c179d9824775d2fac56f316275f9cc7f07bfedf99a9b776e4693d58b8302f6ef88c9b8e38618f05b2ce82beda25;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdcda1824024cb3d76df56aa51c1a8f1cc324b3ed670b6643dd59c4c798fb113256e76d8d01716a6357e4b3770f8f1974508e64e7e11a6bec10da1f4f225b9200fedc766383cd84d3494db0b11104fc87f8165479980a56a8ba502fa9de7bda1cf4a86340b2f86c07fe8243537bd0d5c37f7036c57b7f5bd572df54bacf07c599b78cce7125149044c0c7930cd89cf5652818cd730a6f8e6c7925ba98128f1d47c4554c45759295d532d8c1115f50ef88cda035f588c54cdd6545f1c4a541a6dec2af17551b79ad153411f0d4f6c788332111bb652b329369c3ead9696c3b486cb7d6042e937da9b79461ca97a114480b37cd7e1d799a74e055043074e382c538e3b84477ec3062c1ebb51f918ccf8f8b54caba3dd15f4368841505ac5b95c221993fe1d4868a6f836a22e92d689604efbdc7ebb3ce57c11461f417675b71d58f29bb0aa0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he03eadfc23508ca29cb359e0f62e8878a50a6928f4f32ee8ec4b5a85fadc47cd296955d561f734f6f17c4c9de17a5f0ea0c49ccf08534cf18e16daee4603c4c2245bf6db47fb5094c9d8e499513fe8e6945b034258629a7ac2e3c142ac10a82bd704203c1b07df3828765590774c755cf921ae42bc65be670044153bf86966248a69a535bb030c8c69c2fd9032f22cf8c7d15e01a5ee48e365290ae08052eb7213b75f58e809caf3b39c13e1e7372301689741f9d57c5efe319798bcd74330bd57f08087eff9c640955bba2e83d977ce0a79e1e6fe576013099614edf06b885bc283039d32bb4e7f0c48947f35ee1dbf32bb06d20fd786e1b5154f4c0bcfc205e4a2af57764033e8522ae744eb6b4861247658b97fdacf0a49c396c4f1194a11ce7b36f5bc4d3968ac97de5e1680e0c033f1f871a15a06a21965c246fa64b0d316bde965;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h82deb2ee5427cca854b38e20a50971f294d821db414e0ee3c71c0d7f4adca696de8f50a66511cfe9a87bac98a293cfda6ac24a610cf555e4c9c92bb57a422f796e6308911f2e99e93a963b113d9164af57751221e8bb3fdc0441c7977b2e9a9f2dde769efaa56e9715e95ac5041a327829ae3db268acebc1ed222171fb63bbad20676ee3288e06ee75ba770936c1411d15b1523eb2c9cc1270757b90a1f75c9b7498e85ead4b519e9c519fd44de3cf3bfcce8ef3b8f1387070682fd58b7bf8bb89126a6e027e20b93f944d196506d6f42fbba64d0912e474c8e8633fa35c5eba294ea3941b1ecb46f96670fd483de5818a5380907ae5c53a616edcea7cfe2c03528b88bca7577f6c429d7525ef3c4472a6a889795fba72931b2840cfe64ef7f0092aa4fb1120a931e5f1903f1c1ca9a73a7bb3c908f67cae656d612b8757cc2e98b17e8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h342105e08bac22023103a391ec8973059aff6b25ada0c45668fe863d6983358307fcfde21ef95efc51855d031806ee3905d0b280a03f8c24c9fdd53ddf6226ca20320252ade901a4a60fb397663103cc65e04e72c4fc1ab2e429d9749ca54a899f42570c5a0129fe5f7f7f6d0cd5b34ad14bee94354ea4147dff840f225705819c60869fba0286c992d8d99d8520ab23807ac29534eee558a2e5467ceb61e750549b2e39509ce7da75972cf981661c1189ef652c7f8739a364c0d999221b3cdbd5833b641c4cf665a8c31fed6ac74b3e4558a830fbae61fc8c4d3cfe979a3ded3fb8b6f0c53bde5a29c4fe61ad2db638a2c0ef32c1c172658a51a81c1077b12546f2ce8327f960bc3e2ee9ab900c334649c4a457f0a24cd998890e32685106256c8dd3dafdab74f552acc013b823aee46f4033ac860df37f1af7717cb60bbea1ea0e952a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h94ae6e02a0f60f03ffb3273622ae65eadc4a0f37cc22758d93b1da61d8ceef46842d2a7abac60e9feb828de282499a6a1f0252c5abf0422649748ace217b85d2bc0fae9e76526fd2c4093501c5b71f7a9a3cadfeee01790a8beff306fcc52a7f99b10f9c28348da3a158ca4d2473e2ae74b3ea3ef76072c4194b96fa1183098e2c2c383943fc62942ddaaed82b40cb008fefd12495e7774a4af249829362f5f7e0364c5fe172f12ecb9d97422f46976e179fc0076642f72213b2f563b1eb99129cdb64fab6d669d87f282bfbab1f165514f4c81484db1d6ad2cfbe0e1bd63e1b00456526bfe7825a2d193565ab3b3cfe20c484096d53a3b653b254ee6010b9751044ea722c7655eab57234254233ecc2c08f95cb2720158893adac24c38a6feb9a18a3d3e210a84f0009708e520a1f2fc6ea332d2c458dc3d566976f1dee1c107daedf82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h26a34554bcd46d04122c88dfe2e12496e62c0f29585feaedca1f590b9edeee4ccc991b80357b58a9f8d1da23c90e67dfb47b992d0fd93f96d190e64810dae1691856ad18b85a1f2841bbb6bd2b73e902b346b39e35614fdc20214515b9330d58f63ce56a76f86f8981cb464c116e8deab2a191a6f279ee36d1915f84c39f521c50315bad885dffdd38521804cc36cd5faacf0613ef404841aaa61a78c4dfa7dfa0e33122d228deb018473a6ce45fdbe955bf21fbf6a8868a8b60c2c9da6930a61276ac5402166f0a2338f7a312bc90a85b778da53548c5b4da73ae1b7f4971998e452ca7b9a6f36079981c3124681596da15600d5e4d905e31ae20e5737ca7854b96c12af7c8be382213104718a60f79d5bcf72cdbabf65eeddf4f26038a31f9a396b3bd3f4592e6ed6ce7d8bfd7ad47ba2059ed43c42bb29c6b50c975cee260d3f87109;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h31d45d765f17e341117b66e764bd0565492ba44fed82483e28373a88588952aba2371047b95100401cf8258c65216a85f0efb3dcf94f0cc9e04dfd142a677fb9ed48c418bb09953b3ec12534064d9cf00c4670a9a02338346594fc534ce6c3da8fbd01b3eeff7c451a2d17f62576e45dc5939fa0c1fe9ead8f1472cb82640f6d48bfc3a6708cdfeefcc55db1dbbe97b317294348b061b7916a5757f1b375f570856a7a8b6e605eedd15dab92a930a1473c124c9bd1ab9c275523c0f6b4d9c7b03d3c9d7d54e94f7170c43ca625abc7da08b91c74b675d177961acaccd5e6b26a7fc2ead92229a1fb774bef1debf3c348a6744e21b2de3157592d9fc60505652f1ee812b50d812a1d186c44622e7d8bb822a4124bef5ded35ecc26de47780e5bbf4dc798f4883d81d59b41c302011653f53575ef7f6ea1c3db12d5fd81352060578993f9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3276e218ab8f6939c264ae78e908b67d90473e6ff46c65b7d0bd853e0a1263d07a935b7970b6f10aa29440f9738a914afcd5e5b288e5857798d00551e27814ac2ae7c3aee4ccb866b7152d89bf9a08c11d7e5cc2dfae8bc388fd2102e86879120fcd9dbe8d869704507b3f835fa64f183dbe2f95697967f9448eaf751317251d460c5410095e26b0b88dbb9b6d9fcc1bd555cac0c20f23845587d420baa9eb5a53bd4c1db9a171921ee3eed775be1de7071e2b3c45add78a820be4ac09aa83105682c3fcbd027a0e799f662f07132fb545712b5e06e51a5be215add36e8e04c3759f918490f6726de6bafff76bf8233c316520d40064ac16fd8553f491ce702b01e62d414b5c2712e858eb1a054a8182fa3407155a5a866bcf1d96ed91b54f6639f669ac925d5665978539b1f8ac739ba8d689b2c02bd842553080ddbf2b1eafc55cf392;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd434273207c72487ffce1d6f31dfcd8562f073aa0a270111660fe99df2c45482a83ac51d36a01c4ce856c9dd7a49b1ca80daffe81397742c3f6996e846c6b3fb2b7a7419fe8c6c94b8511753d33a0b5577cc75a56d0a9f93d4a698e22b6d81ca4bc38397e230480b9920cc0c31db45f26700f20e8c32851212dcfc1327b0a3ab3c6ed2ef91001c50147dd83f204d46e904efb6aacc0abfaa51e745ffc522f8f0baa52f8b27dda3312baeddeb8b248740bfb57984a1c6fe59336b148dd5ca7810edc583fded172851bc32d9306ce99d12e98a28f0464dfbca25141fc1ec3cef62539852a25f756e93d09ca4c0ac612bea401289ee9ce014158bc2135536713715768bb37f8d1fc46feae973c83949cc2cc95d9e7ee61d425f642647363ef84672e290560a5d924e599bfe7631f3d453f70ceefab7e858996435f28f1441980c28e7702048;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h36c31a3c2ad12f29e48584c382ba920e5425cdf938fac72dce4d2dc9dce52c1f611c48e8e3868d572476053242fe0fcd32ab28a00e71d0c728c0898d2c78089f57e513a37c08caa8fc150b5479d4b46317c6455d9ff0fb2a37f25dd92dc9a9fdbc6e8bc49eb8eb876627898c5c27eb5e807e56ba4afc8007cfd414faa53bec8bd773de821ff46dd02eb71567eeb2ab2ea78fde8e8a44792863eaf79522067ffcb5a87c2cb5f37516452b94b789a20f9044b95a6b97af7c411085deac79d4cd018b4cad8c5cd2a330113145b3f7974c370800795e0aa1c041c90271e1cd89d553ea8666ef4a4d5459eea7074c2281294351e6836166cfc35eafde4687e38cbd2af798fc28cc51a907acae5febe259f04ab6cbcfe061bd1ae42ae3b721be57ae661eb331ec8518570c055cfcd874858e82e62a54a772a1888ec8b02bd7a7d5f4c8702c13c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h75fe1515dedb8ed40f04f2e8c004a21413da95a77e18a15177bc5a296a0f4a7b155bac4d0fe5f1f5d3ebabff3118eb9fe72556cbd915e5b5db00bd495b680c3e3474b2177461354431ba6cec7e4c287d11eaa68e0441fe666ff832241d43cbe22e5a88aef5e701eac7c551cef8a9f2dc376a79877e319bdb3959e88fcda0fbf42b6fe0727ec9f082c17a9230424239678c7f1bf7ebbd931780b8cfaaca3933599e96c6de86527bf1adddbf35b70148c06f67458a75191b81ff5f213d9d71a460e24084171fd7ab53ace3b4952bed4629588b81286d7daef17aafd30cf68466ee25b9310b71a566c0b8cf51b0fa37ef21f82f71bc191228f080e372a2a18ae1e9206eef967511631aae13b81cbf08e4db676dbc71ae87671712a8bf88c0766726cb8a930ac0acb6565a8211b0409d0e5d4d859f227a6a528947afea2914e6774473d933e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4a7efb185c677b0efd7d02e65485703bf8249e01f2216b5304f85cf397af99250f277d8aab56196b74dc2be2f188591e2348111217972ca05b9f93762a7151ce33288b02a95a241a358df932ca7f8b51139e2ddc6cfbf76ae92923a2216633b3a64fa16a6859046d031c60af1f73d9c4852212df5a0206d70646357fae4fc201cdc10feb58512545f778b606c19ed2201f6e913c7bf48d7bac79ce0d8447f7a99b1be776f44efe502fc7d44a420c4474ecc4297a3f0cf842837863a9205615a68cd3290827174aad542d6c64a8bb488dac82542105cd2467417ec72b8a0c5a0948e529c6c58c66b1be9107282f9724dd602c7d016074af3f565515f9b4a47bfda2ceb81978095e8f82031991479c48279ac0e4277ad49e62a875e8a50daaf3a6418ea913ff737d46af3e19b0b4b7944a8858e2aef1ebdbe54f96410b557cec9a25ccd96a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hffb874bce364da54dd72c2e735965999bf881e28d5457e186f005e520d657af8214a7b000394221636f22fd04f06786263e6dc845b2ba4632dffe3945faf9de9c4b608db777ede2121608a4cfeba68849a2a8ce320fc9d7bbef48b2c6378933b5bb270cdb190d8af2a28ea5c7e005e2ad1c0e07d12cd4599ddf16aac1d19d2654b567ac99143dd1e13988039359206dd9387d21d0d7ee031bb9bcbe4a9d071a1d500bca54f80ba83fe81d8b65cf017e00f8c35228e473cff8d2bb0e85140853a26550a232f80e95c1a459cfd6a03825bf26d9b7975c37040887c44891b29b967add6ba6c084b671ce42386ff48274dc96b418c52f1ec695a206281f51bf6c76a05f4186c9625c8522ca504ce9c25350acb9a74e4ca37cc9a3b3a009cdfcb02fbb0f8bddf3cc8e48baa9a869ce5efa2a12cc1039f34ec74e21a75d533f1abca38fa83c2ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4cf81e2384504e1b8be6d17f7403ea67c4b2370a30beb52658976e0dc8e70e499722fde607f7c1af22845fe1764185df528effaf7b1e92b3e5fedda2cb20f6018f946e2320a10c1f061745b30d7dc1c5cc4796ea18a9394ccf4dd6660707bf1eee672d9cd5ee71518217eb4ace4c855f1389ef2c0b1ab86e6398b7748f508697bfde90e1db1a6d29dd346ecf72247937d304b61c6728d4bd67cc6ff025c42c7a4743e21659144fad87d523e4f15672ca2bf434a9f02753f363b8d84127dad991031038fed06bebbcc1fa0bee5327b62ce1dbc955a05cb662a48ac3c63697dba4f81673c53fcf80f77edc58dc68bc8a9f082e1f06ad717f2e6f4bda2d30c09d07b19b0d79e227b1fc5696668eefe3a6441786749118b7bda5f77bbeacfb04c76301f3bfe4b4f4a80b4c37c48beefd533e483d15e3304b7f871258edba35c66c156d9c63cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc23ddfdb7bdc18d20043b56e5432edc7a7d42965f2ff40b88bbef86ca838f95080250eb76b8931e1069f0c6b57a6eeea62a3c1237f8a50e1fc2b8f380fba9c950d481080bc7ced3dc0583fec1ebe7c1d85d2427c64857616f9ee23f73259b67c4299704a54f56fa8066ff92b2adc2633baadcfcbd653928c01543d615e0551907bc439a07b2f07b6931eb4b733ec0143945d7a907f4fedcc378a6a4d33d05b122b475205d3078319fa8e11fdd9195983fc9a48412a1d2577317be5d03b125ad0dfd1e2329dbf541ca98d6e525eba4798fca748232821af7c1b935b753281293012619377628b4cd392b146fab63c15019e519e7ce942d921950c7310a67e9f4598ec5db6d10c6152ea5166bfce5196b25a5fba9f8921f2e55894e0aaed7755fcf7dc581b726eb21cf003b2070db9b9f735d17afe596eef91a2e3c12513bcfecff2d317a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h61aba1ba99b366d7dd562467b6b018ca84a621b2aeb86fc9de24b5abe4a2a03e2619685999af918157d1df1b33a31a6b4d2b964dadd4dabe55283dcc450ff82bf647789084a227d9a3c3e57571e021fb4ed7085b5483726f82950aedf70206024aef04f838285da07e713af58546b27f7539b7f95526a9a9c89d799ae080344b8e8e50de599c7cae9981f126d16b7c3331a9420121c8d2a0a9ec976e4c579cda6c1156478987d80861c3bb1f6c83d6376ddcc65e7fb587c02a239a346a4770869cb27c4a292fb1a43628e47fa8e859e36bb8d7df2c1cf1121e50af2b3292cc87bf1c5d6b6dcc5d328ad2d4bec55643045546ae03e52a275d259e41d28d1592efa8e5d401c2f9dcdca7724dbeae0cfd7853e55c9849f05ceb1b1f3b227ecb965893fa083ab605b528fbb15964ea85cba995e671d8febb27b31279df804512d17085ebd5fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5dd18b346e16e69e26031b31e7f4eed3d6b623dcbd4cf901c920be82cd5360a96200167c9341be3d116bfe42d07c854a9c8fa7e0a04cd25455ee1dfdf2d232e687fca4392ed1582188a682071316b38d93fcc02b934f170d32fcbc856a78e105e4422b2ed7520a74db784c5a3d9a21a9419b07b42591d3453abf929e16643d1db8e410011194fca64d845070699db0c0a1f4daf38f12d218ab20b153fcd9db542f864fa47084e102a7a2e1b2f19c2a61285dddd96e9dd7aee8de4795c994d86003da6b246e55fc15ecc9981c679392959eaaaf5d100077e078ff24f43128ccadc3f250d4534566eab82a0d88417e382ed0c79ffc5afc99eadc3b98b3f67cb579df6ba88e672b4220c7791629561aa21460062d85a0291d6e0a4ec94de69415232dd459e5319a6b6ad9156f903ac754b2e2c4424741dc1b1c1737a7a48fe86f1f3b98603c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he00e701d75b826215e544266cab9090c2f78dfe66470b28e859c73359802dbda49fe11b5d081ada2b2d7bac935f718f09d4810025a520e4a1753d6ea05cebab8fe2f5eb9ad742715dde7a1a7639f4671f364ba1e007d783da9f14e989922f329dea2ce62e26313ad929052899705472354365d485322dcba890bf4e37669885d9613a1c81f1eab40173d1e850875d452e7d442d4f3010fd20862e648eff2dfdea7b907ecf12244c08105b7e4e4482275ed656660b330f634d3cd58c699b817c34a4354b3a40c0b32b63aeab11766e700e2704396d97eca5516b3aa2fbd48c5f1deb7da22e994851f41cddd1c00e0c533e0145426e6be199f96eb68dd8fbd66ed8ac24c0e79560acf2f40e45c101a4c3e5d792d16d69f00abdc7acfd497f0443471506c0bdea3b30d06b4e506637880d9051ba7b79353082292d98e9bd09bef72e84080b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6c7334ebb5351b7755d9bb15d40e4b6180a380a80e2df7c0b60e6436fd379e5e323f36ebbf9251e024c2e1a832f1154876e9aec963351f1deaf4e129f24e1a0100d1cf82c1b0f7fb5a6316b7ccc19311cbe36fde6a6dbc0d62c9d81ae575d58450a78aef06ed1b2c3dbb895140200a8c5e65f5ffcb49ddf8fe184cd7553f3d2e09d92ce29fba69861e6b364280e6c91402081aad88d2b21ea298d6f7c8768f5adcfec3d7a1a16dcbad6d897d625fac860bc8fd7e2261d730b8ffd3886b6dacaf23bf6672a13f7ced716113e84e68e42d919ad90042b2f6ffe555bd90b15730ad3add985e2ee6d3923418617c040e4f7527b74a1cc63b004a23d03d5051cd9282cee902a06ea4d16a7c66ed3d75b09ab3aa575fc5d10a75dbb4258df799f2491f9d7353f53ebe6cab59ac1f042c7c692f2007bd5eacc12117b9ee0a19e15f850f1ab7643;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb67af1d9f1756693ab7ccaee8762db347090932b3504ee3beb55fabe2ea35c0b8acf3d16f9d7ddb101b443946d1af303952bc15b758345a48f5f889784777c6e31366173efbd7acd881801c98590ab0c279b615e19225e75b71392fb98894dfb5f85cbebed122ec314e4589eb4e16a60886b260d7c09e1ab61a84f0a0a40b2d6cbfdb33bb7bd6cc2ca68ffa4f7c5c59a354aef61bff50f9429878766bfcf11d343b93d8c356afbf078a8ced5eab8e7004b8beea45318bc4e0c6ae75d6e11c3ad38c835868083fafb9ea52046f186716fff6577906ea884106d4121b3eb0b1bbd4215be4912b4ed745e63653e51f3a11fbbb94ce7e54f499f1985c5fc78c709f996f7b9717dc04f76e78886ed3047b8362250cf64e6fc85c4ca992c2c0f1a8a5cc5053f899d43a5ba125f6f6368a98c20cc0f2fe860bd45b2269da959e4cdcd6cf0b380c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4098d87915b3c56cbd62466fe34d84f4e36e8b1c684d5e8780fbb3a6a5ac181a6ac96375a2d28755518edb94a03fb52496c2fe6bdd55baa03b2f4984cadbb076fb007a943a5e1722c9ba3fd2a4a3fedd4ae3b8ccd2681813f3160f538ea225540aa1776450db844e0e54e8c25277c5103577d193d4c53c53c39e22aaa3dee1ac8237baf5e99977c84bb08e0ae7091a00dd4105ca027f65df2753af41ef09c0efc56766b301387f32fad5da37a4902f7f24d42c6deb772e203fad6dd0a81a472706223914f62393c13a9cdbfc011b4dbf983efe47e31ccc59f457b9f2769887893b228caf452679a5a428b29e5cc8fef4b0f3e3f367dbd20cd62c8dff7f6310854fa0bd494f1e7f00d49bb867e1b831e63f6628df5921582b35007e671d490e741122d916f7c11ed03eafe1c0bee0e01e1a1941209f4fc482a07286167205647382bb8e39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1a4716935ffbb6c18a0b9b67688a830a1b2d11c3214245b0bb596889a3996c11391f85beb85ee0377efb0ef87b68c94cc7c88e59a62f2416424e8056fd2d1e58be423a64a0f5dc0b7d2f01d75ba86d2c88d47fddf0eea826f060a6c2ecdbf715b075c204a107ca57e4a1e3bd06ff3d40023ba22029078cc7b11b70c3dd135633b55664feb511231e77dbf1cd59565cd87e47a20425783114f3ef7073a32ca1d14dc7cd37cf49210730c98fbe7df68177e55fc9bf2ac7fb9ed80574e8771fa7785397856aa331f290908a767c905020c90a4aff2d700813d2620ba44b23f323d1f96c13e534d3e6ee8acaed6c48e9d0651fd0eda552b84a3cf837b3895e19d3e460b76fd60571996f12be0e36b610b355ee4c794ce943f0a875a46eddab2dcb0aa5aa557c89ce0a1c2895014f75ba676657c6739855520ca9a37017c38a920295c5779d4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h314190cd7a3afd715569c065fa9e3f14730781f0c6fb9b1d89ec15aba5f6b707baa7b2524d506a02fb7fe0ce734f761e91360c483014047456b55e46f46009b86b7ab759bdf59a9869d710143a420ddfa90a985c7cc81817434730bc40c70589100414b0c0976cc003dc5505653e11078cb6ed2de7a745ebd81eb7b160f8a9928a8293088fb661b1b16ae91084ebefb981eabb5b4836a0bcedd3d9682e03c49a08bbc3ef6d08d19e3918c2c7c043bd6775e09ba10bbd3d3f316bdd43fd61badabe6afd8d2cb96098fe5103a84ccd74ad2ce9ad2918a9a3c72e6b5332998bf02c578c2e84fe3fecbeee1f44793c1b7b240f8b49d61cce87ee60a2e7827d5e9d44ff2b9bb7ad9b2c95438ac90da13525d536a061387974fdd6de25c7f92ba08cef8d0a3c9e899ee7a8afd95095d339f255148decf56abdee18dff6d1fdc3a0aadf7f2fb145;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hbd940316f6d09159e6c111e6cdd444e9d355d481a2482805eeb58cc489bb3394861e163212b032846cd6311f82dd350c4969744a8bef4ea825d4f2894469e193f2c5324dd44b5a8b139049883a264bf256750e1bfd02cfdb599deaa45a8ba88a119d8be18df9ca737bf497067ac0a84f141bd455be46c9794d52e39c912e5e0a5acfbee78aedbbd4043e9982baadefe7174aeb39d3e2db75cbee4feef621e11975e310061a290f62cf09e108c8aabeea8fd09e669bd31d027cad570ca3e404bd366a17512b312be27a14ee1dc88df1cc02ba46a4d74bee5e0c53ccb9e2cc8bfd89157e08fc20484b978d7c570f679d387389b0701a73c83ee772fad7b935e94d10e1f8cef8d94f115815c2cced739341e0319f9fb02fa1971d80923ec77735d1a397e383008a42eeb6b8a1d0c89a15a538a16c47884723e23cac20a944e15def9f32b874;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc124759b01eb9861b3fd8a22030b9cd7b08f12f6a286e15001abee270cc5ffb6bd0a7391f6bd2a0efe03e07d3c1fd0df72c6a9d119df65727a7da0c714afb1b4a3ec1b949348c12aea1fa1acaa971cc5ef47d9605b57b3344a60fa0c47eae81610c7ad8fbb1805f1481df26847b78b201175f44aba214f66240c9008cde82356b4549d54dd09534163a2559c1483b3a43ad30fd3d1309985fc59a0d0954645109829b87a7a67f526f3c15c920d24ee27e3c2c429a29668d119bed63650f0c7c4ca2ab929f5d89dea52ab63f91778b29ac231b41d7db774bc133afad2789e28c0efd6c406ba7c6e72d11590cc2319119ffd3471200251967af30e0f39a3423b280725be8cdea5a666dccc0f460fdc9a14ad6a2be1f5f5efba0594d8b1b250624a3396aced8002de01d1c8031bccef9c1707334b2ce5e9e131db7fa5fc42a6b4eba14d2757;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he459857aef86c9aa71c393638bc64e536ef51dd2a195f999d3d4504e3fbae0ce47e05fb57b7403188664c5af104815b323997ea2326e7a9015aa516e66facabdada0bda0919e0587dd156d261c1c5370e319723c0301cf38d2ae95e3b226649d5d259dbb5ee673a201755df687353e950ed3937a28dc6fcc2ecd0e9d3d61aa097a474e93460a06d19a0b6f130e05d1c8c4a5630fa837c669f4b5de0514ea00b9f0bc8c03ad9d6b27ec660199d90ac385345358b2f6b525bff40e83a27fb991731fa8d955b5b6a41281501e610f0351418857192139e71a0bcf79367ddf55f6ec59ffcbb618408631aaf09edd1649f24a7e206639ef944947f1b0b8475d4470d4aea3c695076eec3a5820dc082c1d232c40402061ce959fae4633f89260f523b091fda3b638b2bad044fe08ac4295494c178bad0a08e0e6cc13aad3e1e0b2ad376a3b74c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha6efa95a33162adc93cae6e677127ea96d41b9fd4b3d2c44f3aaf4366fcc5f5705cd378870feb33c1b0a6214a05c87a3f1292997822d1c10b759ee8591ef79297b5179252fccd358774721525dc1d5e8b2392b64aba3092fb8ec7f3dfa76ee2eddf1f2548b16037d1a612105eaf07975d8b6a464b6d0a5cc83737ffd94c39792362073b4a5cae581491aa24615c822950382874f14ad2e78fb7a1465af4c70e190ecdbe7ff78c537ea317d7ef198cd4eedfc3b43860ca88cc2bf12ed5797e8e1b4fdadfa26ecfe509163dcfd9331429322c9062bbf49746aa93f0783760dd7ddaf6c0345d68de285f0288ee7c7ff2aabe3c02d7ccaadefe03e091ad0e1b718c65bcd06057b5c2b8042bb3bdf87bdfce5de9204321471199ea1c9e0fc62539c6d0294b34cd2f0304ba0df09e5cae8ea0eefffc37fa65aa3fd579be1fba861eb1e7ac4a957;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h24d35df96fb02efe86483241bb09fea9321a750debb849e90ad16e848137d8a263a537b921742907c92577d3d26e240c398b71460e514a1fb23c92ff25f2d92d2b481fb3273e4ec406270d958ff0b1f98c2b367948a05590b71a52d98d4771452d82ffef3fb163c8b566e54ae3e4c1250caf8d7abcb47e14b1f86006c3d8d056971ee126b556c76f1915efcb9575e261b3f905b4967b39b7bafa503363c864cd5d898aad8323130304610adb5d14ad53a6cbe0883cae17104708d5dd1b9607faee761e6fcf6a9ebc2b14482cb808751e4aa94fc18fa342982a0416797821659affaf568e6d2480c8296a9a4f276da203ae871ad0553f03b4da4fea7266c7842aec347f93f66f6d679408694bbef1b4d9ec2722000ce11a0e3a2c8df3eb05d5b2ee33a86d5a4c43a4ce9c977d5afa09abfd18a6f987311cf43ddc127e8bee3f0221c8dd35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he9efd7dced76aed1bd41ac275e9510984f522c7ed876c7bdbfa653b140f50410de0ace5648bdb7eabc35f272c0d604b84bc1b1a214188b3df5261715bf4fc93e733b8550e1b2ac9a5ff85bc0e8eba393505b50b57f8c55397a60a1803c336d338bfa038448d7c53ae5a4d5d0c4052da0e5ee7aab2782feb04f4bd0d1bf85d37539e6a0dd755e99d254db87d4fa060267515c5f14815780bb1cd8125efc27ba35427340f4629659f8707546cd01bae0185408a9c4d99e4c8457a4459eda0906e4f77e77ae0a4b785d672f5739fee8a30aa208a5f5d82fbe4c986f172dfc4d445c810b7ec1d3a9f2dd094dcbf384bb6c3ab785c079a49f72e66895f782169a860da58cc28a1ac4d83e744a4a56e6b90f706ec9c524ed7338906ce747f4f49fa65f225f0b5583b581921f8e0d00e8269ac3e558582fdb30b8a416f2801030eafb95b8b388ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha08d60ba116a81789ee0909db1183f568cc55f5a37e366c4a2ff975c04cea4d5459a6c67ffa3be97c120ccf4d64a960f5265c2fbfe9ad328d3de3204f89835a373d20439f5e7a05e79e7f6d2ba293fbbbdf146390f55ad2c7b77acd9163597f894e6418870afe44a8a4e4257e7640f03576d8cc507384443812cac7c9efba79fc9879366dc78c916311fe5e269c46fd527e18cafee7231de76c1be30c7acfeca1f890b64cc066b63181c0958c1fd0643039597889cc182c30c45d867876530d99dc3cc951b1cbd2992560bf9de796de347968a05a8d40729ac81c35a2eccf803356ba0ebaaa278490a96af8001c36c68ae94a4de0235632070acd8cc6f61f09e31745b907060fb60e489bc2af5fbcb6c940e3194ba3cf1b623ae7d228fe79465447d9b3f4d7433c40f89adcb2e347838548bd39691f6ce1242cc8484961825bd1c5e025b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hdeac6b4a8ae7d2b1665921a9c365b532ea967c766c95161156797bd294886e458283dce7320710df90437e1c8e8756859ec8213ac06bfb198b58346229e197eed1ee9130aea9564a9a80bb1a86d80b25a7ed6756bac81208af7afc4a33ae6ce20e4047c01cb4009d2afc5cde25bc7a16efcd22fd0dc6c94b68b9c3b71e433c4e6144da43f57f9b47a91e7be0481c5a0165642b27d9262331ba139d1e87659c6d3bf8235b5ab0c8084c33a338d9ac9ec186e4cc7d92585570c827846593bb8feb25e9e96aacde5df6bc79d10aeb755adf0159bcd1e0efa67739795ff973f49c10d917ee7df3e46b265f5f180120e393ef8cca6053702f54e20d444d44859f1e5e2c12b7a39ca04cc587366e6fdb2fb037fdb92e84609d455d53e656ea71360f0ea46c40082593e0a21550123587fdb1ab1d0e9fd44f67f69ae850f029f44e48729268404d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9c46b699bdcd0d369f4b44275dc84ebc853c24d5e49132b717a7f088463e7a45e47802b76c9b27f23598e7085c0a44aec09ee767fe98a7b83a506caa2d31ff7ba70be1cac3b2e5d3e66d2ec350a1abbf2c8a4fc5e97cda1588aa137693ec27ae447a62262d73beec1f1146406d49949e93170b3225e10e529442795199794eb56606f812e70f3a95374ec0837f26e04c4e7ea5dcd8496eb533fcb728fbf50f382f48ba41e2faea8c3afa33fe1000c565a3153a1a281ec65e4d76699c358c243577ef4e9b77b98c5e70328346b6dcd379ea60cc695f04fdff81ca59f6548e9e8323323b3bebf4e9dd4fb0e9e59c5a2aadb273123740c691ba605beb9eeace0ba9263bc84b829128968e5b56144adb3ee1b5d920d67ed1b0a28c979d66718307b31b885a048ed2e85805b1c6261912bc12b783647c5350a67d089361ef8b3f425b2a846c86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h79fd74df92f0648ea63c9da6d26fd2c701d8838bdf739a56f1bc2e9e5344e7ceebf0b38ea9396dfa30dd970603f24b1fdabbee4c38f693c48ca4fb8a4e5b2e707a8981f6cf52fa49761e3b27940fbb14d0c776bf03db3c6c9f23a3117f860fa9ee4fa337d5c2d9af2189dec71f39cd46bca857d8f6f70273a531837f44f6de68044b63ceafab6cb8824d213a45452b333370a46ac1a7abe764f8965f73e05a841c7637d5fb8c1be9c835b3f7afb7661c2d85e1f9dfbadc04d8a1a3b6a3b60a92a99a82daf3ca973d00f64234a3f02a5daf2e9b87f4ff874c22366b06634e4552ebb5598ecfa85534ba6dbfac6de54436fe0aaba70e27aaa0a2f3677c6b0c9f2c379b8a0e94769fb9deace523f0c512ca9b171ace48a002e45d70d1850565c1dbc34876a6c8a89f5e6a9ee95465c800936d0f8bf5c317f80c822c5fb1ab5441ffdbc9c4ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9525e655b7a6bf10d5e3210e0b39f521ca3d4374877f07a90f73b75cb65d5b024f8662af2e9ce278da218ed1cdb9dea1def13012489a61d991e88453848be192f9ae623234810ad8ae3796239111097629237d4e0edb39733d8343e62307aa1f24223b8c777abd7d63d1e425e12cb29d9bb7206f2c17c8ff0d4a25eb0839d41e3e2ff3ca4d1f1f1636ada795b4d46d5dbfc1ff732d05b555e7ab0b7724fcf7c012abd41e65e13ec50f8d91d23c1b6f3a3936633f42d872e99e1b4c4f70b0a5aafbb465affff6114c86b1df4bdc0d80d7b6ce46a7e318d6a640c575216b34f6c125e0289ceee4fbe985a17af6098a26715c9019b1341bc32ec2c1604035ff259cd1f2a075cf613329e6d1697fd22ef2aca7a1c38fdb846d8e91eca9a8efa6f31e58303aa469da299c22ff4a3a0c68e5ccf38662037a234c9c03d32d92ba0d82ae154734dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd93278b579c2aa332c8873624042ed77ddc5711abc920f0c44bb097383666e99dbc74f8b1ed957a2cd08621e1d7ccf38d7773276cbf07a424ec0a04a1322ada8f59edd8887d429463e5882ce67416cf289f092a84ff418f2bf198d6f7f0f6d5f004bd5ae1806dc08091844f5ba58eb18701cd1ce583da6e81ac9aa0fa8acc563e07dc68e879ed2c172abe128c69b89306cc54c58b03e3bfc361a3a810c0feda1b4d7d9e49686dcb9d59310d6ebe7462b1ce0ec3c44cd39de507cf42a62eb796a725f9acba089f243d8293eb7563d48b67554f97eb969dcc554d3d5a38c2d3dbc9f3cfa0488034b297d50aaa26eaab791d55e4536438cd193d10c265d904dcaffc3dbd68341599cbc65dc2fdc3746cd578933061a6ee0cdcf83cbf29aff7180fbfaf07367666dbd164859d67229c7713778fe7c6e37ba248f9e1aad57de4d6c5a1ec83a19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6d050bc4d2d028cb032ce9e96c3bf2269e92390499613654a78c73eb8661c6a5c469255b47377b345bd32a52e6b4a43966fd0b84c2cc85e15ce3cd85af4723da8cb9c118bbb15c168156e80a6a1efca7c4298487bfd43e4a26e5527e0adaf64df47d9e0ab9cbe90254196bf0ed51d6d8a8c7418f90b10162d0169b3ab92fdb07c926183c3e0fdaef02411f780ae76c320a0148f0d780dbf26277cd31de96c792a9653bef62cc0af54fb4d9050eb562770b4563b5bd0cf56ad0a2e9398723edba1def554afe00041f78aeba21d90e36974a882f6273c1a665b670a6c8e744e41993b5bbca0ef3da708e09190dc425e0df162f0ddb53540febd8be35957fd7195c59159c4a29be05acd6b6f32f71372fd4b23551ee2f344241f6fe9fca21bed2bbb4eccc8b987ae4cd2f72062844b142a76888992596cd19925939692df4c5839f3e36dc6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hefb69b7574462f16a3c96d58b3574d018b9fc61f1f8b24162e3e01903badabeb2dce27a299b8b7e38b6d30e19091e945ca77e8af7971ff40be626d4785bd823fba0c66eba5371ef9cbcad2ed987b537eb9cd083b68398daf7ff2eefb5f624640bfe7c66ebb1b85be349fde8526a9b11e00e6d47068b9aa572bd18290e7e3f1c9b5821a96d13364cfa676adb020728c6576b15a6384ef9bca8f93481520d71ec7fcfb6842a9bb4724915c182d4ef16a0662dc312c054c64a48718b440b58dc6f0930dea2604ce8feb9cda0e8edf63eb144994f0caf46e6e8f691645474df54ade4df6c18381b1f40a09f6564eaaa1cd094ec37a1dd73edd7a28f21f73b035bacc558400aad93566b8fa675d0c0529e605a84300bbc241e9db50221f8def16b7eaaa53be98e404a604607e40faf3803431b98f3b9f30be6b7215e7e83131ecbe2ca1ea5dc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1a77f71a658106980ed3e627856830755312a7e0ac569eda25a609cb280f55e9a138d610357f576f69b174ec334cfe33e71743fe301b40f54822c4b30f4c15c6176ff12d4dc780cd6d4c4481d8a97f5bf828de0c9940207fd66755c5b04c77351da534236bb5b0393332f9993063302bd85e9859ff493bb3845ab6ff1f3947102672fa3182a0b20c9cfcd6e42f084ee96cac5ab6d42034a017e280d4a1d388c1ba132374ea73796282fccfd722badf2ac7c08bb17686b7a69eacd89b1450df726ef00cc8fceadfe62c11dfc6d50ef12fb6ff12183ac3919f3b6b0fd5de14abd9e2c3ce866d54fee266a88a32bbb8dd4aef52ecd6148ecf32acaa71de10ab9c97cf4f2e59c72268b76c2a205142765f718ce09d1692de2c2fce069f127b51c9ad79b34f8e3efbac8ef0cab3ff356cfb484f01e5fdd7cdde308b3afe6df5bd4f393ccdedbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1fcd4a3e8beb6327d93aaded98e847b43b0868e80ec38d5c3e3850c45255536a85d22ad9254e7fcac750e8391ded88c6af96e14ee5c2c3c27477ede1ec7a29c7e7d4601f3ad42ae15c862c0622ad8d8e60fbc58eb43bdae93ddce3c962276d8d8c7e29367ca3165fb8cb7c5c806b2c00a2e800a1d748784e3e4549da491eab0d018efd30e3a5bb7100ac44c902595dd1c93adf95c7d5a2376796f0466385d4312772853c7b68d20760e392844fc2f2fcdf652e393118a5ea6a32b7e6f0827663db2c086885623fd9a6ee340900d9669cdb0ae761bc78f7f61cd7e43c7311a02049b627fe68f4d2d41cb72661437960c20afc3af9cccce32e5994193664f4cffcb03bff8dd1dabed968fce9936e3acc58ec7be841fad47a6fd237d3880e295771cbc4f1763166e0370dd00ed98f42121caa3897b0a5fdeea1541783b47f034bfaf2a04a58;
        #1
        $finish();
    end
endmodule
