module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9735eaff175a878a3c7864804;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h185f58e35601394df45ae0357;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11758926d282dda56934a2839;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15d0990c5905364fd22d1557e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd2457d05396bec13eef985cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7094a9f64dca7047644e58b27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c0bd95d0b1f951e4c23e0839;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33694898084d54f402fd21757;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa8d0baa5a964b044fddf3960;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h624075423856e3356224f5829;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c3b0db236f1598a218000732;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h970bb0f157b59010e23682c15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h193b6717337a3e23a1fb9723f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b8e3bbd064c5c09cbd12b9cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5793477862cdd1dc7209836d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5be388d3fa9aac685437a8ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e89faa3447d64e8bd1cca836;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha45be9b3cb60ad0ad395112c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68467c8f49a06d53b7d22b266;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f5d431e3e71c88a63e00ec48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc7beb1f1ae0e77b4ca58247f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d9e0c18e46211282d354034f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h367eeb85d5d48e03b91852384;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h474cca4db334f6fe53484e606;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4706160f49a01f25fb835098;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a24088a6ff080c610442e7c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h575b0196a98b8c76b33d20252;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6da01afc21bfbed1afa3bd08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc41607a0f77c7e4503b21938e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef10bf6c38b3133a8121d9c29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92b4faac0fbee8432fe6fbfb1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb54f0f8a08933547c9d8bca01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef9650bc19d74622d29eb6d07;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h659630a76d75b098f21e761c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18b57a0090592de2a58a4fb66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a1f6355bd74ecf0e7d51453d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f5d28c6daf2d075c2faf1099;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3849a28f09399fca33cf6bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h425d0b8db84690fbabacb18fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbc7236dceac371e667109c85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf94d17dea948eb221e2a3cad3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habf8edfbeb2aa530f20c420fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd63ecd2c4f68d55cd4a091572;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had92d6d8447f13e4d842364d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fb4c1ae536e58e38e9b7888c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb18da4959e9c1a38b7870290d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4f369681370434ea0b0921b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92711a61654dc7b51eaf31557;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59c61db7918533e225d98fb86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3233cfcfcfa57954f3c19a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72114201fef1c6474cee7c100;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h323f9768e0fde8262c20dd485;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h558abd93ac7e333422a850360;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e4bfab0b927328f3c0174d7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46dfd23d245d31c007042134;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77bcb25cfc4974c0c467a09af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eb0da636e8565b463b57d10c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4996a8f41cf48c7e6732b618;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c871d11448650f6a6d5cabc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15c72859b69b01362e2f998e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb00c5df1d17c739b85ca3f042;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h751e79b7756e422c79dc5f0d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22e886d7e05df31bc5509f185;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1591ff786213d9c8ee6151a0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58d5015b1b4460cb50730d571;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fb487a16f5f11654adcb48d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38c8a177f7ac601775a0941a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b2af2e6853ac2be222ea2dbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h642d493e4e2e1fca34faf5b01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef744b7332109ffcdb5deb706;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a4a32875825add4cca0aa1be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34c23935e2759e8b05b519e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3458b9b1d723f7d4a916ff15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96dfc2a7799f16edf9b2dc150;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbd7079cff16bc6549bb07178;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca763f80d25c38ee8c789be1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbae80c3e53c3575bd378ed6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f87867e8ce8012a127a110c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf7bbec8d5cdc580318ac9cb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h117aadb15edff05c12de456f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7094cad86861d53388bdc89e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd333b260c701a5898ad40a1f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd99f825af38f1af40845d053e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h845f0c41e91f3a3313ceedc0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ec254d477b5640a1e2159e5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bdf23a6b421937f7ffb89ea1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dbc30fac3833e27ec58fd183;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45cc8be9a6671625b1441fd6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12b3421d442600645ed069adc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42682c7f5c8e7adec89f098ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbabf19ae592b7c9111b7923ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd64f01070a77a15ac251b0cfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h797f52ef7bbc99bad0e53667f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb145b917d8f28c3e2f65cc36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3385fc279c1948536625c9e13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8234f8eebf8d903a02656c3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf12330e7933c437b5c6741fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16599fe27b97fcc2d0ab3fe14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc175c680b51daacfbdadd7e20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d9bb60f51cae09bfad25317e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3a0a9820dce358d7878393b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dd5385a1e3bdece1692bf525;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1074fde3256c6e20e3a544487;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16d4c799a93d71c0741f34ab6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a01d51a5c84675fec4a08a05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha05c73249fcb9e9c6e55d0b2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab3eaa15e18100bc135658106;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h693bd2e4d85c73494b2051a30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb4e3f9a83050e91a49de62b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1223d2e7f71514439da9e402a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc4530a2709c61e1debc3ee55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58c3777daae8478625c65f032;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd34c6fd764beb255517ac39bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf414d572584cc29245bc3a8b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4333e7269388349b7106ef9b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83ac7e0cc5536c4a6654ae6a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7e9654719eba6cb8b52814ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75adca3007ee2b49317b38669;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h516fc21f8c9a3eec04e1d99a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdeee93f0737219414a31f6b6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce99e146f612b1351ecdc19ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51caf7df40add4a6c8710f021;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h771f7cc1d5a1487a8bacc369d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a7bd118182e52c135fc646ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf98d689a55ca453b2128f84a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6abd6b9e2adb421bca546aee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd0a6d51d05b5b0e617494600;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hded5880f3722535616be689d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc15b57f4fac1112683ba10209;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb987195ed8df8308db197358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fabb1c479f1c794464804909;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6cc62e0a3becb558306b9525;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbea55d3c85a516b7536b33f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h888a32e1df2a24e7440e3774c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h658746ee5327f839d210f625b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0c608579b778832e0783f909;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeb914cf8fd9c2a411967633a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6d1042742a97a40280ad9c4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0430a75d7ba9461532368125;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4fa6cd43506cc56d0583215d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf64fabcbca5a6599f7578be0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e8c6dc85144f41b5986a334f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4115cbb5166f1e9ea880cc060;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e11bbfe66a019dcb64a3ccf5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56e7e7e0362afc62cb9ed0e54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61960b900042fd7a1b67fb123;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35e3fc9bff82578e25456b9c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf3551c1fc0dfaab40b6e588f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa5c2f89d966095e966262ea6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b47906d33f66aaa365b8bb45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h993370ffba653cb766db92b73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a75f8798829320f87013d715;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9f1381411eaa91e39f9bddad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h760dd525c27bc9e5c5b8d6c92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd216f902f67c1c6e282bb7be5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39ee10087293aba9d591e212c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37a1efc115ae409ebef185f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed518bbcfcab264bb79855c85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha288a97486f38c20dc052bb3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff1d9914055e13019c82cb9c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d75d92839692ee6514191741;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2dcdf55a430fb1917f08c9af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcccb2d476786ff0385be40f0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1558d531073e56030425dc75c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83b8720f90b74cc9f69b3aa09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habacaa6b8d3a1871e2c6ffdcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc00282562fc74a03e8a3cb84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9694b9825f971bd589c811688;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebffafa86d6d6bfeec233bf1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ea289a37e2a2f42e927ef803;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6d6a6ebc83a9dc25d5b2bfb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6894290a55f0ac755e19154d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61521e4d1f798c6d5669c1170;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9205f9841197e2fa0644992be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1b9efd268c09006de7ecbe09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he54539581dc7cb8581e3fbf46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75e9df53c8c02083399c4c18f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8a5517832a0a96040d7a02ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38a2a22ad7d56457733117928;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2c686a87dc95f464be38e0a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9932b454a977bb06ec047123;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h160e45c4663898f1944649960;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72f8720ace6d78cf7c0760c3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe666eecda7964b0aec7d66e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a9112cd907458b3f78efa813;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84fb252c223e793016f659c64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1a30fd5eceaf7ae23c42842f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6da6d464c44be9abd45dd9c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb0b9e36d34a29df5bd9aa31e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bffaad898ccca9840fefa8f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h626debf64704fabd9f38c9aef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ff30b9529c1120bb2a6360f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62f01a6389a8c3240033d80ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f99662295d56a0e53872557d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd656b73da413bfc04b0600a46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b0c0b6e774a8810e45af1b73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc53cf6236a8996a1c6d3a7907;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbf4beb335e6c58d7aed5a36e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc914febd0e8185a2c9ab0695;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb934fc70bd13313972d7b2924;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h831cc6fbb0902c8f5dd2f6f91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h735c8e2ecd1d2a77a8aae458e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae05139fb86570e66c941733f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h476a5d720569f63da8c42aa3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae2d82009434dfbbc5ceef430;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b8a0759b3d2344943564b043;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he76fca25bfccb7d116a7d9b44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9f4e724c48887165fcda63cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaa7ce87ed5c8c2e50bb48ba6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heaf90dccf4b1dc10e066580d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a409cb911dd81f060fd48a81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68c0cb73622001788fef5ed85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6348d1d354364b0e25c3a08f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893be3a1e37978814c7b9b28d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46f918282a3820c0a36fa7b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he351e3a54230e009836450f8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h898c82038a5a659a9f0f1a3c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h978bbb011180ab455d9872;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1971451e5ef8906a50204e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31cd3af0144fb26987dd39e19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7076940d3186d02e9bf7bfce2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3146fee7fdc3c7aa070739c78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ed851a5691c95ad4a036cec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4827b4adc1c117543bbdfa433;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fa58b6af3015ab989e60793c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6f707b4330bf9dbc6ae7aea8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30de365f7d4225da3ef2c0a55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9de65b9216f145285ef3ec33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6003d1b666f495d65c92e5d09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb77f1c2388f1a5619de691e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab39e12992fda7c74cd20dfbd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he68de3ee76ff9a0b14621f605;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c08ad4ec4d4c6fdb920cdbc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12dcce6e3a8e7da67d1fae714;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3297f38081080ed097275912f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha35082b293b1b1dc95fb15b29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3644873c84dcfa4cd452e454f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf41c32614c6a65ab5e1972af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2627b6c0a3298c6324409ca8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2407408e5f6431fbd9a44141f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9a57c46177609a487ecd05d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4faaca962541440c7f154ef55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81d619c745c76ea1f109059bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f1a16598b289fd2b1b893c6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb35bb7c63f224d43fdc61e6f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71203d6aa1d00ccee9a77fbb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9e9fffbab155abe7ed7c1219;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4d52d96bf6320e60538fc209;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3f0d93201f774e296a86b019;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1034578b6b772c8f01bed2510;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cd3a85843c80dfd418dcf1fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f953d9a8532ed54206b669e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca61f302e2bc7e23ed3e9d14c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b94b29ff4c09164a044cce85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe888b37b7c67598b76639950;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h665ec87a418b10ebd163eec84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ee5815a104fc664e3edba8d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74f6c89ce9d0664cb908edd11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbca0482f1ffd7d6579d6f6b5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf00a849e9078f9e946d4275da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb201cbe325f804a814a381130;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30d886b7b59e6fa36e4ded5bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef0255d1cbb712220ca201c59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17c946a3bc93d5aabfc286192;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e6952455263c8ee95c2bee50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h895bc2204db92d1f1ed271bb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11620fe9723ed04260b2989bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32940dd978a65e543bf57bfa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6934f28356140c47e0f3c79b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a82e2df64fd6a531a6622718;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49eb70ed2d3466fe94d2fd2dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78a6ab1df882b329304e2e0b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23a79e5d0d423a57a088497dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4155089be06dcb0067791344;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcad4cf1c81df757e4ae5c2efa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5d3cd6f9d5e96483e5aaea3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd23a1012d28dd2cfb5f898e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22a98af5c1f087e7bc957cfa6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8d0a32258f1aad1c7663d93f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2149c627308ba221dd4b7fee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83f81ebe04adea05a133eeb86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2de5efc924de6ff52cd74f67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h104c41fbe10c759e04f21d501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e82f3c2bd1a338dd231a8979;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a5bff484c4965ef6fb7de4fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5e44bac637ca96d082ae2d6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e58a2d79257e4ce2e04a6c5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h833b9078f24cb8f4aded539e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8034b28e60761233852ed2e9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a0e04e1337e8233dfdaa518f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0100d94377e68d771e9ae4e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2abf4c3b2d2c3940695a7007;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1417fb94fbe4654cbe8486b5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55df9cd5d902c95828c1a4f22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha06ba5b34018bc11512045a30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12d312884e33d4c379a2ad57d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c0db5f32af8c62efae78bd8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfe010c608ab7b56daf89d363;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3aec6de660e4482fcd88696d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1733ba9cf72127fa44bde717;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h526412db6abaa12260fa3630;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83c27cf253d412a8981e42d71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h662964fcabdfa86428adec00f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2bb8a2f1f435f81f3387aa17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71effd6ab439c7060e0242477;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb909cae67a2826bf25f021b6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf88202e0545fc30b705a2eb8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb59006c3981444001aa2edd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb993d7fe589b8825d96d46379;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6875df088be5963fa9c4f901;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5bf3750eb912205a130e673a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb29c3859f31b1275db1014ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h553199cd29d6e361779f5861d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d0df9f9c4302af430c407b2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64377380a4ab8c3783ea6585d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc22d6b2c1ed8f279871cd20db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hada8525b1c557977b69d9ba95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc19c7c545728bd09bd92c85e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41f4581a05ec95a60c4fae216;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h538128ea4c66dfc75ad3afb14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e923e751eaf3a57896ed9a4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c054a87d58afd7acabd91457;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e08ce994acfe259d21b6c3cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3ce69a0793aa83b4a7fc6306;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ef5177215568834cfdeec593;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he80b07cba67b48c446c622b40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef13776c7184d5f02eb199476;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc1bf5daf75878964c1cd683d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87759e3adaedf0b618182d491;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h373f3af4cdde030ad33654b3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1d81bf513d41a53b37a8c513;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9eb398855b328b8bce16f2b4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0c35c453b94424e9447af0d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he702f0c49369c54d5773a17c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d1b5b8b780cde0fa87a4a4c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77f13c1b4cbbb213c8cf0d050;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60bf4dead7eb7428509941014;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf29102c2ea2e844afd868297b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99bbd9369a76b51ccdb11160e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11fe9d232efdda7895cf55090;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habe4f0cc98f794be46ff5aa11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7604df4d53d291cce30c14dee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3af63c04d2540a740a88d437;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h331baa632538ffeb5681e007d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9030c54034eca432abadf3bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9fc95eae89a07ed5a54c96b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6644ebf0b8891f268e958f4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64ebf5f94a60c800d0250ab3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9abfe797db5f7f5b23eb3281c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf431cca4fddf73926fbe61971;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59ae8d8dedd47c6bce6ef79cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1e52d7cb24ed61782496aa0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h756209aeb4da6d0a5a8bea147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ab64006eff90ef55ca967c68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2dad8afe83c04619b7f5eb44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6742c85d8b3f4a8798ee397e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45434a98b6a262dc5e1c7486;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7defb54096508cd977cc7862;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha620c93710650f6358f167171;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4877615aefd63ebaf7fab8fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf2eecb7f8a31f96679d3330b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d9e733290df05deeba7386ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38bbac5ed64235081e6d01e92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfadabaf3bab69a1f50cf20f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h677b7ab688dd6fba814c31bbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba963e040bb6671e72def7669;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc02db8ad764601890518858fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d701587b1a4b5410814ae37a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39953777e3e6b58da3d560c2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h416adc6578a8f6d1075f31d24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdef4bfac51ea3c0fa7f8ff24d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a3e26e259bc2d645cff30501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h717eca4157a5c139ac8e45fc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62aecdb5a8aba82a6ffb75149;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72cc17915bb7dd9cce5b62c4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaa3ca256a9ab10be2d728827;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bf17e55671b90d8ff0620c73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h199c4ebc822cfcf970623f496;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8c262da746fe5c4e068d0e2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23c6eb366d1c4f35d6b4db87c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb82233304e0b97c20567d407;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedca328e53c6aa6975f7c9fbb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8790af839e9507930ed235ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c2932532a5cc01238ce8f10c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84fc9bc785a36bca832806b9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha78f7303b300efc590ea6c349;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2806d79d5041bbd7d5b9c558;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdb9d71ce5cefeaa6594f15d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46cdafef10b3b14d2c1e92c92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8c7fd271a5f159720892322d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb50b4064dc57e57ace242c2f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9717137a2aa9862cb3f46ab4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdb73f0402eeb0583881da8d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he71ad4f2ecbc53069cc641e09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79d0f91d8ab7c86efa72bcb4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he87bf071d8425f93495bfe23e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h192a5ad70a35e3529f99eba37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c5526789f3784df061984c2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78a58b54fa74563190e2a535d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87af32319bf286f9591c45e3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fc0e54b9ab65cc2b914c909e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h101d9cfae0c5c20b1f9cdc2c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b4e2a68b5a67a2c0665b935d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4463df2fc66d009728eb30853;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3dbcb545b331f72ddb7b0a64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc599e804c18ac1c79e47c10d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3340aa1fe306e7b88bfd74223;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39c95de97ff1ad1b46dd7cb6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ad782089da50e32f83d495b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcebf9a9bbc267affd3d9bc6e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h262130953bbf9764d31a6a870;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bbbd09241aed21f41f459536;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd25776d44e89bbf951e4b39a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76a40fe0a4df04f378755ef4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e3629fb104f4e5c23da8ea09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf82d6475f242e9e3674a75094;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e0036c6be236c339241f8f87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1264694318dcdeb9640318395;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed8b50e6494a61f188234be0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94aec802b7726b1e6ac78c664;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf090ae0eb8d3e31a564dee058;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd409b78c996dbf4b33952dd6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc34c7c3b87621d9152cec7061;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h412f51c84489cd8110de61819;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1654fcafd97a678e67ef59bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d93cfd739926ff863c922e1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31549229d12e26e0188a328e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf27b1ce84ec35079bf103b0fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcb3d8eb774fd19282ab8e1c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76825f329961e958eed04ad99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27c8ac92ce89c5038dfbe601;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4316468616a161751d3335ad9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5fb3e42945c9cdc9e3022ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48d09fccf5c38236e0765bd98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c0e50627061d863219597783;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2391f85158de4dbd7cf431793;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha02d2cbc1fe15e88cba5e69d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65a137c86f3b6faa2d467cff0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb1d6e728aae0461a51180539;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb57584764f553a9c84a54fd0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h990a39b083e77b23012a5bd9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87b1d0c834ed05eda9c391032;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70644f399af06f136a7995d26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54caeb6b69e83f859d9d8c3a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70605bb8858b0a7b3fe4440a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heec7c902eea037de1c5dbab72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7baa9df70f81772c47af46af8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2a0ea270355d6e5750bb59ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73eecb09518b976e1efe4c336;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc39d7fa17f0c7656d9b84305c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9e4886a605490d204ab9c920;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fd11474cdee7b0709f75eb96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0facb39b244a07528d806b7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f76cc3daee4de26738849660;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1375f6f73e710339f2fcd2d57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf311d908909439b8f9fd58748;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h459c2e175dc226369f59f22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24ae1bf0cd0873ebf4cb9adff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dd9648fdc3b73fd225001bdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6dfba9c773f57c0b56bccdb6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2387fbbaafad1cee47969e7fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hada94fbf562ad07a84e2825c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h989f39f0736a3a7d4c06ef6d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90e4509c35ca474aead210507;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc757253076bf78b4146c35178;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadb81ea97b1f84bbe283b225f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedda9dc5c0a87b54c29c176b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdeed3245f49255cb336f1761b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h598f6b82aae613c5424999094;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6facaa5bf86972edd0cfb67b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda00348619084839c9d23f672;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2464f4dd26b0904fa9d52b4d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ccb88716645a6761ca9241d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4279e26b9277cb50dd8889c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h354c8e5f97ba3d9b6b7cc9c8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a63e06543f88502245249a9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h457d13f09e07825110ef51644;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c5ab055e3e6073c7cb178055;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h774186f82c82dafa1c49b23b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a46115da0073fc93cd5af5f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bb55bf118d51ddd71313c95e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bff7cd91b2d76691b0137355;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f8e78d306cc67d9c049e3f19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3907abcd907c7acad4c56d358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b83f4c728e513fc2b89a5bd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he94d9c00f4945c67f09296a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h995a0d5ae4a5abd83672a50ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62a98cbcd55ce6db4ba5fb088;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a466dced460ea0c71ba6a026;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h376022d80cc4412b7f414e474;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbf8851f2797b34a2ddf65479;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habc5d336a5762691d8271ac8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1442572292e93d7d087f53b51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7fb019dfc2e7380c9532e6d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0c9dc975f813635365c10e53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb999d9a4557179ac96bf7d7f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h248e983b7bcdd33d71ccac87f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h482d6d97ade39d9968e319126;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29e55e18f405f406b0295fbf0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h587d22c8f2371a94ab2dedae1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ead8be206e9152e5f81a6a00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7daff475967c51a7538cb4465;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7972752790bf593acfaf922da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b88d41917bb015796d281a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h291f1afe5fa374659d6c0389f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18f64a637f57fe6524d3375dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb59a36723c7b54d9201810468;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97d6551c2a90c76347eecbfb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60bb36300f3f558969ea85412;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f87a212c32a3df69b763ccdb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c975cbc33d14b15d3f0d7456;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f7d02fe724962d64783181dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bcbb8d277c96911ae05c8a61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd08edde238e5cd781d84c921;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4956be23dec03daed357f065;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h594bd268fa6a8158580db45fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9930f3c3b624c9a8eaac5ceac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc54a65b8ded02abc3a0284ce3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa53bce4f0c3824021ba94d03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77855b5d3f8da7b6f9d4c38ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd35b107fc4f6cab25828bd56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ebcf7718f97bc08ee1b2c0d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h375dce3ed94de1c7640bfa636;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaec7409fcbb9e9df3032154b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd06cd19b4001059c917de383;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98135519d710bc2df7da4cb06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a4f2f94e3980a455de3a1125;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e1f6748a01b79ff4c3a4c575;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h775df65e4f701ff08bdb558b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce85e50bb0058af413d3319dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha967e90121ad593f3e28f2c2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b9edf6c84b9dd1306f5afeca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52c24a7a4255fbec4324d4c5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67dbd8eb257f4ee12d67b72a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92a9beef92aa0d70538f782d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80c9842992dd988f875edbd42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e36f9bd5d7ad7bb484ed9569;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf343653a006e9a123e302307;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80deea8185648985a8aa4fa3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e44294ea184d770daf2ada4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e63fdba4a10f2d3de771602;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1518168b65ae4d52c76982682;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6ce5efb4fff29cab65025725;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb54898c7914feef03d8ffe74b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc40beffbd12e588ee115aeb71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d1d4e59887233710d29c4dbb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5f6c18bbce2932cfbad6e0f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had906ebf4120525674883215;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb78f7bec5772c221a74dedc52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h434d80427ab7ea56de1c2a18e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5324c8136b422121cdcfb71f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a9c377066262d9bcaf0aa36a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafeca9d0aa18420668f1978a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2a5ef011e04ed964361e816f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9b92cf3b2cb818b3dd45b94c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h664f2bc12f4019128c32d4192;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2e19a4ca9325d913f1afae80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cc11a2bb18ed13e1b85e733e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2eadd3d8e087b82995c165a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35a757306b31d5e7910fdc2ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54a096649d95bd1e203e58184;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h209d027c1810facb1b9caa5b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he18fafbf28e31e745bb470b46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34dd93faf3fe4a82f647df7c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a205c1743980ee6c1ed16d04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23f230f3146f413f058eaedec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h220874313414e8fa4b0420e3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e22a848647cef73c3625dabd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8832644dc481b34ba0b32a4b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16faef0de80b2be5d0c5de15a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4dfd9907180fc4e162370de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecc5bd348c678278af66e97b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18176760f5d349f40aa8dffa1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6badfaa01e1b4c8346801e8b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd81acd7c98e08b82619d209b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc39f5cd2f55b43e41be48ce4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5398d214a743b0bae84dcddb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b706b859e521d8690abc7edd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ad78d50961f54115814539f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a7ad5630f1c3cff14eaa1502;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a7039fe2dd68db0ff8b1b0e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf303abc013c5365d777a6889d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac1dd12b2c01a9e7e1689381e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ac5c643c685bc10dfe954c4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2799455175233016db6a60111;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a32d7ec53d20f93c96a7e493;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b473da28526ab65171d2722c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5840bdf56ea0659c4ebb56426;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf28653b554444ba4905ebd403;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b11bb731727e30792bd3aa09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8b46c1df01084f43e1f1566c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb677f162b31d9ec49b26d7be6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8556849de151c8dcd4f0588;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1dbb4698c514c92038a5ec82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee6e8978e451985c843a1c1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4768140b739f884a1295d22e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dfdda4e6c9bfdcff9b7ebe91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfee8381285b2b376660305d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f2756cdce66698c3fbca0b29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fb2bf9e7e75b903dd7c2b93f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h978dad5a5cb286e503625ece4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88d30c57033db2b78cc744d20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h308d43f52f970e268b2f05535;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0dc51cec6d1f22f98b0a37bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2a956286676e3e71a717c264;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23fa79ec1bf68e77a4302c12b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4669c51a325acda7a8c3c90a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8b117675a06ece7a2059fdfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ee9f1aee2a59b3b8b454bec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfafaf4f4f50967b118eab6eac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7675c580b11a696fd55f0332;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd087bac287822b18bdde5e46b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10eabd8c473da2460fee898e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3a7adcd77b4f98e7a79f05de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20337968de189e53f29ce4e03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb50634d5f353ca6a45aa0b762;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h766f0f41777da654daa9a1791;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e64f7bf07bd267d8e1843b11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e433f839f8bb6a3ffca2977d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10ecb37de2d4097ec4e4b486d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0ad93150e188477b38387ab1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc356a5ad73092ee166e1aec8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc8e996c815c7fd984eec34e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08bdb5b19577163624a6cbd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e0eb4388756856bf31d2a9ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf8101ae1e825df240370e1e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d629086a0d9012638281c062;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67867a9404c54a7f300fa3144;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha355bdc2f1f498c02d83643e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd82c2f4b9a818821c82b28ed2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c1600adcfb6316bd6032984e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha95d1f090720e09841ec4dce4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47bd40f49bc41effd0c4c54dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e26ffb4dc0a1377688b24e20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hace258ad91fa450e200af5dd4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8e5d2ccb249fbd7ae075972d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbaa49f2a8fa39d763c4c550e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb34122a114d826b99d5de42ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c84a234ee90e52d05da86882;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h999aabb0a4dc137a138d0504b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e24f90e8ebf6c8b3aaa5d5df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48b12421cd7f94a8e743a8e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1cd737e25becdcb646bf7a49e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a0cd78a8256ec177f073f2de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haac280638c7a91ad6ae6727f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2a659ea18e82e4b7fb722918;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7c26fa6793af99552187b4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7845184340cb742f0a72331e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf53daed72e396ffc2cd0072e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a32edc917e252d21b955e5ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91d2b3d62803cdf224abc6d0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb265b4ca37fd213b4ca366d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59b0c5e5e04241c27f544629d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57aea9f2ce66ff5f21f73125d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8ff9f39335bcf488ac9d22d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab7be36b409e7c2321d22e419;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ca71cacbfa99b04cf89e2957;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58a64344fa6a8ea27067a38d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h190c98e8f08769c0cb3f8ab29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb74511ed1c6468bf1518d0a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c2b878ab4fe2002f570924f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd06ce53adb67d3c9e80d37d88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h839bc058357f5304939030b7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67ab252a46a0ddba8d3c904e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6eb5ebf6fdb76241372395b83;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ae8cbbda4b7a028b9361d65b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e62ef42577b2d496d03f6060;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h190a82ad11b3b7a5da2200356;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bf2a647617c835c5a44f2de9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ec252a309ab5bee7e3538f27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eb8a358e34fa8dc4aff0d388;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he92a455a13021f3e449b798f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee59cf4cbc50ddced8bdc9af5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h936786c1ddf68fc00e81ce655;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h198213634439edce0795ef610;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbc66f4edf24611d2766c4d18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16ae20d5790903f05a7cedc13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66597202de037947a885c481f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11052d2ed97a8777936ceb35a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9c013869c20adcbbb85b7540;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57af0e29529f02e162e21a41a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14e727a78a12859977d020ba8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe00817311cbafb65f26b48bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc90a36dbd7027f527052d98ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24c807269595b34ff9ceb2169;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h889a68553ea5c3523e3f21e0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17637a25bdabbbdf558ad3a97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha20665a77bc37a8e1cfaf737;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7dae28824e358cca7dbab87c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0b4d1e9ddaf1790e3635d553;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dd20bbe75af267214295155a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40e2d89cc0e28379ccd278493;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f4741489f89be74c4a5210a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4e54beda16531b889474585f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9376c81b7cc4a896aecd9ff2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf22703c68c9a56ef7a65d431;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8f9101f3035392c986877183;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92f516c7cecf96f6b606e312f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5c2e9560d0c12e47842d5637;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f95fd1599ece47069f3c26b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc65373789c112c8f5f329e47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h821e62d6a7c190e5e2ad5d612;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h119beb3f44dd0c6519dbb72a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfb0a2d9c33cab2f09b911a6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1db2c0ffcad55811911c9618;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d2be642326baaf06c9d11a7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea71674cab00bdbcbc0bb146e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11bca22a7d287f14b21c8af99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27ea5a2b222dc959641a8c996;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44564eb41ef7263b6bd25f48f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28ba9b054dc02b3140b895aa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf96d8aa6fd96cebb12104c1f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab98d2b1d2cf2b06413a72e8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6319184a0815f4cf7d0aa7362;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee894443902313615b8d120b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b028d11b83cb143c50a81272;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h189fdbfdae1fc2247bd6594d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5c023ac0dc99882808d378b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e482cca33d5a1a4c0caedef1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha961ca78a9bf3c3b475c57215;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cc9bf88ff0dceb8403e5ca7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f8dfce7ab701dd143b642074;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbef571c6e0287305bb83e6924;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h971f2d0a75c1e2da4ce692bd4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79493c06bfe925ffa6d827602;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h213a9c034e2c6661194888a70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f1faddf9186f00e8fae536f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b73c32036de1c52401384281;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93395a13e7c6962e92e77d182;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7ea23b452b0472a5b316aab6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha37b27622ab550ab8e98bf080;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6659305f2a714c79693f109a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce979d16eda60245ded28a64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0763d9f3bc1f420f20198b58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cb59e61420b6b08b8de8bbb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52cb04a2aa0687f3c75eb86ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f5132f44233d1d12dd17a4de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe11dffab31658f2c63619057;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56f6275cad1ced8432ddd6459;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h916c664aac4f57c5dc06e2bdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6406f43e844fb66025fe95ae6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a58e0a8d4c18807df8721c03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24ef303014abc63ad6b719ebc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98b9327477d2568b391ebed93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34a985aa875e9fbd62aa44bf6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4a6d6fef5301861c487f4bf2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc07e5bc0f21a6bcbd401fb3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74092358f3ed9b840ec45d7fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f2adbf9b44106af868230698;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h701d73b9b2e85eb7501d028fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde30d3816b4f0bc803d26d586;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5d1e220965d7b78a9e50787c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecabecc69fd8b178efb3fe341;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e7695fb2ab897d15266ab58f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbef95bfe9334262602b3b166d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d303cbabbe8f6fc5865e64f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h966bada3ce0e384629ad5fee3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46566b750174dc3a7ecdaebd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbd8218ece23fd6de57a28c4c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa4ff6cb2de8a1d48a0df3262;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6f41ca1830c9ff1b5311b01b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcc64b116cb7bb962a7d9429a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c8e2491139cedd16a0eae925;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8035ac63be154742c9717f0cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h481c92f4cf7e207a7bad73776;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3916319c11ccc809e3caf56ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h488c25ab37f65d7966ceb73cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf38e45e5a6a677d1b7f69e38f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcfba0a9d8628ab00f7e5d35e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc6bda654e157e9dfa4f292a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd7f07efd185092998b114f7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5d9c7e29771792680989e103;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf829440039f0f779c0224586f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0e4279516ed20c670f872640;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1785d87e524566fc0f15672c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a1b28b5938289040b079a5f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47250b5718d9df8db70a31be2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b745356c490e48d6cba6042f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6ef7cb6b1dfb9f0a6abe78a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee1798dc15aa5e062c88dd246;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69fd99850578acbf35c09df95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h165bd7e10b803a0580851cb24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10043a0198b5e4bb6e1d0c90a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h841c1025b7df1d17f336c4529;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8871e73691baec3e11b3fd644;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4022e6481c72118e7961cd9d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2ee47ea5f2916a7abc3a2d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ba0b6e21efa6b6283bf41335;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h346b2931e5d7ff9c61274ea57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24be2d02266a2d61a620bdbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h201742308be9b2ebb2839e49c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94c98f0c6f34aecd3153d36bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd71cb8345db7582a98adcd4d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1142edc7354b0ddd7fa56f221;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4005d87dbf4c59d65a4a7e333;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35cceb8c66bf878b57f797c76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12d9c81ca7fe6d347ca7641bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd12f4fdb07f83135dbf3204ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bbef94e7468f7ed953cc44ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1077662fa4adc78e88e31072;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc12658424f2fc949f0dbd5f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ed13e274c356f7e750df2224;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d61ca2650cb5b2d1a5e8ab47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h940abf9379e8a141dea6f94f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h475cdf0b8e1df857708d40e3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ddf4e46bd62b1482887971bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb711ff409d058c37b441c9a5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8cfcdc256939035382ff1ec7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h430b169671618938c6e30b1fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfea7060affc4033d324b7a02f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6319fb85c8b0a837253a96054;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae80bf590158346d822b3db53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc19420b346d9395864c415c9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12a97dff1e0a2f525fcf06d5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habf7df2fe6c5a0e836bad3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a48bf74d51a03010e826667f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e9cc1b7fa953658436d024ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cd70df65cb088b85ab2bd656;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8079225cdc0c19bb5ce99bf7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8387d6ea16195baa97b540963;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h819edf2320f480a975ab60d74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5475d8f5908f3374db6fcb1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45833c6df47d311e561963e75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdad8c39824d55b04dc4b29bea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5769eb9eb3a29c5d1e585fe7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64673b428ab63a888584fdeb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21a53118b17ce2fd3f70399b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf15164dbf667b67324e55cdee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92592605599c8481a18148c09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79e30fb21d1a1eebc4b4fa0ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd94c4ecf287a5c430ad942798;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfceefc731bdbf5fc5e31c5e7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9723f47d4f7c3ccb51a2b8a9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaccfc06b8cf7a4999eb3cbfe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h276849fe841524227eb398d77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ff628ef718330c6ecc8195fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49fbab01fcbcee93be74033c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5e3e7434d12c7797722279b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a13961ca86c76b9313aac326;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8baec4968d6ceb5eaf72b3e77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h110bfae95b41eb74570084e0c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88d9bd26acec6a2d35bcc02fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2899d9b3f95b972f0f208ea4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655299d3ad9ebf763ee1a08a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heee4a3c73e0f3ff19b446dbe0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce210550c0ff1bac90a5236db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h502e2c3635863b86f2fc4b22f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5602d60ad32f31f670ca1b2ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd188a6fa2eb1514e1b12c08f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1cde2f9d9f3ac4d10f13ed41f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8a5b4786cc9a8c5cd611f8ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc23a6e2072a995b60d7f4db7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbea3968075f853cf7e2752cc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb974812f2899c1e549536436f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha233b25808b096a838f7d2317;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cca8f943d512ea4a9462579d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10dd68a6eff6352eba6e816b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dbf24aed1ef4e8f220d91942;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee47555d702f85d66ce4d05f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b81653af0e73966d183beeb2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9131528d46ec22c44baa7a7cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb955d157fc2c04726c2e7a6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf35fc9b3e683913d74e9e4acb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85dcd63ceab25448068a77686;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a464eab29d297ad383bc36f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he55949f0e6992ce4c6e8844e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h276781eb377ef707ec417526e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38d0c6d8899f8c0a61485bdcb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c0f561de0fffa3e3f429aa47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18f8a9de6d2de5db623904add;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h804a66ae259277c9d940a85df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd371c2f83b56027224f3928a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f1af693455552cd65b37d9f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h492d2fd5b0077dd19205b2e52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c72144ba5b28375966162730;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd0bd91fd2654e1114d75da27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71d95b599d6b48a15e5547729;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8abd5c5a5f851a960c33ea87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdc7d6fd9f243b328e5c567e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h451584da0954e38cf60b3e194;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe60c8734153fc0cc533f62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc59b8568359ba49bb78d2191d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74725fa4446a31666c6990f63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda5dcf1671195136ef05b5f40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd90b9d0a45b2936fe73d0467;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2ac44cd7eab6b3e52fce82f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73d5752e05375cc64c296898;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbcbeabdb3c38dccef9453aae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7288548eee0655e8f29e13d09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h669332731edd5c5961f818a84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78922354c3feb9c41ea380abc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5df9a6139cf85060d84b0b896;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ece2954ff3d41951ca1e110a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf49bd8619c27c32839a0a83f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6801846927e0d83ef21ceff0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63bdbcbe718f0d8b68a342472;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe4625e83d69b7263c6d7676c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcbda353b4dbc9e63152a9b8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he89770e5a02a6cc9555b3805f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcd3bf2e190cc733f1134f378;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88b9ccfcb4ed8f91b4fab3c2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef6a15057083409d1d31e87aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d5c801a297d9fb1b841d8f35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc3f013b669609cb80f76bcdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c2734eb090c3f89526157670;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h536e248664ed164df5c0130c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b64553e7719ebd06c61835f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64720337d644e864bfa71a785;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4efc72513ce14268c9be5968d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a494fe4086529265721b3827;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42ba5695afbb36db8a03baf7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f67791dd7778fd1da1336e2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb06718890ba172fab19b834c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78e35dfe6a015c8bc4ed9b117;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7fdb9eef7b805037cd305506;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde438aeed79d6242a15db911f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c94e578fbc921e6c2c0b4950;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb4d7b6cd4344f010d0a6246a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b99c5d9d30476a1dd47b681e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2b139496e296756384a8a424;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cac6e3feb59575e93c731a6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h923d3edc232521070747dfb05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46749e04922fd0833cc58e578;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a1d0c3e1a89ae25cbaef3a5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d85f174c5e1472f383c5a288;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h770fbcb70d20771dfa272e78e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he449da7242de1c95f555bba6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11ba445a8596f2d2aa923ad22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eb9344801e93e81288cca381;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2853bac15b216dec04cf27512;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf08ee81513b0ceb09476ba2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d6a9dd1e8429f991e994671d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb39335905c0212a0548a3707e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63a9b39fb774e49af1ace59db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdabe24e46c73a2f04fc6b207;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f89d3b46156b397561eb3828;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9aa28d4f38aeb30c8cacaa3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc69baf221111c474ee93519e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9a8dea6c88138668ecde96b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d7922d216d5dde5c18d421a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha500f088ac38018ffbcc9fc1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34246926e1c9600478e2013ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae1622bd4d0dd075df0930fb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81497df5a80d99303a8032f2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9988053d34e3ac4c228a2070e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab38cdb1bffc5f725d867781;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ee11d88da70a82f6e2a3000d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h949698feb7311fc5cf5e1d85c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6570250921b8f2cace107264;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff7b00441ac51ad0b1903db17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff0f4e2ad59c9d985619e6897;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2933a95edd3bc2b8230ba289;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6da9411bd32764da65b1850d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h295b403789138a17a58f766b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h571168d9548b4a605ecf4eacd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcf400eafee1e4df1bfefbb08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd47890264b7dc09db1e31ee3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12660492e311fba0a61509e64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb0dd2255b619ced13cf6ce95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a9ffbec68fad94aaa33122d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ca8fb0e6bcd008fe65e6a5d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h887ff2790931383d2e20e72d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he32d8acaefdbd06397715ddf1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h140f8bde61f7361a2d4651cc8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2aefae4eed67c6f7e4f53d4ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cc2e699d6db1882a49283aa6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba2fc7282e93a6a42c24884b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5bb0202ef8c6e5f19bae0902;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h831488ea4ecee389c260b6b8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h904c4dab0b334a6593ecd525b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3921a40dccac59f3af8e0e1d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee490fdf8ab8acb6ab84f4937;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb14cd743719cdc745a4bc228;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h920ad513ce37e77656faf9dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hace914a13c910ba79380064fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb396f955fb1102b2787e183e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e5031559ce03342686f93902;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h961e6dec44af9addb8cfc3fac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ab107bbb44bcd5c6ea094b63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ffc2e4f98b49732f0fb7b22e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60ffdda5292d1f84ce70fd256;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a94201882fc3bb5eac580713;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae1c911c2a56f804810b6092b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26332a07bc9a309ab6e5c525d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb78153758f13aa211b5511132;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8482998de88a5cb2895d3d856;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d901618c1603c4544c2964ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18cf94203c9c4ea0e335a0560;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8bc9b583a990fbda42bae9da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf32357414932af30a3fceb6a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h420a12e5502792b15003ba8ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e319194fc82d434c19298434;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54e263c902e25a5c4d75ad072;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63e941f29c22ab960d676c03f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57d4d5883ce2d45cb26feace0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bfdcfffa3d403772e566b5fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30ad42f1acd3e50c3a47302ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h278a6d4ed143a3fb383ee51c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a73499364f67e78fdfa67b95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h563cadafd53dbad8f7d39d35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6b1c4af994ac4b91d6813175;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b2c2b6ca5e58d419bce6cbea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7640c7a6a3e964e245cb64528;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h501fd3dcb13dd8f2aab998174;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76b14fcbdb4c4c616d93991ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc2a4c3009673f29c70d26c8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55b1fcf2596a8c4dc3645467c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcc4dd91e18f9fc301b06f9a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h608ac3eab1331c749aaba845d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h611a96283e1ae9041fb255ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dcaf016a53597ce186e5a2ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0f7d0078ba9bcffd23b1bbe2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e9017a9a449f1a94329a59cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e36033bdffd45fa6618dba71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ccfc51bc4fc32980a25bc126;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3af781c0a77d8b27d23f27846;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cec674401d4bbd759ec4231;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67e10b2b4f2f09a5db857e9c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha79fce7c2fee414b6fb7e3792;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h719237c9a51050e3b44ea1210;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h998423a685410d7994f16a0da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77650e2038a305b335991bf1d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ee7b3d61e41052f09d4b41a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d0d7d0e6e228bb14d1c0f1a0;
        #1
        $finish();
    end
endmodule
