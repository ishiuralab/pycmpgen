module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [26:0] src28;
    reg [25:0] src29;
    reg [24:0] src30;
    reg [23:0] src31;
    reg [22:0] src32;
    reg [21:0] src33;
    reg [20:0] src34;
    reg [19:0] src35;
    reg [18:0] src36;
    reg [17:0] src37;
    reg [16:0] src38;
    reg [15:0] src39;
    reg [14:0] src40;
    reg [13:0] src41;
    reg [12:0] src42;
    reg [11:0] src43;
    reg [10:0] src44;
    reg [9:0] src45;
    reg [8:0] src46;
    reg [7:0] src47;
    reg [6:0] src48;
    reg [5:0] src49;
    reg [4:0] src50;
    reg [3:0] src51;
    reg [2:0] src52;
    reg [1:0] src53;
    reg [0:0] src54;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [55:0] srcsum;
    wire [55:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3])<<51) + ((src52[0] + src52[1] + src52[2])<<52) + ((src53[0] + src53[1])<<53) + ((src54[0])<<54);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4ba3bcbf04a65590d1fd7d9615b6bdc8873ccf8ec8d5327c5ef118d992a1677316bf3c224078623bdf71f58ec594c30d6b5331292896814254aeaaa5fc02a983f9128ce6679fcde56644e1b5ae2806be9fd9b3d7a63d3847a7b8c24a9b489e5d895;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3fac03a043b845b01f2db9d13ab502e934c427aa5ff476d763c064572a6a53b6cd3a053674b5194acf8d8165ac9dd9f9c5774ce6dc8f2d503fbfc104c77a12f5c48f03400b00988f98755ada52b772ca7c226fabfb58f33a50c9a9a222d79f43833;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4455831a2dfa2c6657becaa1e89e5eaa1af40eab8a764d80756ea1a27c859a9136d36d8786a76dc0ba836a7264ecad3d09f7e56e6bb514bbc368202909736fd3b3a183200f81498a41ec8ab810dcd83185ba8ec2c1ddee8de617ea838f7d7f4c5b98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ce59b9c0bf90bbdc9c2241cdf1b211ec37d618d91c235ec80cf84332c04c2689777a0947c4dca39560799b2d48c3812764e770a876d0b0f14ef0f6e9bfc60ded16acd83ceb5b0e26daf94de29674286bf6309581f6fbc08f62455472ca8214d697;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h610bda52d89f915160e059da491953d34ce5668bc45790620fe868175b7d2d04580140ed5f5de912e4e397abe990f50b19f43c20804aa8c17f3b3d60187ce48e4b553e14670eb7f45ef0631419241b6ef0936e4c002026b7c06879bde5d51cc49aa6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb03e36a823b060aeb8c63ac097d6990905d8262403c78f7d9f59b14ea355bbf2fecea94c25715c35a70ac7c45f07e3ff1721669a09ed70c9faa508ae466359085d2c5ac430c70c3d97214ec47cfb11a38f5e75fe8adf8cf8a46391ee978b8d933c96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea186958c62a20dcdcef5a1306db6b145b6572e68bd680711f19c692412245ecd00294ad98dcea47195aec16af16985343467691e62cd661c0e761fb548f171a882298f60129355bd63f253f0b47ac0a764e34da2a33611a619e74bc3be730e7d432;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc40f98b966e3dc1ff693658ab6dc8fb4bd389a8e99a910496fa03acd9a17fe7af0a893af4e8d1e65b1f3960b61edab6eac522bd1e3e533c6881f79788fa0ce3b6bd1216ec2993fae0a76dab7e9c6ca5f5ed369f52ea62194ae3864016b25f402c502;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe50a4e6a3c0501a9cb6d757301c74c8d3d617c144436ba9f59985d2c240c538a0c125fe20229459e049e3b3431ddc366ad68dee6484a52f69677c6de5d209467cb27502835837c5197fe74a10b1ae6af3c7d3dd4b4c8a507faea070d3549356d6e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he407b777c3aa7e1e7f5a8561fbfd78e479dc697a5a6c102b46704b115c822efa9a784ad801017d7d0b6dd3d3290feb1c6830fdbdf4e7aa90ccbe22328e7ba0b4b0d7e00a4dd1aa06f67be3f141b8b1938c8174ae9e7b6b78ff52057b0f1dfd8700fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6e853dc6d4431d9860231374f912c540c7378c8a9bc691627071e13fa1abad8649abfd15ddf9f4fea675cd829ce546de5ccd7007c6445ae41332a8df474264716bd217668bc65af58e5d8adee8850e1f914dba589f1ee29720957ee6b5adc95fcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82c851d25865f302dc99e4245fa5ab02f5b639080e4b792d953d8c2a42a909a7bc510f64b743848e428eaba5264fdb0c06094acde46f36fe5f74048ca5521d0be5075483929f121078134439a52ead43628729d4811803dfe67f2c326bf53c01af71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1abc357d0c3f7979d921522b355102679c6db4cdc8ab1ec3e36d2f3580bd6c7044bf393619f5a2a08ea49099cf3968d9db627010a5ec93a812b15e5740cdd93b623ef5ac37cd600553126fb09b0d8deaa0cd4432566f36ee9bf6315a0ec0e6847073;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd75f7ae45bbb47192bda5729043fbf5ef2b7c8ffdd8ce8d94d70085495ec20727f833f7f676e3a0199a9dd7dfdf3a28799b4887b7d84d37658e3254b83128ff61c51e32b2d2cdd9fd207a400cee05aa321744004bde89e46748fbb9f6fb03fcdf4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h619eda5b992794e8016908067efdc25c6fa5d5fdb2211d36869abba58f7d383ba87c3b76703a011b3f5c45cc432d133c3573400bd9e40814abb1136eb91b1588cb42748d18433d07cd5dce76b7cd0e6338003f144d978a1fa0b05b1a286b4effa9ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha51a4d36647b1a49ce0e0de81ea61f196e5144209e60ae743b8c0ee90b152b28217c60a52575aa5899ab76c8ab313cc510d07778c686892c5721acfde7dc59ac54bca60892a02bc4f52d4aacbed02f7d47a942d7631a60d09ed44d9d9dbd56f6142f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d661016f5e6085b609666549b1025a00d44b49bcfbbdf5fd4eeef21e9a1d39eebfb633ae8d4b29665cf46e819557d3bfe5f6b30914947e4992e196e438ca1389e9c941706fe8ad94fda41337aed7624a3c7e29800ef0f991dfad5f73b67c062b768;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bf61faef4e47c5c56c6a96d9927a17e31360a07642caedf199ef5070d1851898aad3c0c8aaa5ae7f3d109d06fbc15b93fbe85fc16d33d771f6031341315b8acde1bcaf5e2a79edccf02f71a2e6ec7fb4a49435ff15c44a78d56e685f807467bc768;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16583e872c09d4b39cea05139869767fa84207b2940750b9532e0c69861ee65593c4bf88716b517f40f96eb82caf2ca5aa9256ca87098710b0415b4f154f9eb82869b275cdef5ae2f9502e913c6286d21f8ec3806b7c1cedeb51e6eaf2ef70433a9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76ac2b6fc141716454d7c647de54b90d0fdd85f304b2974b2182aaadd67ab833a7e9b718ed6a574bb50cbe548bc27a6193e4c8d4a5748bcdb1b0383618f0f519eb853873598be733eed8090f0a3165edaaa783475bcaf51b13a7ad731c2cddb05e36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb16753192c95aa55f4d867c3589e5bbc9989cee5a81a11bf28688620b3abc7ad2f53efad5b35f8e2a5666c80ef991ab664ced1a5fe7058e983802ca64e049ce6be2b7158f3ddeb0213fef175e90ebb4415ef07c5c9348eaaae6e4a60024ebef48ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dbf5284a0b59fdd19017cbbe3786016567854a275210715b7ea612f17606be4824f61ff627670171f18f3feb1d52270699a219d7f04cdc642c633422a36a799514565e70f3a1d6b74de0bb6f2816a48dccfd98a39bc46f7bac0140357a3376fc0b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f7800f427e79215c2c177fe4e446e42a82a633bf0f8f6dc6dc83d0835143b4b4ba89c9fcc9a65f1d27648abe055e229a6a1b13d2726c89812b9d04e526999e330e3d0da6be8cff6145cd67a8d7f24e350aa054e983ca7d609a71c84453fe156fc44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5cd7221e6687f0c2714fa9ec2b02458431eaf1de619b7275d1e3037d5e141b2144ff05ceb4f1c984fc3d5a5ba497eb1acf360b59d6a48a65691b3aaab938419d56df511b461cec941949fe853f4d69c49a14d64446be1e638f463e433c0ef38ef3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18c5e92788cfd7be150b5a066a732cd8673e9731def061c31aaef213c57855f13edb2e974621a9bcae14552336aea8842e0d94ce073f486b6bbd3ee6f358a53d574d222beddc35b4990007f7e4a36c889e04159b8b2ebabdcbd21bb4acb419f147c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c92c8f7e1fd7779d4e91cc6f2130fffc670b470a835235430cdbdfecae41ee65335e19977fbb9197d466de7daccb0ee1b05021bcfc67a1d5498ab83637b2236411234cf3c0bf2dc6e1b35dfdd80d12a70311614ab7cf1753cca391600d5318e340d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb41a229646aecc4c6837d3830c7a0762d4ce339e5d8cc0ece6dd660b95a37b4a65daecf288f0c0b1392a71299e84f40afb55550bd3416bd290ed1f46ed8be3cb978224dd92595fef8a00241dce8105779500030cecd6ba0b87c38df82433ef4729ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h315a7dcf171f1a332bd36bac239d06f8ff07278c604bc33e38dd75744b83ea366f66681cf81e00c6110c8a30c85122057f7342320ea5941a6b180942e47077091a6e1fd2fbb033663e41b4a8e52b66aeab6f1ed95a6d7e9cc7622633cb33dfdbe258;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddbe93f6b24adf7221a4b64c8899a08f276de838659b11b531a9d8be7c2b1cab3faf7b72672656c3de182b4c4fe652701ed685bf11e938dd99f3651c8e0c34959a91281b3a7d8611d93c47e3c4720c03b5beb0a331b0e7d4a3b22e1a203a0dddc673;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ca9e7b81086310e4449197475e9e3ae54b8c144f2188ffae68dd23444ad9766fbde9039dc995622f6bb8c2559e1bb8e65026c43c949e3ec5d990be10acda3ed447fe6855d00b4a932e9463d854e063658e78a6fc36df05b38980b55a97aa2f668a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a0f781bc1b029d0f27334770b159ccfe91e99919b56c7cea134fd6f4496a8cd9d70b1ad90b8dfa71fb66967a664f4035abd27a8a8f0f49e1d6f1a51aecb526fc1a07c2cb2e345d90f5ae6420ac7fcb15206feef183d3378203553cec904288000d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb1c16f4a58e82fc4fbb72bde662607e656d423eb35906b71efa0bb73bd809655d473d96af42028758265c998a8dff32200521c6779a808b303f96777efa4c645f3de2a04a2682e5712ac2a7ca3119eda960ff1e95856addf3e6b6c99ac0c25f01ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd573a6b440c5be8291262e96da88301ae490ea4e79aa408264aa0691ad5e94af354ac438cfda69eb65bfe6096add90658be927d42785e321eae9ab95203d4a42f95db369ea1323f6b727044f94a8f651938909c84112a56dbddb0eb8326d83e77600;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed78df12289c84f2f1086922304839d2bf34cef45d8f7c5564b65f42da51db6d30bcad2ec6b98e5c65b7442421cc62d3d41117a9561fbc739121ae0a7c6b2d689235f3b23a89b2eca1e320dd8a3c13f9687776908348e7c95f3ac5e1a8354827ac7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53a44c18709b6a46883dd6a13c619059483da9cb60ddbd00c220996d36adc82d726cd86c0d6002b399875e9cc887fff3b85f2ac479668fa3540946bcf7a8760e4ab6fb15af5b5c8d467653c1fbf25aba5e246ca38e33c8258fbfe222312b8a13f07f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha30701091b79105ced089ca4db3eb82c49f74b0f813e595c4a0e24d44006438bc322c29f9f5f639cf294ec37fb4c36823e2f88ff66abb924aff3579a5d6e9ed475bc63d1a16c53fe94d0839708f4ee8131694a6319832027580f0fb4cc8cd208df85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7dad8692780120e1099674abcf613c123a127a0c99c8f9bc8bc80ccf4762501ff8caf798cd4f7685d4fb304934fb56eed3cc0c629b2d083bf719309bd974d80192cd6515ba1b1bc2fc1e672574c869fabf027e2e667fbfe63ea7b6a916da53d6995;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h902070efde251d46a09245083ca7624748dacbf3e48df7deda187962af7ec3649928ee9a7f0e8bb13a1a1c26ee81f9cf31bf0b50949d2e8afc50cda1ae98acffef2c4d00f2239afe682a75c131afc5eebbffa014eb9dfa7ba1fd5d653a9b58fb4561;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9101f96a4dfcb9cb9f117b937057447b99afa974845e4cd135510f0898c116f7ce97398fdcc211fe779c5434fcbfc31449500d6234ba5801f6db191805c0383844c78baed160860ae5576c28ff414d1121fbd52176ed95ca7898877e52780718fb42;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e01e1e1f6f6be0d03220a5290a0759cfe5ae594ed6c10d24e1e3f111390fda54ba60c58c09e15f9d8feb80481548a8d417e4bf9f29346fcfecfbd1df651c9a8c37a1b2668f0f3bb9ead95abc448dc64c789e1ec150d8f560ca9c464212551d104f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44046d0460674062f23072b793947d6c665b91aa5650c4b80e1ddb7d71a502eb7080f00442080630ec7100fbda7492f985603e5311c9f516097fafe2a8120927f66883e9c3d59d53f2657141537d01cbf26a5bd37f7d8783e0965fe7745b61ac5e98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb866c6d1446e98034e7274a6ae54bed24cfac7e31ad667b4005feb3eb7a4d627c81d4002ac8e7b9845108e0cbac92348784cd2193aec6d690ec5fcc01b7602e849999b08f8230d649a47959863e0d069a25c8613f513639c784863827aa7e4f17247;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5526534a84e084e0f0d99ec5bf754cb3122d305b65fafe2e295c2c948fca7462e0084d2c01a6a36c2b5bb27ca5fef20627a984454b0017738e43e8080047cc269386ad0e5e01f88272d5ac7239d79d73b61c7056af361c74168cb776de3b99296712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f3533e927ed85d5eca3113543961a708ec3a0c8f32ab8b6598ca5e455329485c60a3c57510b27ec226dfa314bd5e1808f8d4bb6842138d2ea81fe973d1682cc3812b5ca227c4ba491eaceaa6f680658feb6105d9e6e32923fb187c4fcff662ccc60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2b5bf889820a7db8a6bf8ebd5fdf572f3a328ea199ae3f24a2f9886094cef29c84ef4f9d764253e331b078f337c5874ea37e8d23caa82cd7c6b7864205a33626691db3905f03481bd3363a1cb71da22fd9665f9a0fca5facef16e88746cb100e4e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd67e517ec557de6ac9f815ed528c8cd14c042decbf7f82c6bf1c2a5f473b1014a598654871c202a59a387dbcbd9f104e6946de51408e3d4ccc9dba199752f42bdc13ccf77481b048954646b508b46d0d42ac4f57a8deebe617867640b5acff81b886;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bf545af3562b1c248411c17061df0dd548cd8640b946fd044322d816a4094eb5b66a87ebadc822cb480ed4df9a2011d7a0e13409dbd3f5a43a344d479182f3104888b93ad3d4ef429a8bfe1d6833562170a3441fbbe11dbf618be5695127cca187f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd40531a5167ba784f4a5cf99384714da36aa16950b9e314af17a144ab7e2510a4d8fe06127afee24bca032d82c6feb805eb7e8a494a5d911e40f5811c0a4bf9e1a61610fd3067f4e2ebdc7f873336b11ffa30088e45a72ad8ec464f29dcf69073ac2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha33ac0184f63c5279d85af418bec0d3298c0a88a8898787150a7f019e9882130d37141268b8cf1aba5f63da8ae98d358ff6e1f535658d7b241de7340a915c593566da745e9a8c31624a4ff47608c1cc3b16f370a9a5077f098f6499c8f7bc1ff8ab6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h873267bbfdb9a9a7a80970aa803c4d72b5ba1feecd6237a6342700699d0be384dccb2f6f476da9c17d7bb8ea09f8c48807e0381bdf9cff2935f4bb0e4cb83190d4e96f2e28682e7d781bad8d737b17205fd0d09dbc6e30574db47b4382c473837257;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h507afb70943115a7d96264c6e34b9d8904440d52a82b44acd5128646ccd012cd4c4746d6f094ce919eb694aa3562b6565e15c2ba5b591131d6c7a07279f0c2e129552351165d277dd5eb89c05b388bc126ae165abe399a9f48ba52aab67c63e64cc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24f2e35d7e2728bd8f218797a73f053fd58e39b86f12687f822ca783f434d950be49201a1f426944d6c948bb0af03ffcb1aee89f4fc6f1dce30f1ae43118bb7dce260f1dcd4e6c3846d5e00ccd125fd404ab8ecabb45e68a81e5d41818296b36d40f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h951016220ec962ecabcc3f11201ff79554795965708ee8b5c17397fa901432c68feda2fc561818472140246f76d8749f7ee60d43b503b9b732599ec3073f2130187badf70b06ad63e8d1888139b6c965031b51c36ce6a2e324dc29de10cd0c122081;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f7cea353b551fee51d2ebc2a53c4c1c6f8aa8ed37ebc54b3d17da80a1f8eaa8b7093dfd43f9a4927b08625a69bc78e236af3477605b6c8a46639815221df103db84b7031aad9b4496f8f317d11c14d1130be745fca20e37552d47c746f2488f9369;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h134d813645313b8369cd81d2cfeff5944289a287429d0e544319593573779c2a039193cdd89d4a3d6851a3ef53ee3e3fa0b3098d7bbd3459d72daef3b730501ecdd0832af54bd0646a117cb3d1624a62a73191fca68a5b9d4fc014e5956ac343c583;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb16e685923f4c0197816bf12524abec9814411786e04aff8c812ae58c4601f695e8b5c2c4e2f291326fad3d8bd854da30b1e21b234d9b90d161adf731693eb808548625602e283d0eec07c63a838945bf3fb436e0c223f4b3b02bd1aff1122c42713;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76b1796f7aa5c1d800cb21552cc66aee092e0af57f4955ef72f173eb05acc5078e2f7627d2ab3253478e055224df030e10c2144b1adc8f73fd4e18e96ece99b6bd3275faae0b2cb3dbe2925c60e4a24fbdb8392a6a2e4459e83cdad6b9c4488652e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec104dce4103d9b0926fde7909aa162b019a5902932b480e589de23f06b5360eb826e43fbef3e41bc54cb69def37cb21b466d13e9da92bc4c282deacb9106a8979c5de882915a3e93049f597b43fad79fcebd7235f16e6905d0ff4187714c646ab5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd008efb5bf4eb5a1b678e50cceedf2550ecffcdd95fc87afa1fe7927b365dc437c63d60a2600ad73cd82c8c3cf235172ae1d6d4274bc1f1919850f204aa0855fa84f9f2a274fa5967e9f5a8280b6df631161490c4636abe62fb2c801a819d351250;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddb6750ab39b4e27c8b8d9a471d1a269169f62e0f76930af610dde7bf57dceeb49ae3c7ea196ff9fe109fb4541ad040f80b4e64dbeddc4978befd5cdeb60dea15d7e2afb95b44b4762ca3edb3725410f52d8ca63caa404f1196f2b57e677a86eaf7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f18890efef4971fbad6a301d5d8459d6eda612a14ba5a6da420a22bf8fc6d9eada4b682230de461fc092103eafecf3d27c95ddfe8506b8e781b8413766a9a2296054e9d198fa0f1ad420a3d0453348c9d6dca812fb947e67e1d398a92b9b8a613f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56f304ff7e601d3885c1669818ae7d3075d6a669f96b6a5ca21df2cc20089a39ef19abe74380e99e473e9ffdcee82841fc1b7e506a24006de6184758af08fdfb4a4cfb85127324f985a7ed3a184cf4e03e724e963aee8d9afe5ca7b7ef997021ca72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he128b5a651510e9bc26e342dd24c4dab93d7d17c750ec600910636da9f94360fcb85708896de254b9353c38c08d47edbfb21ad9b5cd599e54823082742b8fcb7ef7bf84a7f516690ea8d8f5c6834eae8043ecfa366f34674e75965812377ed0a3d44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h778f923b34ffbd24021d005f002fce48d6e7a5f3546f355bdbcdb357a37c7d8f5548897729175fcdf94bd9d9e50b9be47b90b9b56753d10d47d9be9483ee31a2184cbed1c1488932f714d1c3d217df68cc97f5637456381c86ac696abac819bafa0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf55fb6efb69a8f31adf6a9f34258aba97dbb4a2b94eab8bbde40999a3302a5c09d5c551124fbb20bb36a0816fab934606d93503e36df5ea4155a4821c5b6343d1755234ddf3ea13f20cf07b90789f5177fe43ce30d0008720c9ef19db8d90266e8a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f4d6d868cfde7b99002ff42dc538c6c57f020add054369adbd474439356861126804c0216adfd13b2a54fbb4b05aa4acf6b14846ea072efb30671b0931224b97a55d9c401bc25d43028a48207115309012cc626d4a6db66c29f3564d1becf25715d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c5c25279ee5476176cb809081049c372003c4e93102fd9e7f69c966579904a39be6c1ca4e911e5df092df862be5458544d76cfa4b8ef4e9d2f2a0064431058b7ffb0dd3d643157226e2cb17b00c96ee53e60e337cff753c689a5d612695d8cff33a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e66125bc19af7d643dbc639608107ce6275ab90d8f9e7536f7947be7c2cbdfea4c366197f31acd3dab83bcec0d213e418a8b0dd23f322878301d6bdb79f2b80a66be0979cc33696ff6c0a7478a042872ae35ef79bc62ec4c8acd746f6d604276cd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h930b201d9b12470753368615329aaea16a967204d251ebd46860faab0b2b0bd515bd3106396a0100bc127d5decf39819af82248ebaa620ec85e50c40adc705af1274f298c738cedca649ccb758a469bf9264016909608dd9465731a0bb48f2f4fde1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1b13f34d734b4335bc0fd1fe4f7067c41b2494500d8f5d9095e2c916c4438b5a95e1029f3ac95ae5fce9050635385cdc70218af768f17cf41d179c4b35f6e3ab6bf92d046eb5944715a7c78700946b3b8a4ff8806d9d643ffc2a97162c8a2fbe40c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65ed6d3f456440822bb648cd9ebd6f8e7ab016bf41c234a89813dd89ff7d149fac29d6afb245eedac1a2f71ef2eda0dff55b116a0c2e6a09568d2361c4a71638e236c995d8b9f8c2cad0c27c5157e058ae5281e3f00dad8e4fc36505a7a2c0ffeb1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b0221b99ddd2cf461cbd8c7ad95178ea936eaaac70dae5d7260504d6b606c03d44e4a76b1deb188681740b2cf15fe0cfb16ae138f5b48c355d84d3bc4ce54dc9021dbfccd4096dcea1c89a396894d49cad1b351a50525cad7d4b11cee21a364706a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82ce684ffc6e93db293f7683d55e678a5f487bf683b8fa09df37ecae4467e8e047c8db5f00156b7cc6ff41b729eff6d1819886a4ff636350b5400c87025b399fa833f59bc7c95ed17e990df87fc747e34b371e10a8d16a99ce1c84ca4962aab0e316;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e851553cbbeb41792688ebb36578603cfe86f1bd202fdf9d6b9cc9b967736a2274125113b9bd2f3aff08eabf5d613fde1b9dcbc4f182a4f1e6e7cf758647dec5075eeaf64e5442fbe6818c7d3b2fd94e67a69e9d56a4350ccfebd9993e2f31a2f36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdb108118dce72be02fbe6986f5c5a2ec730be696b13cb07f2383408f45ceca6746406b7fefb8e802bf33ddc811633136f94b8e31ee576be0dae9781a24aaa6a12ec9b95002a5171ac4f8302166ce11cbb0d1e98dee264cb7a167a65fea9f99460d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7e5c01ef547ea31799fba9d11fe3b8133e095e8cd5757aa8be1a7bf6d444c5e377b5efbeafe78a75046f5bb594f6ddc6dc8c1333b2d2005c0437ebecb2ffe3c352b0ffb1a972da047d39033e2b4b7d926df4324ebbe51bdecd2441928a2806217f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa5d4e0a78844d6692e133b5fe0ccb19be34667b9deb699f602e8bc5f69627fc1c3cbc93b5f3f2f2c3cf266abc7b20c6821b98c17133fd06a81f3e7c0cc31f3a80af23e3ce3f90745afd937a421ecb696f032137237b0eb34d0e9c58975fa756017;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1749095bdb65939ff4db7a2e438516123ffff4cdc11d326cd9de97f364c6f0ababb5b16c94432c82c326081dcff671cb667551ad14c0283dc765371985ccd3ec812cbe566bbaf56164f0d3b000659d0df1924a87c0bab2cfa059b3185a153c754fdd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h760312b7890bbf6208b380e8dc4e3c0b7854c492173d69e968705eff2e7d989ac0c2bb9698f359dc278e3bdd0518ad2f88cac946a7d5e7f81c17e281fe59a6a4488053c80eaedfbb6e336fe8ab9853bcfef96ac2b8131fb017f91bebd0c2d66239f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4837463f7d6882dd55226323ab4eb4d82cfaab34d2b479c179821b33bedaa2a3eda3f59cb8b06b301ef8832d0636cdb7511a12b680d310c672a14f183333b2a55513de838b3ea4355bc782b83cde50bd99bbaf4ad7def68b5b002a53aa96d6c883a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b82afad50eef33081072d3b3f5e3266d2b46b625e9439e94b96eb0a1ea4c524d8addb98eb35824dc59c690eff81912983bf9c05f1f557b5c85798a9f0c4a3478d7b3ac86b084ed3dc1a0fb8bd55a6e6eedd0f778c5744afe68c3e28a615ee0f07e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18d986b1c863ad3c647774952a50e14b9dc26b6a744ab5516fcc31fb24aed99b76c715c3c6c7e8a7b23d298541d129b9136a4f1b002983e30ccf6d825f0affc5febd22ec3f130324bc7f548e0fa567429d4f2fa312533288d5c387643931ee36f715;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7e6489172739d1e89b0e361193b6c33a855b975e5cbc1c6ace88fe3215f803f3e67a62a1b604b039a213defd56e2d1054fc2073cf92cc5e7648e102f1c8b5171407a10447042b95c49d7ed55b3ce563752e09597dedc2f5ac48ff7b32a054f0a3a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a42e928b4b73d15eab883529e521cd283f89595481519c73cf2e592a22f7699ada6df727895c1f1fca37022219f2ae3ccdd6c8541eee110515d85c1dc339e2f3dd3822afc8da64dbb8da05011a6a70cac7ed1c134349dbfbecaac439e1751da3477;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c4acaf361ddc49586fd29ad05660c7023ebc2d60831a02576a4b80455eaef0248c263b09870996ccf2be53de30f7e2a006d285b7d1699dd5d4ba44f660d51b7cb36af8f634c7be9bfe0c4261ee118adbc9671d1acb756672936d5ed7267b6d7b415;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had524ba22345bee764f726ce347cd397cdb232ca11d2e7213d33ec94b59e1c0d1b4fecf3047e145cac0f12c175582cc4496b1d06417d1c58077e510669798d6d0ad34edfefa77873e07e187c91dacf94f33d4b569b871d2adfed16e1485ea8d39c03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cbbd21b376f715f754530698d6316d37ffe88cd7b789587dbabeb83bdb8ca4955f8768e9d0ab67884549151ff5f945771324e523a55557d06172b3efd1e035cdd0d91e75ddbca1166726324ed56a9027a4b772f33f052b66b1bc631c6ab69431c92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7aad5f53dcec320315f2dc7d164d080c1c0612541b67b528ac96de1237cecee0bd822c6c940a533b9cfa5be0cc2690e43b3f98a6918f53ac2be65699d3a661d7690665f5e3967f69dfb086a80f956e6a19c0eec51a30b3433e923613e9ea6ecd0d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33448c254ef2088b1194929b5aa93aa369fb44578798483c62f1182a21b547f2ff645166a99603b716f2a6350d7604008752d85dc913432d2b3e9be31809460aa0b4d97b0077702f9640172946d24713e278b8d78a8246a829439640ca3b54963267;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h984442a9034667b49bde42405dea6ed4d2694c319cd7aca80c81fdf118fba524704934e00ad31b1eb2d0bc996aee05f1c6c647b4abdf22c3d4b9fe5d1345c69b12c47c761dcce7c95923c5d68a3994ebc54271dcc44a35b3adec7d5cfacea7c2bc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dd300298ea1aac007cd43e564f220e4a3b81abebdd4b4c2f66097fea60097ea813f3d365a0a8d899f162f056083a40156a19d91cbf3a6a290d35768a6ac904231b1bf8c8eba2ac41346565a32dad207125817a57e28354064cc08f250842dd6bbd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d9d61a53e30599c54128ba3c0fae9984e322fc088b1e9ffed55b21dea02eaa9fe0ed4cbc63172b8eb5a0aa0c948803e1d0fa1609403561847118a1e2df55b8f23c85d328b73ae9a4e872211aa10a3951bc8614868604d851793dcfc494b3ec6cb6a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd68828b2530622308d68ab216a08e55577b671331b1541ac2a5397d64e94b803315f3366aea536db37ae43d5735dc0d7dd7280137348f9aec35b822e6bf644a50294d4f6f372c0961be035b34d4ce9c43fd8933d5e48c5d9c244ebc0bbac6e9e05f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he33ddb2ae3a0e9c7a973d7a50e4b53dd78de83ff06ec463eafcebef7107f61c768058e3ead19adb14e3f24d7c0dda45585c5446a1f6e65bfd1ab90a7f245fecf4f7bb3411b2ba966922e185f4e9f4f0df78f907e65583a33c411ced6d6a526f11080;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbce9323bffde5a6bb9ecf60e71f4a6faceb646eff7be2ba229933345dde67d8703cb3a00e395e536ef0ca9bb49c62c1b0fdc5bfca2e0dd7c5ae58f35085d809177a4cc30093fc87a7a80227abeb2f03c2d4a923448bb1f80c271d2bee1815b6e0f9f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a579a81957214cfa7ca245eddcb6188bf540ac9a37c22ad52d9d946bf688e0fb97ebac583f67b590266766dd0eaccc188ebab12904cdc205fefd2de0da91d4c1b9c1a1bd7b841c0d536a34fa4e62942d40ac2d5e908e2d90daf338ec91dca87e841;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7657325e61955a978965d0ca598c9977913fe8914313eafaa6e20dbd99e40ea059ce908de3aa0d8bba70be2b8ec18773091cee6fc4b41a9002c164506ba03b6595f167a611b28f80811d9968dfa80d2179b0ab314bd282dab28a1842e4c1ee3b9505;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1c74b8a1ba23f9324d5bc2579b01db48f08f184c60dc009e9525fd6c902fabc4fd6acd36e2c8400d2e3a5ff5d1ec1ef67e707fc89ec3fe516bc089df3e752318621c8cb4537db9ddb393aefdc574b667fa3159a9f761b94cf71de6234a309c678dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeb2c53946637e3353dd498fb28f07ef9353d1ae43de795fe81b924456c03f71c7330dcef04bd70daaeffe69eb5f4fc314a2165496b4fc6b26d94c5e184e331a658257502eaf01d5a2648af51f4254d83ccf38de9adab42b8fbdf55e2e723aca53b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1c2c02efdb2cad47f199e043ee68c11ac57af718ad974c57f65d40ba4dbb3559930d72fa23ca3b502388f122297de2e84c993d97c2772a33bc9f754b4ac4640bc14d608fe3284edd06ca35bdac589d61d0d74561d89106a5cb171850809c962e6b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h580656423b0b8d35f6946722675973b423c418064c06ff653692f6375c281575bc4ebe75c8539737f78b904865cc571dc163a28687e5bd8da6e19c90bde4f7d986ee60672a737972e03d6c2a07b594dac32c5ad533362c285361e500f57db7299775;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h431132446043581111c04ec7384fc1510b26ab5cc8e8436f395b31c0924089e2e970675c5e2b7ab141b8e3cfd2f5c585e0ef328f230c221f0040b346478162800d17d8c0b6a9206ab3aafc48a4e21128a9f073ac6813bb8be9408c9f0d6af5179f82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf4755de14b13ce825dec82d53084c09640722ae40694f63066ae56a3e1d3ceb2acdd0b3367cf6ed9a5d7b578d44fe306c60f67259ec5ec34f3dd07fa87a4227e7e1d70fd1b2e0e3d474c675b60fc03d542cfdafad383b56c9634dc9638d1d2b0374;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he741252549c15dbd3e01705dad56b759c55e89881713ec333e2635f068ed13c085778d9fe6b6707a344b6683444d01d6b9c3d116b473753c1510897c752b9b91c1a2c32393aa1b7eb90ace21e1b7ef6b6e9ca1f400246ea2c387c593f660d8f9f17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h232df30a285734519044db45d6619fe1401f7064582bc6cc554ac07a547b77d7d7befa5a8381720cdd7458391037c6913e9251d2d5dc5794a59173cb4d35aa3ae72ddfa934749970dcff10ff6f8a6091808b3c599bc2b661d019285c9bdc6c46f294;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e73c29c8dcbee9b6cee429920cff150fa1534c702ab9fdfe9b66067cd2b30b09dfbd27113a20ef2cb6ddfbeb3f1acbdd6ed5acaa06cc920915382df096792d270732412d3e547efda3f9bfec9b0ffe6266b9bfdb839e49d47591b4b25ef3caf14ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b18bf9c31eaea23a5bcf922e4d89812d56a2601540fa0f03b2b928850d5936c1709852c03c1bfa4a508a6e6a817dd7c841d5fe81167a453fbcb4a1cd058e38aa365c8307db498b9383a1f17a4c6d47cd9d945a8e064c80703d03ca97bcba46559c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8228a3bf94242d6c475c545f2d35f239fcf6e91aae6a37ac9bd255adc3453fa7abf30e5fa04b5cd7dd8a600b2e079a437ca132ca8b8221db38a71e3e8a411403d7ea79748c92e952fb52f6b37bf03d72d8ae1082e91e746d823ba686a08581078648;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce430e0e17996fdc4a277793cea848cfa03cd3205ab3dd9fdef9050984d96120b90649f3a4e6c84ac5c6506e9a640ee693784deac9b7e248257b7a2234cbcaaed8a0a0bbba754504412c42dce1f0a381157beb48b0ac2c4f4c83728e7c0a0d82b247;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8990794d07fbc68a07e1097ac37c66495ddec15ef1deed70373c9c8b856ee2490bde5377b8397a21295ed45e86b31f7438b8b61cc320d0d4547b0159c074d4fee38fd1fb9ab305ad0d58a138e448639c2d4fce122e39b78c05ceb1ab271e77cda90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1114a9b0275137b60aa5d14d0a79c57111c1387212cd9b3fbe129ef4ffaa4f1c16558e1446bfa064166f349755f276074b46c865b794d23954e76940371271ead721f96bcbf8ee7596193376827a2874586c4d9a9359add4968e90449bc839f62df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c22fa321fa2e7cd7dc93f4278e27e18e6d08eaa5cc9a09c619b0c4c177e7ed1fd52647f52b493746651c31f26f5adbdd5c2641426164c1b4ecf5a3113c18df43fbeb7aefa8c0eed0600986d15fd2e4a6e4d4faecde89954e37d5ac4cab074f092cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4a1e12c0dcf1e3c87a8e6a20407a243ba99b7cf0d90eecbe1780e5a9361ad578ce4dca8891c255484e4090ad657d72b85f191a14405f8795df89da8e7b17bbb00480f1c1ebe9421b4fe1ba68a5b1846ccdd7e596da68910daa63660ec53d2131556;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd57e00e2e932299a131b04044850f4e4360400534381905454a841602f81ce4325948e24c4dde2316d5e7a0ecf402f9cb4825ea12757ad8ea6eaa641fa094ad4120642501be646c0da9ff444742bcfe3830187448868827a640256c503d2480c17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fed20dbd9b606b4b946e2ed4dae034f2808eb650af47c5bdeed5a24873b1b83077b16c818b5d561de968b543679ae3c8f6e4830eae0950aa1e673a63b5f44cd633e7274719b207c91c6d6909aebadabf406b44a327cd835b44aa59fc4886b08ed10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h349adb6d6bb2e4be833293874a44399bd8227d827d841c737219ce0575262d3e135831c76c7d8a967c8bb2d7b260dcc3b25a4b68754d77b50818cf666e97ae7f0b85663f7a9d98587b684c83bb3de5be97ed42fd099c8a477f407a7ce30762f61d26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h261f3cbddee39979ed2429a072944403cad4828508f37fbe1c5da115157495fd589c0f391894ac56280f70d8c3f03e29019c478b3ac4ea4e243049b4e4dadd32eed6bd4bb8117ec3ca8468c77006828210c0bcd9300878b2d96158f93dd64e43dfd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1375be62e80b98be0584ed9cc00821560d06903ffc4442105d0f721323c62bce47ddc837f99d51fd38783fbd6a8051b37c30e62626335441ad69dc68220b177831227a568ee68e2327fb653567c280b7f8b69292648e1765a333a87557e60fd1d84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6135d6b6936237af97df7650b06a2029af1033d878213ceb43c9ae433b2a346577e82da603c8b94b36e1ed580d9a059da7dabb951b0fcf0a101b0ff2833c54cd883b044869fd49280745d07d95cfbd7629657be05cc0010ac70cc4cd9784ad720a2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h765fd254b9838b8f0e55b5d3a8972f365856944a521bd62897e5cb456fe96c703c80d1bc6e26a06481224fd5ccbb617dbcd111ba8bbe375e8799d8716cc9d7358c6ce0c13a11ecea9551d47ce0b32bbe8e3aabfb0bd924820bf836e062ae6b84c3cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96c50087021764453ced6bacbd32579e59a879faab3b4bbf9cd97d9c5a0cb1c94c5e8de03b5ab0e5a7c091b8c35c9d0027feb2aaa199a84cd6376dbbd8e4d5f818bcf360a38e6d974d7be89795c5aceb065178cb7d76cddd3df6bc20fc2ded29ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71b4d1d9d63e2fe0a8b00570b14796a6ab0896c6162bddb67c1af6c56bb9b54471565f8ffa6678d68674258265a16f527e09e05c22d61c63a96308870fdc2923b73293c5b94d0cb9434667f9a0a4eda42713eaff1409c3648842ac680e9614130101;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84a1e2ff715b97ffa46c0d5a6c6dd689abdb5aa69282d24db25e9e8a6c15583ebca9d5f7e126d4aa451a5c27860db4b6e66b09f9edb5e0fdf1261116b67b61f65413a0b9be99c420338c3784c237afcd18f7e40129998907144932b22983d3fa8b17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c0348107278af5ec04332e361a30fa0da99d356780e5ab0c8974b4a7dbf044eeca7ba61d0a2b618df62a6f81867355cb0fd78b27c95d09567e7b57c933c3c8018bd74dae1c9cb20630ba881bcd24be36e2b93989e7fef1a2fb6c47f234a8cb5622b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20f172b57ade2d06322854a67d48ef7077b33d3c90f5f8efca6a5816e21f4cacc37ef436a6bc3f86e52feb01247796213c6c15e3a5846664574b0000f292d8508881341d0ce47e7407e8e0589f5ecb1ed25bb5ea39b2b93b4b5d029dfa6068eb8908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf274c01b5c7e2fec4327aa99708f06ef681d6973df0be551997ea1a8a6fa9d190a198a69db875bcc29c3d777745c43b5bf4932615530387e29322af3c7d3e4590aa4176bf9d0d3cc783cbd92aefed40e08a1df3fa5cb1aabc88794871e3015d6811;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdc10f8934f530545ac221fe956e694eedbe03e0d4aef7d588b611b04118e9e6aa9414f5e90eaae205b47df0826feacf9e5064388ef0b1ddb099b28bed21c4ecb9202471c4ebc78a8b4b80677c53cdbeebc67165530cfb2cbbe10dec11e2c4c2c383;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h717e3c5714030723a3782fed709b992e68efe6a9e7c10376abf99c73c991614f9a77218e7a4bcacb503bf45481c0a8568200147c800b7d58959ddf49fbdf573f566abe279f206b9c3dc1088859de5a0471ce7a8868042d79dc1e80eb8b813e14878d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27e21febf9a517c6d213d6ec9c59706a00aa720dabf7650d2f4277c336fc27bf66392530a7a37b5d69673acd11a0ec3e1507ce2e4b1d984a019ca11e2bc30f0abe955eb6e79ac085dacc29422f2bb3698a280f6da87da9c0ad315b18a9ccc9bb875a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c6f4f329f9957308e344808e7646f27fa4615c3ed63ba5fc2704acb8465d5c31b1a3eedfe1b2fef14508705718ef1d196737f90d92533fad2629fcf13772036bc4e0dc13d28422bdbec1bebe04170cabc81ac298080f0eb9830d59381434b35e9fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ec979bc6b58fd1db4ce13e1d748036a214813a1524dec593c53876febaecd9297629c617e8ee91316d14c73734925cc674e67f587ce31122931574043c0aae6627c1e64a228035ce5b85104c029d6ae4f7830cd75d7af90c496ae30f23e0dc4041f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd87a2e3f751e1e7adadd6edc96e8f19f9bc5120783eb00dbbb31f86995d2d8e20bd36d733ad4bc3148131fb3e6db0edc7b9a48a225c844c57c4b8c120880676f32e2b8cd459272226eca3e3615169a372c2a4087e36744efc51e8c0003b7d1e2956;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf750c6525ceebb877007a64bce29407b940bedfe2a92c45acefc04d7ec222e51396d78f5cbc9c6f28d40ea449a0146e307b58652b98ce7effee85970a49e8e9dfead75bae4c498c9a4121f02dc7231dd027a25150971bb37bd3454945ef1af22c0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf479e27fa059270e3bedcad02ab44893564dc27c3641e8321140f1b59bf9f9ea303878b7ff3290d752b48ac31a36bd3586ee64b0173be582ba80b147a0e86e8fa7edaab125226d0b4dbbc9d8fbbec60a96d4c9165d8d208d00d8c0cce13a89d8489b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4fb9d1c7dc32eb07e588c4f3d8beeac82dbcb2479dc8369703329a5b9cf96e5f436e7912c71d0609f255fd00d54f5b0f96401927ce7d350ebc5ea25d3e9d7b754ef0e777be55e6fde875040a3b50ed20b36769b6d80d2a3b5288dfa7dbf35e975f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53f29ef899b3e0cfdcce2b44336b9e6ecbfce4ffee23564b9a76e3c70b4d6255ac1b3cad71823fba85074bb7080928094ee5987d994e58d92baeb89a24ffee1d6ff275f6f07f9cb0a2f9e7f3dc464788e4ddab3cdaeb9cb83b5ddf2ac882f1e5919;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a91685479cb36725a1a490ce6437fd17f94c06edd2849234be51583b738fc9ddaab34a35fa36d1b1fbfdcd9a302323a5043ef46a02b9ac3f3874481597e41031ae3e77118da05969324f166e68b176523c0bd4c45f473a904933029c966a7725feb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf54d4c7693437584d286769b70fd8e9de8c9780170d7ee0a0e29303abb2f53e75f6577667fa250a2aeaeac8fd0da85bbab16becac4fa68d52ede07c4fa13715cf581bd635febb6830645eb6b230c24e57fea1ad6f65cd6fc96eed7f40c531130c0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h481aa85616da41f041264f63e6e16a46125a95159900c8a26b5bcaadd8637fcf67f65a9d44e7cea42a7443145d5735fc80cbe8f20864c1d1b999bfb5186d0091fd597d9f0407b0d2c58c7e533e46e0098e4abf98a13c15d39beea34b5e64767a2299;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33709ee6c04ffeb157b2a381cb0dc0ad3ee9fe16ef0cbfa250f48c6d3978ea678cc16da05082cad285921f005a85559ab72abb6c984f2cd3740c5beb346abbc0721204f9558fc8546dd2db3ac6a986e1072811f80f847e69b0f09ec69a251da9a2d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9be76fe3b8ec87b18bda48f431afef612b4865d7b6deac6832ea08c2503d052c80afbd6267761c8d815058981185ba9a92187f99a8636ff46371cdcc23393b87fe8d745e8477163e9a955d142bb7e0ab1111d6c0202961f3ecc8b6c706e85953dac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ae909f4047d5905932ab53de8feb558b315ca702878df0b982f7bceb325cb0396c730225b7956ac8f6022b6b9f3df03e0e927b0c7825cdb0ee899172f1b466c6bc9c5b004e6c24e9cd08c4a96c0529bbf58b3548fa51231b21bcf0ec01d1c1c736;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9bd2f0b8bfa1005da445695c1e7df7bf6a0966a238d484bc2a8880ec1d9679dfeca50a5c17b2b76185f0c6111a20f70f1ef20b5daaa93865843e00e89ee79233a652167e4cb36c07748ff29754a028a8861d86251eee9a7f245aedc1181c4e2ea12;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb258c064c22bdafb70669f7e4bb9dcf35e8c26b781d97265ef1378c5ca12b2d054e08bdb5b509b544e293f294064037716f266c94b0ed6568af57ba8ddad948fb661f22eee04ec616d5516dcefe61915bc93c4b148cbbbcda08cef9a0e18b98cbf9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7877d13ae2be1a1d83b542557712193929d31b895b460fa826aa0eb327895c3072d8304ff57e5a08dd4b9145547baafcc3560d8bb88961aebc4c78539475d44eaf2f9a9100c0b7ed2c4290c69ff9a434295b4369b9b914448374de9895211a1d30f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62492bd72d1388078d8ce5836ded2c77112b2b039d79c51dec343e302dad9fa3e537d2857f977a66e6cc47b1dbeb4b398a8d652b2c09787851aa2e1e5e1e9a819cc0402c9c95f5bb75907b654c37a71e7f5c28e5933338b8f8b122f9aa22e196c75c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc65d1793892c0d7bc702c5f237d1803934c044ff8c7452fcdf617eea97ff6f4ca591072376fa8256a913e37ef3a9e337f16b48a448ba57bbe50b6524a493915b55e0bc29eb18a71e420dcc6b9c1f0b07cd2450e272eff0f96419d65335e16edfdfb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he234f21a0bfcc7f23605d47c1aad29cdab89bbbe0d85856b044fd30824fc1f239ee534c4801f0b247bfdd2fd5163725d63062decb3062f20e095ecc986ee7ac65da0eacd81d5383448315466cea3f1f5549c7edf90f2181591350fdaf744133f79b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h609c10cb522296b25a939db97144a6466d438e65ee6cdca3042c92f6abd52702c0e107acffde8d30aa5ceed80c4f40eea0269d7cca97d868c10032fce90b637819e64427ae60901ded8d4acda32746f6a6adc4f08f91fcfeb8f124b4b109475aa4b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca7b0b82f41d4a2294d1a41795af1eda4a52703bf4c4aad1e37001efe49648c4f354d6f509aae2563e4f1115087df027b4ab99164e8d972decf13e99fe5b32c09dbd822df6505e94d7054a9de0977dff50eef2fb364a59bb2f9c474d90a6fbcf1646;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94a72c82d2dac6906beaa06475808a76cd9783a72ae5b1c0b4942ca9e4b56439ed935c9b341c358c40de5434db5eddabfc21733d211ecdd6aaa2b2ffd939a5540e891f49c1b5f9a1baa3db42c04e95cf05ddd37fb7b4164326242f4b9ec3ff09d12c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b5918d0d84a0a84f00a5dc4bcd34c4b05cf651db7f6ed412920dae02869ce255d2366f09a1ce5a3d790913aa28d10d578a5ba338e11bbc430784f3056135f3ef60cc08141b165190c85e0a559bfa12c8590b4198beccc33986eaf60d331b0231ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbf676dfdf0575b013cebaec2f861300227aa876fcb2e95ccc6f659454c6b36774f8f10b16e031c9649d85df4432ce4da174a48dbc63bf76793a4b3712f62cf0ed9d3320b38f2ba28505b934b033caa7392b5f9ae4edb02fbafb0910a7bd645cc800;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f58666ff53779554b44aaa7ea47aa10d10b5f3c41cdd58f1ef989f2f68f6c30c3aa7a3b6c0de10ab7f64ce93996165dc3058903d0f2af4850daf61386c322e771cbf79d94c930769a6b79683e259713e12f8fd7ef91b57544b116e58d9a4d810e71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16a029cdbbe4376cd49e3d29d118d52f0493ffa1b5500d1d7c5107b134a2b6ee71e0be850c104301c3f615f99d18d10e0826e4a21b3198c94e818705876eba03b833ff53786e0d4ccd0861f4134e33f29a4d77022a571d7262b08de1bddbb6cd56c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3bb8e9d104a239050b02dd4dc079d9402bad6fac0558c3c9889531d5b3d793e91c86afd6d580a8841540430429ba70e367ed24678f8d2a806320dcfe9cc10145bd20e1591c92460d1d84bfe56fbcb37aea8df80fe8226ad50cfece6e278807b649c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8764f307a5a9a6bd610f6695747419438cb2d01222afd87208588c554f7a95be150a1dc1947c0f1f2df3f313e2b1ead36705a39f442bdf0f49a8cd9277e52dfd878d17b3bc3c010cc099e53bfbe3a099cf58deebe834d7106de345bda44b951cc1d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99d6853bfa84c3b1fe2ad03a5e7cea30a23fbb138924236fcea92dcbef03aa8db5b4c1877b21dc1273919a1078ef6c467dd28961b448b4b8fad99322eb115e0894e437a8ad4dfc92e4f27cf340f35884f3b117942e223df86b563209a680673487e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3c3e7a404a2b1af8f3060a1fbf09abe0bbc2e67ce7b8a3bf500c637f1fa201443040559b6947a63ab5971f5ad27ea651041d5a86f0f96f9f240a456e6654181822f2a052163151bc3aa0d2758068dfc4083c92312c2856dc9ede238d49088238659;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4405b1f3f5943623a0acfd599fc8fd3a8274970544ea4f17182f4dfff9ecfd6051727e4612b0073490d4bbdb1fd082d6fac1215d3f943ae95527fe71f9b4a1895f3970ca574886f7151176ef1800fc91f1cdeae1b785149dc114dca974530247e347;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafe1a102460306e7d209cdc06e0adab49676be7e203632720adbd292addc72079b4973ff5d6db4356fb4a7d766426322b6368f883009dc968d8a77b17f919036f9a46a1917923451cc91575e4278c4f4c0cfab742b58d8c5204865da9cfc36e9c6f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1294232cb1f04c9cfb160295644a64111a1ff6495371504b54ca9a5690427a24a7d90bbe04c97347a227ab9d1d2c5508796413d4adc05174565a9da613b66ddbd309571e3f2f0812eb296c6e6b7bd62600b4f9ce50ebd16f81c2f0267f922bd174d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd406bf5be785dae8bfab28e10b4539fb89ae2a611ced49b59d40a1287d87e8638d439778e3b6141dd34569aa5f688da0b353dc3b48727f067adf8397432886e1949042d4302408753b83af1c8812997a84d6b90f502ecac8c88e31623f9f8dcd102;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42f10a16b53745f5444ad6ddf7c79fd80e60f9f1cada986c4b47498ae42eb230cc60c9f0c693848cdec42af7a4875009031a92df852806c6d9e2d577a2e9888c045c88860c1af203632b15972a830d00dec688b02050274027df43db5fa752345168;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38ba66f0abdc60767d7402ba59b3effd4d1110066336e0ef90c990863876569fea21a17f7f1f00411d6722903981f528a1911f009b7c4dc7c35b19d46f97e3cf8a54a9c00af3ae0c6598d7461e08b23b4617442894e912df7f704e2e7eef9e34d540;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h144a1bfa0bc2cbd6c834447033f43a1965e3ce4d7233a07d49112928e9847ab2a8aa204992972bd61a0a994378b41ed73a6d0b3ce7d74ceb0f5ab7c6bb12a97a1dde6348f078de1df1cbe2cf59e03f7fd992e9f3a153593843309c0f79dcc56fc1e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fa741c5afe915e1ef0827b8c97fc4ff648745e4e5bb2d2b95ebc2610cc802d3f2a3d8189f490e0e46319a6e1f62015224ec27762a34ff048e81130eddf0692ccf39862d0b7f42353c1b81e4a656a3a85b2dc1dbc431547cfd00a8aee21753e416bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bb74edc2b4cc24000e96da0f731a4f45efbfa668281d74739b08e636630f830c03e3cb499a7d7c94c66c8ca28ce588ab093230eaf81d324d06f942a5f7d77c2cf4f89ab9c755a96af636f0cbd46dfae876ed226bc4cf5314762032362c165921e52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had8a62a55f1d91834a500a93b6426c30187c57b3166c926447f2227adced95b3e27a0b69f2512b25167eb7bcff9756f83bc052043eb0de6fd3b4b5c487f42041cbe8f4aed9d11a9a14680ba3bf78397c1cc4d9b7246a9dd0c182d58160b2a88dcd79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93834b47d933b37f8a2d03a5ef6ac5276060fd73a66f07126a4c907c256aee1fae6d4d23f428d25c61d9b751502c77e8d64021f291ed77c78c6ea77b2b17f672021cfaa5a664f72e6479ad97f2e61126eb64ee70e6023f8f3392bf06b91dfa472773;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc777800860b37c0f866b8431c0f19f40843aa1bf91243f569c7b1909f107e946c84476f7be81834e74b25ea71c9e628a95cd1cf9f46b65ad3e2bff0d3dcdff3c2ddb20d059a9509167f7e72c23eeef323f3fc33fbbb44b29f2156aaff4bc14f6ec18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h110e4f9cd9a147b25d6abab00866739b38443b6d256d2f73dce2989e72f2fbfb2dab996e4dc006f9695e585ed764fe58a0ef3bf2b5646110487bbba4890c1641cc7ef5373494d00c712a7e6f3290e082c24339228b3abd0d73b16e0f6f2d472f904d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h139b1b8df60014b8bea81b00b3bfa30efcb97198d5f9ae371eced74d91805677ad5a2047c061f1b8274310509c64e23d704a0ab5dfc4a2f88df6c97c06c36d76df450373b8aebeb7464e576898a01bbe5da6cfa2e0801d292f73f494df18feff1073;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ed89668276e862dc9f312f000dde29bde15eec49dff6aa59912f1f483622ec525e50acc153e29fc42ac5a1ff8ff84496821d2d874284107b9464802a7cfd78da6f39be1c25fea62dbdef32b380e897eb0627240fe1cfdbbdc4dcfd7552eb8a2a1af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a17547c6bd7b2531dca4593b80a3f723c0c574fbf1105dca4992775410c23ddc9d54520f7521443134b65e48a7bf2249aa4c2ddf95b3f3ada9475ef69255add4fc633a9dac6d3b3d777d44dc5f9412531eeb03e4faa0556ba208d1bc0399a012af1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde531666ecc0fa03bde8f32985d213b53374e39ac0162fb3d9c50caaaa98df4b136e0fbafd569291d698a4937c9b4fc21ea9f170f529c285a8ff2a94ab04b0255de2dfd90bd11328d18ce9c86f6aaced46f36bc48b7496c563e32f25fc2c77183dbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19d246976d7072f90355cd30724e3441acc5def15dd9ee02f0284467c9ccc69c5f5ed0a854853b0c2e3b284765d73e9a248a1e07eed8e1cd697bf6f3b18529b08fff5f1a3b250f9157eb4989cd8b42c4d6c2d595e2338d234e66e893fe420b27fc43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86fa3c9108b0baf3f34d9d80fa7db56f35b82f5c676c82833dd8be17989babffaf91f72d691511a238ec664554b05ec91f7a5d27b01e173d2bc254e122e8d5e98a26994c8dff99c344f12cae1c69f4d0de13a80a66aa286bd7bcf2c835b6bbfa6445;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36814c98d26e845f6d171480d888ed7e74d701ed47d4b3012eea90a0f20ff27dd202343bc11fb5ede04bf925c431c9bc2e8f8a5d26da825158cbf52f60ce1d180e8650a1edfe28fb698d7a1633e1a52239bfc698f03a3459f7db6218bd89d5a47195;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ee839457222edd2bf71c629131d823c59e19fa5a7a9ee3e996953151c3339fde08e9505c2106b4eb586cdfd3eea6e13757500adc303d225a3bf08cc12f0d55532084a45183b4fd393c4cd50431328665c13553c12816668807722b28170ed8940e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d942d02ed6f2287813538f964e6183ee9dba099b29fe3871c7b743527ae74a256e9dcde92252763842468924df14f914e6f20b661235f71cd57ad75049f53d5ce605653ca86106773bc1bbf2b7656bb55e340148661f97199d49595bad8c2955a36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e472c6e09454d616a245bc6647694b697b511095e0b5ebf5ac52d374e3fad04b45ff94243da6e5877a3b54844e6a5f6248d703772c2cd2bed738589ce2fa1d87d1be476cd199f458a62e0edc9f024030980a8fb16f5bb784929d745d23183a3420;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5c7e59b634e2f3301b47fb77632b9eff6e6c5e30d6949aa8c5b450532ea02d9138e075d74facd585c7c02781e015db306bcaa9a3bba711170f6a3f78a0d4bf8aa3e982511bb31997b891436be924920a64c4910ac32a8ca4834f313051d61416dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3722159d8d0a90cfc23e03458f9f270f6ed1e01c29074eb11277104fceeca7102eb520412587ae99156cb5e42a6977be2c49b802062b723a20b0f44e438ea6662c3b06d1606a4412bba7823ef44f478e37c7b00837c4da4eeff5195d9fa5562b9f02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46f145614d9254ee355903dc79a16199ff93a28e422b32e5e8840d73f0de13e04888d00f494e5eb010603675b29405a943bf22707bb2a55745a2f31d5e9f6b602db23a9cac97e415bda29ed8e60a3019840a9aff2e303bf53ec65d1519ce3dc7cb5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a1f2ff4b26ffb1680466f8ae5ad1e1c5fc0037f61612893a7dde9409631bd346f87ada1d85b435511c5e22a9aa73cebefedbe9886c65d592028527a146c00c5d67bd84a1874f3897ef6cd78c26b4c84fb426cfd899057624bfcb611e94bdb29f696;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4655ef5244786d06b7601f83dc09036d584aa5d19b66065f93f02a0ceee4bfea6f295fa5716194635998d81182b0df7fa805b6ed668e97bcf8551dd5f6b05e483fd4454ee1f4499f933e5596dd4d7e1d8045af6fc3a6ec277bc6d67cf5c1bf0db1c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8e145fc8ed7b84fed5f620a3a73e60f76f602743fabd3d521e0cfa33a0c4cb0c6295567649b89f917c35ad672b9db7b69a0f1f5d47c3d01a8408a9fdcbda5793ad4f40105afdada6f172458c89377dee88a9a2aa220e0150db68f5f2e0777c67ed9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4eecd1c63cc13b119950ff433521db1084b6850a111359a04d54dbd8cc33284269360eded55a8decda475406994a8b1423ecd66277beba7f90bbdd1d44234522781beb4eca20efb493c0db71f9ece7fb0aec14ece9bfe4a73c5707ec2c35a4a7b2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bbe606292e62742f3135ec2fc4ae6807fcf1b35eda79668480925bd4a8b5d4daabab8e848004108786a2b04aec3d14d0d9ebe5a77fa22962512de4b5b74ebfc02a1018d03f6caefa1ae75c0a9c9af2e0bc4a8cb0ebabd4fa0c3a79735760fbab2a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf13fde5c14a03b7bb0120ad040b6e576a3db3bc56bbf8736e7ea93f07556d1af4a28d20e2312ab7e28833f4988c928263e40b7c5a6cf1038f8ccc5a64bba5147c97bf6afb32fb4c82a21de08ed0ce30dd342d10e48519348964e37a98cca6e63335;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ee6c239d4efda196a084eadf637a93d85b6b4ea48be79f45a3296c232dc5193caa795566fb79a6494c0534a97d02384e5eb949b26318cf582749add6b8220f9d03d1c9422e8e91920915e95416008695b570bbbdd58688c2fadfa0833b95cc39d2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf025c2914259815e7839b8cb546570ac55a804193542d4cde4de2595d4f8698d1a6ac2b88ccdc3fed0bbde5637b867918802d789a57dc648aadc4e2370e3a4f4fce755ec8011b0cd2423eaa64bea704aebc380370dc51da48906bddd4c69df9bec8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1cf0fdc8d6287f1847e241051d2a3ed83f33c3ae28351a8a0d26066ffd3daa369346df5244a880ab8dfb3aca1d6c423b647a1d339782310834d515e8bef8e83a54662a2e63b15773f5eb5a6a9197b4dc16872d9718b4c48a77029c388d1f127a97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0a2bba8fbb49705b5c5cd2c3ae9a5e4f4d65678571f36e2d38adeeaa36a17a2b898adeb5043a18f92adbb50b6d49e498ffca9d4802554cda83238cd6cf6b9bd418e98a5994ebbe9c49317c4d8337745548a1be86740715c6c81ae2312422b8af752;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21b468eeddccdfedb21634418a323eb58d8951feaf42c349283fdc2ebef2f28300a8200c64cd5781f815343b86b6f63521a4db3bf3a2dbadc7232db1e351300976a5bc789cb87af39a555d153deb5a60116995720a67cca033b6199f4ca04b01984c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7727eae23b79690ef96060ad1bbc3e0eb564a3e9bf9378f44918913f752cb2e398e0f1d7c46f78fa995cbb377a7b7fc297b3157ea0f5071d97576a8254583f57e70956fade9f7251661bf6fea6985a4b17a428eb53311a26bc8d1efb3fa459741d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b0b9ac09010495dc6fbe13e35150bb2f14314127aad089c7477649279aa109b75b4fb062071e83f3318e60655a2c74a43764d2d27366d319f0c72eebc3bfc3f52c2f5913eec83c3b211bf2eb11c34da4f20d9c56c272894a59bda4b69e274756f60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c7ebc0161556699207ca5e1faddcaabfcd17fc66903e3e0d7a9f7a60559bb7013acf0aea2d4f795486cd1840639e8dd140ab33b1cbd11ae16dd4555d23f6cc785cb41ef96f6398af87f61ada237c767817695f91822abeae7dce0ca9550764eb495;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbf249ad833b37fb0308c25e11d00d23fa53bbc22871ee2aaa7bf2cc778030567d4bc5c25b19d5d4f4e1a37043c16d3d78fe1997f98dc61e5bcde5cc1309dbc76b0ca83e06a3ebdbc6ae04c413388220e66b4172912b1c46c523b9071e86cc338d4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cfac17c4fc2bec1e909b5ccfead4163f67bb60ac3a36424999abbd5b296be7f21dac251da4a48852aca87ca3a356607c0b12710ee5c7b862bc973f6f6da967f78c61a5f0a1e58f8023d054e365d6eb9ea49aff2f0625fdb10d8717dfb6a8ae452e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd5034cf9c7097efb2524fa23ad69e2f2a1bf4700eef3788e7379091d0c1a2a31d3394902dfc5079193709cdcfd8b4d70392530606478e9fb16c12dd7c743d579d354629f0d1d1dd2e4b8080e14324db9db2d563005bf4879abd968c7939a20ac181;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haca2b3254c696484aac879a1ef708d432c048a19fc62e770696c6685a0bd7c3e34034fbd8fd7fb8bcd3a4dce3c53a28070e4d6240be60050be018a581f1d6ab2ae4b50b03db18130c823d191ac5c0ea74965910e7954dc4c4fecae1b67b3748e8fae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h808e94fe18b1de7922384d688a534b9bd9c9c4b3f7e562a2c3a71c9687c73f0a2bd0498d92a97a73155d0749ce234cd9668e4aa168ebcf0e4826783b33035db3d5a7be4369bbca2f1e2e05cc667818e370e981055b865d8623142cc52a13e7bb1120;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e0d60b657eb9131cf61fd9cd1c105c6faf20584f4ab0065f29761995ff5d47a2c1fc327d7609fbbde59b851dd51c0bd739b68e64db8d3ab16623ac21f47a6762036c90eb4e87eec6e3d05f341db8efe271cd66fb87fd686c8961c4998047ab96267;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4203dafc58a8ef554221b4d0ef5a15dcc6de003545af44baac87c1251639190917d38571c97afb1672860a287d3eb5fc06b707d604e496df048f9c0210faabc83219aee6bfbde98771f71b10f55c4261d9a89b5317455d1721df9f85298ee9c66e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6e7ec8543c1e9baedb16172c3f4d929fcb6cbf408f1135c9027c76f93c9f16748a5571133afa3b856f37cfea45377ab3c7877ae5d204dd89943293e516093d00681babe0478faa71b9dc7027dc41ee86ba1b568042ce570a85715c3b3b8212c8e6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde1f2828ffb758cf1e1a811373381384d672ec231a97370cebdda28cfadd9c55584f8cf8bc750fb9c30993bd8b1cbdfad29b1dbdef0def0ce01d695319d06d8fdb3886d8f471c5586a43122c7e73235c317f159ee5c155a99dbc7b57025330053271;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e6f40b79c47e2138dd54eb2e1910caa5bf56e956bd2b3efd9a1a8dbe5af160c86e6fb2b1790c5f6f5d7af951e9149411d890902b244925cdad1f72daac6c5b46bbb4f575b61494694a81a5ce8034806a4009c928315e2b23de97c0c5efbec300d7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf43d309f7d7833a1c8316570d239518f7eba5bb3e415871d858fef8f0877d430e32cb7fa57fe4080ec9abe83ae42b79f217448265b68eca7262c56931973f6d9c102e13cf198e7afd5d84155cafb69dd362c4d2215bc2da45f7448197200514f208;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc451b09c52cca0aa7fde6c6b997740bcd202f2e612fd0ace9487f1da8a6d07f4ca8370af4475df16c85a27d079536b69ab729c82d21a4358ac30fe5be8cbe120c4d91a1ee622677c71bdd9874e335899073395745eadf7d8509276718a2443e6b99f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bcdefda54a0fb9d042ca7a8f0cccc82f637b35470f533894ed37cf8446e4b4570d754afa294c3f663fe06b6cfb35d13890104229d36ae05b6bccb1a6df290e89d49594e01f9a7302fd8cd3e08bff95da56ea4c7ed18f879ef3e8d63025d8de8de74;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb89bafdd308db4b7ea868d9dbe71ae543620a106e983f842a8bdd49e2f9198585019588df1d8d78f24c8c210171c6c6b515628ddc2ec0e2697ddc422500db34282a0e6e06f4f83daee8f37512aef793f80aa0b322cb0b6be1de927454180d99c3daf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha51d125eb8d9a06afb1278b1bdd97a65f3c4ba2c6f331ce66e440568a4039b76cfa89ead392d6c84acfc06188d58288ce553ef88807056124f071c0119bbc34479da3ad78c1d4f4254abe666f9ae673c2f718634fb2bbecb356e291ca2e452abdee3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17841d841b5d50157eee366b3112c9e6f5dc1e1ce0e534802a3a1cfdccb9d67764f4f5f4e1e3335d2e84efeb8e23af0aa7cea093d84d4af6ce0154de7cec31205e97255a644bc1e49c7756b5f62caada23b019555dcb6cd72f771d85cc49408ed95b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa6bd13ef2b0a9369864cfaf3c4529871a5c8c635dade648237b5f4f76ada396358eb259561831794ad0d76abf2b41ff712291746dd31070ec8631d668186640d43de146135a49a923f807cfc8ca718140687ba7337f56764380ffc4d2a8beef1129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44253b04bcaefd86b280ef8bc8e9d4f99db52736fdb10fac525d68e80b82a5f26ac123e10a56b9be63234f5bc37f335c67aaf77dadee72dc680c7427b12457d9e99c61d2d8cde076c3133c535801c98235d840e68b457f515d1ee5ed8667a6206094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h584042866c60012a18ccc4cc617f6cb1d944e326c6d804c6a46502b907e3c90c5ca0451196fa16870b01b397eba98b2b38c136ff30dbdda366a8abfd07d0315012bffa318427aeae7661ca09dc25676fa20be0e4f1a57b8eb00baf825da1e7674cb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e9fa15de6a3470f1970bc1544c9710f69bd7c8ffc184d7ee907774c090c143d1863a914a065fb22620decd4d6421abd475bf890e4996c0a63ae54f2ce2abc71509ee5dfe98a9e3648cdd3d3915d31957678cbe329ec3bc67f584188c979f813a361;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56da349e4f3bbcfb5a489efe31c00b086cfee9ac07c1e32f425384bb1c24934b3daea8b0c0df63103639c407ba6306626aa0ab562a36c5d5255528239f26f9baa4b0a718420d13fae27e6f2e4ff0f440633b6ae67199ff4837a90a91a97e65e257a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c89313e1e88da6100ae323ee4c9ad871d6d3cd68cab8065286227f415b2dbac2004cfc7c16d2796719e69576a81e8fe83997fa21fc1cd70b8a18126af7f80eb7699fbddf83b8c587e1891dc2c4b2e90a6ae5bbaa88aa5d89b60afb5f48447f2bee9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbac927947ffe224770c132cec3a87118101a05184753b63257316db4b01726a494974a29b9a0b4614a917b404778940d6edda4de8698639f4f2f61fd2a43a83653caaa956e1284df1d76fab8139084af3975b8d6d58886e42f015737f2dfd4957e57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf893cf1096be44bc3f1a193d18bc499633c2b5b964158c6a4362369c12a5705bea4eb1fd29a8413d4cbd401c108af744e6406b91bb15d9a6faccd6e851511ebde72e1e699f93af36b949211e2978ff5ca1147b0689fd1be1e667824dac5f7b50d73a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h648341422002dce3475aa9a9c2ad225c896e35279881e608c8083784d773febe180e882f6cf0c21d9cc81f54c80c5c392577e03d24a332f7a093abf7a3025763143bf2ebe69c9b28443c8270679be97ec1832a3e5497293f3923944ab990a1d1f21e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3527d4c2fee0a20db2d290ea1f80c248f5d7b8bebd62b2d903b150a82f9e3efce33c7d2d21a33b7f1dfb82ec156ec114ee4ddb25f274ba39276f02ae1cb989c70ec660376b9b80f086a94fed5b5946ffed41df3b46d2f3b702f9ec080de3551d1575;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ad407d327d0c0222b918946592203b6014931ebbd1f813b628e52d46916808db7b60b3ba95a2137805b8bd499fc56ebff7bf7b8412ac8947c683ef4417cba954adfd108b1631352a849bebfd29e152516003db519df423d1ddc10dd130eb57b25a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74c7a1deea5f5620f3fdb4165ce34679a661d24da3075169eba12a06fb326c1acdb9e07e218f7287d2556581527ccd1b8417fab10ea04ce0ed4d93a3968f30937e566cef9daa5c755d9b548e0dedaf008a183f92f64be4daeb6ba5d75eff78aeccdc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5e89084e1e347efe4980440420f076a477ca324b6373f2ba2237e56938605bc741f602250f7b126e6a2a5152578233d0b24656fe62fd8410a45152ebe38701cdecf5800709a41b136aaf7df5bf7b0a6f98ea0bb557f688a16d8df6722e7bd6b36f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f0e0ac969a586c14c6fa78302b0da510e00acacc4731e6023c2e84d19d4306a08f9517e6d7a6528a711bd0b18ac9f95a20178d3cd19ff8f2100200006df1f03369a8f93b5087cc174c37559e93f8a7cc40a106ce92f88579f6ed7a21f8eeafb791a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11e52448d178debcfc9e3ca546e7e0a4fc25ec9aef8d9fd96d5ab53360c0b46891ec3d573d366e0d6739c65b7f967f7eca71ca153d5309c8cab4b743c9023eb156388f4a1e7a17bc6da2fbedd33795b91c3bbd77a3ced40c75fcc7c019ec518eb8ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcad5b18cfa2c362ce2c5155577db295f6eb02812fe6204448fdb44d5598fc1b742a435fd7205f3e97186afb97622dd60d1add42f33da5dcff2f4f92b787cb9d1ce522d614216f6d891ff5e74f6f7d25d6f1de18a005c92961d93e3304348bf3600b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44f3a2583d65c822a2a0c6b9569c10dc3e0b3bc4185fad784310714d9cf6d03beb15c97ed85c51502e616292fae6046eeabf141a1022152cf37eee76ab819b311c46652e8457c4c01ed639009e757fac453f9697831c17dd480819c9ad020bfe96c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h319a921b9617d8587e0a75213f62efbf0fed9eb49a1248241033e15046faaea3754e30c923f210c80ab4ac30b3d7513348d65d099078b0a5c3ec866d4352c3f899aca52eced3c29677c8647859e4ff1ad19c5b7baf9ed3445cb3b40df836a07cb1f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf072133a84a6f4d47e7c6ff9ce64dbf3c1f47237fb8218b8a894209825c7997f9e5ee196b33ec3ca431859336a0259f30cfcb9311abb821bf6455fa3fd7184076ce9b858b3b9305afa31f1b983aa96a49ad40d50343daef6f5198590250c07462102;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb44ee6db47071c2199b1ca4dcb1102713754a129beed29d9a67436b6aadcf042657890fa6a5a0fcff6e22229f07c17d12f25bd12c14e65568b2cf8abb1d6b1a67ddb063e9dfce7c00c26d9ab7829112d652ff36580c904b1085f3f19f62910dea89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5141cb320f2092c4e5b7cce0f8157e29e5ab80d776c8cc57a7f3844134147b9cd7ccac8c773edb8965c02fb059e254b697240386b94e5dc712780ade8b4854c0035bf9eedbb698e4f6158c0b00ba81eef407143ee1c83250da7e50cd4803c21933cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a3c5c83566e60b8f65cced5ef9ffcc5ff57375b5b775a2f0ff72168315a3a61d1facbb90cd84ac42f4367fb448648b3c2d49d6b26db7850f4f1da8ab5a9e33819856f6ccab9f7dbdf4806a80888bfb7193b744d3835bcf9f7e0469ec3b5495f3a0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h662158ee8e45b58d973709612b4549d43b4f74b2a454679567c21a4837437ce4ec0d9da5152634e1561c69146e67bea1f034436490b62fc81f3cbc4a0f8b4d7fab876b2184b1916d5130403b3c6b0fa99c9bfb4e072ffba39c6b7932733141815b4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16291f86230677a6004a5d832a3c449ef5fd9e83c4fcb576b6ad7054e86332d6b9aebfd5bfc7b2179e4188e9c16efcaed41c730140dedc05a48cf923019860e6449b8a12652f839c39a390077e1dd886195420a0a4a6c919089ef2a88ad1558a8923;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc58c85fe0a807720964ba1163f0979ff51cb1f705c10d038f72e36619b3ebb8a24660278cbb433eab11ff197d2514cd2c27ff7e29a89c097998c9f69481c051aeda8a4d16f4b86e44d41e15bfebb6c4c0715ab5bc3b266591414d092a39f2a230096;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf21e7eac255e6c5d09d516003f6039a3fb27d712df315f717ae279c5b66a37cd0dcd37976bc62d2b99f6f9ec49bb7d9255af312cdb64563b5d4d0d519acecff322d21ded0c5e94e0888278ac23df860cb3867c29db3206939ab1f0b8299e063d01f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h668824509c07357cee625b64149d3c77cfb0dfc035063a420985e3333e04b71a04e2fcb42a13efdfa1711e53e66e21071e1966a092a6218e07b267cf4ef961d4e1a77f149cdce29c0086dc9b2709e388ac3cdc1c1968cc9552b2445d69b990d7d241;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4063f254003e07d1d0b5d0ce24a58343f8909251a1692d2f5d0ed434ad79a3eb504b7e0a8953a4e46e9f800215e8c8f5d5f9d58b9b54ae7f03271875d9900b154f837504f3150cee4ccad8b49499c0c13150376964b8af3417e8ef1c914bdf56e557;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4217da4fdc2a74472f8292c9213f875d4ca97a29cca4bc680fc404811ec681de6cd1a35163f62b2baee85df9f3001761ecdbff95f8e8a68eb451248af9bc0bf15037f37a4ea46949928ae26593a5dff63db5d57a0dd11f997ae1e85e7f1262b151ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd65a94620872e72e8318410cd4ba7da653351d3d98251914da7fb7042f9708be58aaab7a915864b27265d42bbcc13fc5b9b0fdb95aaf571ab477f2940ae3d487988aa6ce63a8e30f7e88f124b347337a6db233c4f4383e5f79029537e09467d177d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfca4261169bff78990f458398ed0bd1707fa0719dececb16cc79872c02ebac6ac99f99c4df9c32f6d4367f3d33224be46d178c070f08e4a2238c2ab489f8c653216a96e7ce0cfd2a3973e547d33dc196b7324fd0f0ebd9e0c7f543a98edbff6c19c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0a950e503a684da57b0f55e9e49a038a8619330a8366c7f9f586f31e413e4383ba61133379797a35fc62f9a96724542fcab026bf6240d325bdb12023ec3e939b44caa4b3d2407ae835c392922b1ae903129d37b17ffd60961891c0bc930d80bd62e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h367921e9127c778083aac1c1bfc045bdb35a77d68b83dd01088a1dee240311c37ca6ca24d53bf2aa66ba69cd5a7a6e0f4a7cffd11addd4c9262867ffef9b04dbfca66a414a70325ae9cd0b043826f712921da9c362296cda3d0d6b88713d24a147a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85c873c91b22be833c78e55882059b777622f5c017a544f72dd96e653699617978ad1e296b020a08ae5a94106a3b77276127ec1442e5aa54414a60c8d51d4451d1688aaef8b87b747e53c89c9842c14c9b756df5342ff9082bfea14e927f0c9a39c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b700bcc5b17e72ab772440ac5a8abd19c1084142b96a3ca06a24cf408b51c88ba9ac9043eef14450b3ee50af769ce5cc3f8f05ea55bbe143c07ffa35c9ae39164f159a079273ad1fc742df3bd98ae4e7b31fb87ee114b6ce32c49529e163b1041c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2829be7e7c8000fd9f5fe6a8e4ef0a019ba42f09d09abd9c75d2775bfbf87822f2f57e051bf46e92178c7077970db2519091bfd82724166e015795884b23993b9f1e143fe8b1f5261ae1e8ddea6a78f78843b98d4f23b6e17e6cf528e7b848bbbd53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c62a4fa0f10cd27f571560708551018ea0903f83dbbb7cc4264d8f190334939e4231e0fd843961ba8c9bd40cb1dc954604f3fe4ff1fc705c2074c86e4f30c0ed6f019aec79d95a20e9c6b3c5cbf22bce4320d3ce50011301743170ce59a31eeae3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd80be880e056fe9427a56bf48738aca787bb693f27d08dd7c80732d04fa8fc1881a7e80dc8f88f984c5489c8168be4c417007d2198cf406bf5d179093064aa514749062bd0856d1467044b3a3182fb809030c88324b8e8751e6ac02a9d719a73c222;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb793bd651a40221952eb1a8a5dc4c4bfb4b0fd029822be39cdf4dbbc540d49d65a6910065586714caa050d3253edd350403865badd65d4e4f7091a9521180d85dc439107d1fbab454782bb633e1233987ba0e0932f72f41b0dbb6c9d05504432400;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h167c7f5c5614ffab7d3151facb9e989cb196d6c60b49492ff1ddd98587bcd3aac1da3809e5ad7960b6e18ec2f46443833275327d240deb3d86368dc89b23a4a9ba02f192f78486e96546bbfdc79453d50a16013beff687b0d3e1211e4ce33e20dc8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1dc4b2f4890dc2f01eeb5696314cb3836c7d782141a249ba53fa2c7ef1cccc1c22473f4294ba082835912b0f53aa3ca06235ff95371515376a4163ccfc84a1f48895a2fbbaeff9d6deae67ccda6f1cda5969dc536f1082aa66597ff21691e870bca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3513209a349a99313419f7eedfe579c099eb23398a4ecdb25fd19f77b36428ed9af82bf143676b053eacd141064593dcfe5a431a53da4058c02df81a8a8300ef3453c77feb80c34fbc945862b99882cb93cba1df16920356c00dd6e8edf7181f5929;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f44f77a6878205900b1a89413b68e70c01c3fbf94f449ff7150541afa96d832d9745d95573b2a599fb078da15400b0b9f3f2fabbf6d16f8c78d52384f61120bfccb8cd3983afed5be605adb57617b276d030844be2dcd93a695e2f5cdce5285a594;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc388913845823a0e5043b0b6d2007dfd192fff8103f296e160c5c292cdf0d10827ffa45560b6b068cc47fa2b61e17e7315fc58b1d66aed6c5797281d9bf9d5679d2eb4ee27c8bed1870fdedb694e8d77b2b87d9302731eaca48afe7fbfea05c1c2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb98e20462ee7e1c029a366b825289cd1b5aedfe7a0654d7b77d4ef33dce8a1fbe6b9023b55b925aeea99b98587ffefd4548aa34393b872a42fe84e47e5bffc4d14f726352cd2b4d81ca35855fb0852a91f161d849a2773c108d17aeca985de9318b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6061cc3af8487fefde25ede7829f7eba0ac448642d555dbd63c9bc5f0a86baab27f51e756b31cc8fbbc33165caeb6bc5d0f521659170ee8470d685b3665b7996fc9277b443f5184dc476ad6a3542493f5a595025459d5760425e6a6c95d1e1419125;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48e2a1238aa4e345363857375ff987a8db68d6228e4f5c6f9ea07f8d4f0c1bec52f710110e6e5daf4863692b70249494349a03432138ecfba76fb070c0b96cd53adb8e3d529ab96d9c2920035d15fbc5a51c312fb8098b293543f855150f825789aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6a570844fd5a9d2ecae76e168d011d8406e20326095013cf07ad6367c3c33525a829a71c2094f83b0bd022cd5d3114ab605c25dce4d3a9fbd38955fbbf8a51ac52eb6fa5820d749aedcb2665bb5628dc9bc7295a89ac0da730b6421fa77ba4ed114;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3db4182e2a86fdf1ea5e2f08df0ec67c7f8270a6231dab4ae671ee68b3b3afb4ab22d59183417438c41fab241d55d876052dc941850d82f6ca403a9540d573ea9f51b166116a7e26b955b33620a62a141aad1e6f9cc536af28aa6a8c9bde0710a4bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83cab4d35b9d5346f7a42b24332aa78ee476e9327a08c18c39632faf3d2d8b5d3373a944b1135674b56edb61b2bd488bf1a2b3d050283f88ecfc7c5686b54b1814cd5bdc16a7484aa364ba13629527cf2ce688df05976239020d207be7a5190ab2d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21668a34c6f2d48d287c404241620a0ccb8453db25104e7bd9cd5f1361da14dd22f505b5635ca7803ba8d3d6124e1636f8728639c5c9f4a8f802a7ce2f55e0aae671d3233aa3e738e2be2e0accba37fb82edbb739a989f93ca228ad4f50923c9330a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd5cdad5f344144e8d980d0691f6ae901a402410e5be1417d54dc84c4e70d93e37e7228b67ccfa847de7966f387f658bbecd0a55d0151ebf807a34772d1cb6cc05653e36ba7d7496de5fdad47758347fc7ac2bb180dfd8931447c3c5c4221f6de1e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40626e4bfc00757bd6e89704787d35c53230cf2f12a0969705435e8ccf1dc227482fc9e7678758fc081295794b84e0cbf73bed3d6cf9829e1f10b1e189bdd49a4dcce96e5aaf9f540f8332a475c6e57bbd43de30590fe3d1eaff8e15c068753a116b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97873f62717e086eacbf276ecd309f3c58b8c9e954d7deb6a98c1238a10e941079ad93bf25c5d8a5b406e39ec6f21f56eff6c27d860ba3cd7389fd734ab20960ac78e37b33d2e1625fe4790dd09a17f723b43c0756d3a329b8d30716ea013cf2d522;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae440f45fd70314d4eaa67940a9e7fe06e7544f31a7dd3d74fbd13d2e1ac8eeb08dcb783ade4138e5bc141c0f3b8f0bb662005a95a4817b912125fc3a4e8c498e29261f7e0052fafec7983fec0d707eb8415dfe0aa1adc01d9f72afdc495e44c3e98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9133f6f05e035b91f5cc76b001f8ac1f94d51f17a2284cb1364bafaaa77ed505a371e0c6e75c93bb15a855e00a3267441cab2b30d6f72cbd36dacf77bbdd0800057735870b1c7160713258bc702f1094c6ded006cd6f65db81e503d9dbf5ea6934ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd388eca1c59581e7f0e5262fd1cb6df4d1ab3232877b3fc116a043a6ffa3bc6442b15991e96f3e9e55bf3203594f0c0fdeb1adfd620bbabdcdabb7932a33a977958a736c4647678e0da455ea856b9367e3e1eae43f9b4a2dabfccf81832c5f000bf5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb11fa0246247523903d07e90e61cdb293172f4b63fbbacf1be28f355967e9e94fcd55825b0b550a6ebea8c3e67a9f18c1606c543f32b1acd3ac3d3978a5e940a2865fa667e6a3669c91d7ad76bd2f28b1d11d78ecac00af5f4774e0ae89bb2da73e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2313ecf56ea6c9b6020ece7ecbe7f04dba49324e21131a455fc9d966d992551c20a425ffb3f80464363ffea5988abed17119ff76913b4614ff3e0b904537eba2067e3a1454a62bf2685e89b7de48157d4c4363628e8608f45059b7dddaffaf1a8d16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23142dd8b36be824168ffdfceba8871bc03b4c5f3f023c077b714255adb64d29a2b4177fc084b9b14e6b13172f2d5d7da3f6390c70384b845013a9baf3c30759599d480d1efe5a836ff361921312321dd45317f3795451cb3ee825ea9fe847819476;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heae45e7fa1494cd370ea06d05de482fc2925c9fc9cb1ea2a6d0a2364541bc299168b0901c3551aa681c20dca7addeafd6270b049a631778f6c59a0aec5be7e3f9d936d20940aec625eeceb445d1832e74d82be4491b4b90421c9ceb667bc846a0f50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h295555ba81cdbd007aac19da17373ed0ed8b73c452cb8f094b29d28d2adbeed2650c405ffb57a11116974cbc124a2675f3bdec03f6033f2c466a1c8e4b15a8ea14e903fcba3df9d4a2a04da7a9be3e1852006f30849c0f9469d058a2b7e7369bd330;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65c426259660b766656b206c6b4b331564de310c89be4caa9dc99a3c57a93f47dd593e7c985ecca0469c45efb0b664da5ad540d89c76cf3326fa784e47083f88ca4e813f3d5622eb83b375939d7a639561ed7343fef10b25ee50276793aaa1aaeb19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3e752bcfe6c7f5acebbbc6a26b40cc93f60098526657ef4f6366d5b43f57ef2b937af5a24f198e4bcf87540934d8c1733d578f22e80dc628e79f305283cf9416e6d80c633399747bb0a7d48092c8916c251989f302f2ac059c11629154f0dd7d86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h210e0ed2e8a358fcefe049fc668314a49a9f1128a94bd696839fb550739a8b9afa6c3db87ebb11f53566ee59fce45a496864329214977d026e9693ff2db6b9eed89a8901a7f0b7950d3b64d10442a2e6f2b9ccf2cacc83088ade39d3fc6b61cad494;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb81190fdc7a2622da8ec05403cc153afe44d4f0c4d86a50710aee2e3e3ed770d0ee1cd40e7fbdfe5677078cd780c6e77913d2e828902b9fc4e5333ca7e2ecc4a4cc16be349b87597f7a38640dbaed64564081b813cb4ea53b0037df7b5d4cfe21fe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h987507cb160c35b9e7609044f078693eb3573f6188fba76d4c42da1065d03cb67c17f3e88ca038bcc9965d6c3fc137affa2af1fbb651361b1b16dcf56a39cf1a9d6f585eba9fc464ea6455bfba1c9f804464b49561eb0ac626e620cf3ef6c686be19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a00a5162af6de3545806db98d2b8d0a60c0d3d90a04d54fef3d30b2de70f1c9f5c5b738cd9987af1d2c6caedf9bf8e6c8b5394a690336bd5d580ef63db7635e96dd4b6d7884cac0d37b05bafd4fc81981cba1a30d258e6b0ef27341f51cdb85c80c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6969252f63b402cfdde48337d95cc64ecdab1e2630e59453d5ff0ff5d58a573bc6efb4f173e20908c30083df7b396afee617879962741616d12b2c037e9dcdbfff9493bbb1b0e6f27a76beadb05d0c6f0eb4b7b2c792043a9d6383eaa3ddecea5665;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff6b5dcae0286603ac1c5cdcc286cb96537776092fc3bdc415d21d115c0a20d21b9c2e4627f75b54ae7572633009b14f9a5ebafbc64bb4fa441fe4533b060877a425468e5bc3fa672053fb5a8179f53c0e8748e9dd6867919dbaccebcc254743a1e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22da65a814ec68643879966da41e8819e729c9885615b08e9a402962ef086cebe5b411094a5897a48588e523cb9a36fa42574b40129cc3f699bfef4bcccba1de11282a0d8334d6c353a274795f388fb0943a3fc98ef19450858d3b334102b7d01d4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fec7481a27d46b8426454523ef942da41d3541870dec0313c50ab6cf3ac4561719acc0194bc4093619cfcf96fdf9bd139d5cf7e01e52a37474176e559ea5c4353d943f472f27c140bc078b15df9ffe26526e8472be728c77b9c6ac3fbb62511b9d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73bc2fdc492285f10eb8d65ae16788136d5087fc1d4537257f00c522f9506b69fd8ede245ec96acbfbcb8a91572fc8dbb58ec8b6951bbd81c8015e084162b65f1907b6858c78464a2462e1986632e9046aec919f1188241a11cf4d59a1363796c995;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e5fe4e94781ac6f0e9103ab02e1e7c3a02d6f4980038bdff4c1549e02725a8c6b1ff87f376d0ad610f2eaaf000d1f59a2620b2daa2ddf2ce91dadc2426a1f7ab395494d0f59915c94c1eadfc774308d62d9884999d414364b3d772e43a1647fe55a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae99d96b3394028fdaffb0c45a806db5f749cf767cde703fdbb74cd8a037b6bd73b7cc2ee4e7e7b67e79cf5f9f1332bc9fda25d87dee89cdd93ffadcbbc09889df4adf229c22d0a5ef242a2ceaea59ed875e11bc7318cb1e9a6a80751f14505f24b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffb8467a8199d3860ce85bb92761bef9fb9c00a401048d2af1f7bcfc4be5a4430f19c42fc8011d667d889f7898a115b56b3ac31808e00932edf77a3b8e283a8d7dc6b324bf3f3ff159f958f0c84153bb93b1142d70a271988104ca6bc938f2e4a8c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haff610cd4b3be34ae26165b10fdae945aa8012e90a472d92f35c521351ad2f22d809213d8da0dba005303a140221ddd0fd03cfac52b58e7ef75547908c23db339ea9db11f2dd1edc3982aebc8e6229100e2f82d8d558f931781897a3b692ea9194a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd344bd9b7d707318b15bdb9997932ba795a519b1e44214e6d9ecf2a74473360bfa7e5f772ea137fd0ed3f7a1500ef75868d908849f48e702572d7492b44a3230f2bcf8835dab3e400e3f35c2f7e22370d8e332149070a01975bde90b214d73d685eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8aeb568800d01b7a4c3b94230e09cdbdfb5d4c3d5917c309878817a11ff934cceba59c88f117b04c43fc1dd170f0840c952090563fe7fa6dbff96529f6603a3c3283621091c99803b33ad28adf7f3288b4fc85ed598028e3a6d02823b0d9195a8982;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba3dc052d4186795e88e953c47079a8cd7a914c8a43ba9b35e712c524d2df06580b4a7b123ca2949a50ff7fee1be80620dbd79fd7cbe336500208e4cae7ca63b5ee24dcf64591772ef86e9e9afd58e3c0d7eb2611a1b57e976891587e07bb2145254;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28ed33ff2936382887c9c0b00ff24f3c8a32d9af993700cee15bf9c400bbaf5014570420bbebb78b2fb0b43c514ec5f18d68c614e2ebbe6723132b0a023428614da637c2d9c3ddd86f180fe8c0e1a3be795a5a7dd8d70ffa4148abafa963368b565d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28da680dcbaf2a4f8c5abede80809f62b60272dd4b466cf978cacd727c9016a1f233f2452d597ce3e32cbde222b30aa936adbfde1d88d0c29046c0a2144b686bae0eed7bde498535b6f7ec72f24fcebe9b78f47c7040e2db290e182462fda372a960;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b31ed29ad5e207c9334ccd5e89dd3a752d5d8d450f2c0e2acc194160ab719bb385884fe6cc7e6a87d31de70061ba2471bdc8fa01663786201d9938a5323e25f1437c700e703c1ed3bc17d4277d20c5b9cd49dc7325c65fc00d76a72f76e572a1255;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h146d0322eaf8934245f1b1725316727a4eb8258d8c6fb05399d4e20a2c04710189c1ff99801d980ab0c0dabe31669e75f6b1be84c76c950fa423a01d86d24bbece7adb1a3f30d35142c7b8b020359d1eeeb7ba198d78e6363b10d4147eb278ff2d9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f318b755a75a56ad0ba0aa20cf84a64be47f7184f2251e41d727ddce28a0c5efe841a36f7d2fdc1d08bda322d811108b3603bebca890cac9a1f9a829c5c6e55b4388ef5a7aaa79adcae57b4e10d95ab0d16aad732751ac5c0bddf4f2c14945d97f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h191eedebcfcbb71c09ec2c372e2df25408ee0dd7d038a9687f56ba265a7c041d228e2a6e2d033ac9a2c0ad44e5aff342c43e5f180f7bad7e8702662b11b978f3dc9508997d2955abf790877f63d4412eff140cf4309b661c4195840ef4bcf4480c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb64ff1ba2bb77a11cd522cd386b58a74f036e240ac13057c026fa331e77d6d397d772e3dbbbef5dc6caf2bd0db5d2b2ebcc93092100c531da5954587aad0718377ffae83db98bfa6bf4d045aa510f6f7050ca38e60b8cfbb2a3ac0d3859c4450b6c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha628c45e32b895f590b239cdb8d8549388b199af6ff76ae8a76ab494c03fdedd96b5ac40e4255dc7e0b4eb1d7287c5d2cade4d026fbc40c9d691acdc5ec56700fade99528fb9eb5cf8318b8baa59381ab30341e9b63fcdf0446fa2523c058645c27c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4513cb717627e245f97f2539e46448a60dd4c314671357d24af3fb90adeb0946ed924864980bdb9a917426a7cbb8c6282aa560235179a6127e9e25eac9c391e08f3b2902309a855d7262bef9ccd4845c5b56a3452812de75d368e1c91960bedef64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfabb40f3a0c631d3c82ecaa0dd7b17d5ed19ec12f73a6feb82fdd914c9b46a0ca741bcb86832f0eb1086e3061de79ecd96b7a116d69e889a9eaa0c0bde86bfc8772865e68ef558964996b349accbc0bf26910f7041132dea36e65b66ab57b5f12b4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d3e9a5ee7efbb35f75ebaffbbbc0e5054a89e00f9ce1252f42186e824079e09276d12e1c592a5cdf610566af48eb00e0a24b7984ed76ee8b787ae68d0dae779ce858ef0cfde42e914520d97ac9f9fd150055f085d1d128e80a9ee9e381b6687192e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84ba9f64ee60e0c3c9c4cf11848cb2a62ddbda6cab3b42c79bba6a0e6d6f6078b720163a8479ccc7b75e64924f7997b3f1d2e76a803a1f75217ef3f5b3ab60291eda01b72fbd1475ad3ab54633ee24dd77774f6289763a76e8b5753ddb8cddfb0c78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbf935632accf65a6b4bf2546ff66196b7dfaa08e77ec72de04b88a4c4daff7ab31d5940edca49b3767b29cb8566bea487ce8feac0db2d6d0481657811fffeb8fdf84d684edd60b867b2fba8dc7a97c8a12e4d4ad1c4cc97e83b1cd294b5927fc71c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27b2567670dce599bfe6b4816dde7e16b0247b60a330c710033de43763fee322281064697afa7660b395d366d7de86515d8d982af08381a285589c5e5cc64ac9fe658953f9b5e6687b8b578ab1ae4f8cc4161c3bf4a67a1b07d8a2c01fc07ad0ff89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h272a7a0c2635b229852d8a3341cf630549770e3b3545b4a150e7b34ae3b9a14580595f37b03a540df86265078fabeb2b5adb3c57d3f587aa622595edbde4f0513d25e3cfc3683bd5d4822a831c494fd24b746b26daa6499753d09d99d2f87ecadbf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93d8a42080407b95587bf807a1524df23270b2a0ef74c2fb86f795db316746f27fd31993c4ce88f73e13f4f98629a4562e1521e29ffe059de52d1de135e31a07d6bad241fb1407f0e89bcb079fd5f0fb92907edb8b33944a79ea18653fa8a121ab1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedb8471560dc3fea186d617d79feaab1a94c98505684f05c588289dc55fdcea027fc7c533de4d98b32bec93398ef971c992ab6686374c591edadd686145e9f22cfa6b29347265f618ff773aa366992da82ad14439c656715e601ebe83685fe510320;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha43ca896d15160a3d74783390078153c69d8880e7e2c867b6f850d11a16ada95670988cd2670e8c8036315ba0c74e24fe248895d38ef6e7537562d75d3c2a8c356f9b488cf174379f3243619f39852f455100f542971cf66ed26b05aa2884e4c1cde;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc35ff7dc18bae77586bf2201e747a2cede80bdac516ad34dbf01a91a70216332d0fcd74faf39dfc574d73bdd9ed4b529ee729e4f0ea8b3278516b4be922204802fbcfafc7198914677dfb29b278eb0df6d2b87962a877165790249c6f8700c2e14cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb53b7292f109fa2239adf46e4401e99d61eafc2848f7a84b9352f7a86715d1e169263cb3be5f4d6c9e673e16059cf3b631ca43110fb3b40c8dd11ca451396145c773d2910ffe82b7e3912d50a842aa340eb466ae2b4c3caf20dcb2afab25c794f15e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19b905f9c9a38b4e93791192443f720d636ac592a763d29ddefb3605f85403efa19ddcedf7777ff43ae3ba1c8f8b5757f7872fbfac35edd73ab60de73643a23fe585ab421497d8ac1d7b8ef83465edbd6b78c5aec15f42c0885100029ea02e084dec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f3d84686b5bdeedea96677bb744e9cf51b5174d4fdc2219fef1fc3ef677a917cbd9254af7a848da8870cf2877051326450a30cc0875af473ba52ac4dec9fe1886974cb3607facff9296f604110c1a8fa3a4b17c553857104ab72f0e6ed658d96ca0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68ffadc92fc06845ed819eb650d3bc6560f188c1676511bc75bcef2d0c2b59846edad97786a1fca6f8dd56e5f374bd7b65ec8ebb18567b70752f3e9c68ca8ee62012c9b313329ac0228e1bb27f60247f8def6dd961a7129a19d4bd8d8c3d2b930620;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c778154c947d8de5a10e4e7cdc8e41324af50b9239be5222a1c8679af42a35026eb6d35f3ddb1ac9801d90e0d817625ac0325b30e20a4523b8d56beb0ab6b9c5a94f25dd2b2fa2543051136256e9ea9e7b319b839bc5586d56af09285633fc7b71a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfa3e0235cccad7dfbace6deb20103da3154888fc72feb8a002fed3c9437c74da2f6dd141d57b01a630eec54c216a9bb59ecb1a152073b02c66dcec19f2a8e9e3bf10fe3d4276ce52955e47842c48aaa6d2349191dbca4d153fa6e1b964cd18b7e22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h829bd8e70e6eec567c1841ad652697bad7c3cdddf963e04bccba8012a5933f96d8665d0bb22e8cb73b1c9095e81e20a5a561fb5a87f86ad2bd5152f28fcf43590e51f8e2a7323b38afa60c1d19f13d11d7a38941c2178e58b8f9158039978ec76cb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b107e1c402fede07f4ab49d9925c7a41bb7f8780891110f1555ab6b5b87270b8996764cd117610845de4d9ed75d62f6665497a4cd46874cd02fb614853ee6e635e7800b06e4210d116c42559692514b4ad31b0238472d86343b4100071341db4cc3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7defbc491cc71a47bd1be9b44f04b81fffa488abd7375a3b09729774747f34db8fe8cdb03a466e41b32cefc9241e8d2b5c25d0478918b68018cf863326214065b1a4c74773d3c03812e5005500002559ff21c09def5fd83f3ad455dcbb0423df4fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd70d5a0e156dcecf87a5cfddcdefc1768a2c6bdeaac69396c3236a369d4a3124e0aca50dda9ed950eacf0b7fc5249b03fb22544a70528397d2e21d4cd6f4e6722be338337ff186a639e4483308e0ab3a7968b57789c855cacef2398042e79658d314;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h535de4e24bf2a30d1cb6a1a2b0d30de8e562ff2cfe5184654618041ed90fc9c19db4845beca81a023891e742807b04f9e63e35fc2d8660a585871f8259b631bf53a91dc202fd4808779fa6d008320d2cafdc80c6626c0d6aa357e616ac71e0eaa1ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd0e5da0868171697c5dd70cab018ecf1da3ae2d1161b1759e796c7b5f21702b2796e09333f3a1683d1260cf2b32a318b4a7672667e4ad963bfa8c0803ed2656b6a95fb9b770ea1ab8f1f6ce20d61f7b267cf7c29b0953a7229a54ecca8bf66c6a45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8207e9c16e9168e3eff73216331954c0c1a760462866a5379a71fd6f1e019f6a55183b9e1f76cfb6f3b137bcfdffcd9bbe23c74c29d23590b957ff02596682323809142ffb84648c81fbe6bd502c8913954e92654d4378ee6656f4ebd2c99a3303b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb35da9d005ad8bd58fbf037d77fcb4fed05d80a7d62fbf8cda7a1e5ef208ad732a408ee507225b4ff58fb8b7681a606455ad81c1e426a071d6ce3bf76cac763c7c53793a904eadfd898a5ebb79b2254bd581bebabbd6ba1294a89fb4b219e7859273;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1e2541139e6f6881202feed262a91ed5b770a53c2690c5a654e8b1e25b42fceb6d9cbd296cec9fb949c0f50734be9fc10613ad4419b11158aabf596f08d229b3b313a44fa303e8ed8bde90f4162d86f97e9d821f4f5e043f0b818cff550e50c4fcd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf320f92122d4318560c8b2e16377dc35c4284771608b3e7d93dcf1b9b87e960e0b7a257ed29ebdea865d990295f812394595d69caa54c38278ee6ec83dd3d779909b7c6638e3d7a34ef0aa5148ab1062edfae5931c1c750ea582fd369ff79823915b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5c887033fdcc0215f6130bc815b6be840c09f77151b2e126521a74d2a46e35f7b523a4a35149d4bced69620faec71877299558e7f7295d0491055a548bdc04fe6bb3de25fab956b017287450d3825dd8d8e38d7512af3d206f0d9e8e97b565cb4f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4fe96d5690cb4913a7c78334de05e56e6e342e1681fcdce54c0540de382a8e7f5b97f3ae281a609335f1da3ce0c455674af01a6e1c778e20adff1a13aaf121090b06953f6ae3019a52e2c4161a7eca2b2e40c4a25540c50290ce5c60fc8d13a250f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88c3ec1e58bffe5e5b28d1d9bfabf1e0cd9c53edc286f46c318c2a9cc6f416e68a924a079d43093f8777b3d2bf716061bede32cf11c1adce9589d9523f6b331459e85f6a34fcc3092df91cf80be27877a52bd60b5abe8ca1fbb918492a86f93d3eae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59532a7f7a2b62d9ce3ee3d63fb25c87d78d12a0cdbea70f0d597eb107ea97737c038127494f3e68e4e146eefe81ee7ddb1f936950c2469fde032fd011d8e7260045b24ccb04d9d5cb0ea8a73a197e87a3ee9443533b1bc3ff13c6e6a5c282278e41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha651f2f1528ff24a0673d78932f825b5ac69c525bea214b0e9055ecbdf55df3ca87d977aea51a295b0e109157bc30c23002f7433b06c9d443f503990f9b32165bf9245b17d65e996048a2117ec44e27402d307ac4608f83d554b98c076559221a4e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9eb72df0cad7f6db235e5d2b8ea0ac8dbd666a3f61b1363e8c90418021aa898a68ea38b2369e5568916d14482115b4271bfd6722ceacb1ddce9e70b0f64a0111ac68dc9bbaa07924915a88982f1e14f123235d47ea56706163e4e7b6abd7333221ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea93f9e5ce0fca513d0afab92d7671470b5671693b412ba4ca66f4b3c4a95e8063b266878b1011c6dcf45362fa714fdbb908327268791c7173046d0c9a187cb835c26ae226781ccd9594024de15f721729cd7538e8c75e5518c164b7964faaa30214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e5c57ab218db4ceaa6a63437211c07efc56a805d01a23d030103de922acd87074d28b57b639e8a4baf23e284728d9f4320ff44b6868265c3ee5815db56628b5f6fd1048ee1dcfbae957da830a1437418df5acd402242d656a1ea4b3819c3b353333;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51122a4abc9ca62d93a644e7bf56de306d781e05650957d9f6eba6d9654b425e6f727602e3def120d529bd0217d0bff99574ef325de82e5085fabb673047f3f662162758d67c16a261aca91877a332938d2ba55d9c64e94e0f9e40aad40a2975b9da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c7f4d862c8c70f58e366a7e795c4cd8b71b21be04f471495ee2ef2e1cdf5bd10feea4b0315b234d487a2ed1621a16abac3d53176fb814d2f7a1c9566ed5a11184e88dd7b847fd60715c6652d3f723725160d5fbe527fa253e69cadb950036898457;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3135f57ba45f9d3639be5fe65aece5a1e6949f5ab77bf48f635ac923e1a0a47b529d78a5bbebee62aa592c722c0c55ddf797a6c07c35c4e5c571053c631e5dcf9722c590c4867e1ec9480cc176fa891f0c2fe68436803cefd938e577d1a66cd50d0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10f6bb6aed497376adce914b784c13e4c853e09246c865968a508c3d5222da019540e61f1b073332cb2766fa000e6efcad9ebbe17e8ed1ab492502740d6d1854840a8492668df2ef3c95e8a76a331509541461a0566c7f848696d4476e90de02f83d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19e13e13565f1c40163cc680c335809274e85ed39293ef80b66483b4467e0fbc8d2aad6484712791e1d92eafb96114f2df279949ba0ba902d0cb7cf9a4918b3f79298806a958102b3c441eb100d654c78e95a95a4e1b33cd4d0f516119bb8b977c39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9354c49750c49abe21e5bd164c1f69d38d2ba213fb9b1ab75977a0c63b174ba59935d53ddff3b5122cdd2fc74863bf61ca1c8e78ebc13f7d971b315bd6fd528f97d08fb37899b52549155be0cc2390fd5d34493d54d4017e1607f4069da8e4d048ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc945a5cbca9d5df567f8cd4f8614a1cfee20d180c9e4b6a275e6a45b92a16aa6fb2cd77e714b02cc7f40480b3593bbc2ec5955f9b3537fce2f3381512f2a5401411e9745ee8f38f1a000ef38abb5b2e87871345d568dcea16e3a8d84eb64727eb38c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h505af80427e21e930ebc11afe390e5264d22b3698f778a1c1351cc132b85644d8cf6a80c8602caef7347a401e2b790ece9ea38097c5338e8b52f0871271e1e68d6fd91dedac4d349ad6b3fe52627ffbac01a1c204e3bc3de19f72efe76e51c0f5b5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1ce51d319a7a0cb2242a579e8021394196112adca280b996ca96399c4266a1d0f37b0bba33e122e016b50d8fcc0005885807691e5430fc108385e17525c0d5fa52a1d8c491b2bc2e005f976b147db8402213d4d69d5a9bea5e4e5978cd8d610ac2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5647e58cab3c79dccca850e1bf203cb8127660ccfd4d23abf7f04ae117a09ee39eacf6cefcb89b39a05adbe718d7351a5fb8ac928180f80cdcc11153db974110d312c70ec75463278fe38741e88f65ea2496e284bea22172b5b991685b261c787b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52fecc4c42ce33a0a5bf9472eeabd507bdf58d3c82d1704701568e23c6dcf7eb8b939c19687f4f3aea8ce02782574cfce1df96104368156863a62b22da68b604ecc6622431d85ca2d2e01780f7e92c7a991ca6d5235fadee790026dd34b38bf8d086;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h793030f0d6386f9b0af67924300a55f7289a7489ba71ea459e66e36af730b467dc86c6e0cf067d0effc309d7faf347b4e6f26126f12165bee92f809349e3074459f04e5c70b624c17a6494a3c4f0db9203f5e8db054ab1fdeb7b7227f7768a936cc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71ea591688b610a0b30fd498f850cb625d90dca4a43be1d433b3129eb77e174f1ba7e75e768dc8d6ce15713e7f7a25be54ad767a6df44fac7a43225a3db34142d5290b55738a5c876f9c3c01afb3fd19770efeab7649edf55eca9a2e275351baa725;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dae1ddd03ff06651687054f84fe24729bfbac29bfd7bd04225f29284f126d1ff98e651246711fd145eb189d51796540cf97b6bfdddbaffe084d2a0045bd9bc42c0ce071ce107c1badeef77af9a08e851e5ab18e4f5c3c53110ad06d411e79e62908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h852c93ed4c734e0f8671566ec6274e42b2398c3a7bfb485356bfadbe3976a494a35017910113418b510e5928bab4f16691debf191790fd238b005f522acba4d19b7ab222105781f4a4f120fa99feae7ac3ff4d7ae5a177f67fe1e08d0ea26860acc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca2523ee1631267d327a3254801550795f9769b0f71022e9bcaf91c33127db7bed1ef065f71bc5faf6b75f9c9eecfbd86059bf923b409c128174c24c5e8d5062663fdd9fe5a7ae9ed2519ce92abff1722f043c8e241b5e31830718cc7522408faa79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8304aae95efddcce329356f00ef8281d43a20a6efd7c577667b3074a33f193fb64543d5246481cb31f6793441411e0fc5c6657097ae0e94dad88653efa746d314d0bb30b639939417001a6144864c040c4ebf08c5daac1d4da432997fd6696cb351;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf084834640587c8f0c48197632f1804f6d215f326c4e8b3aa8077d46362b538e793b13c5aafd9a1a1994fc29e7995ebf9ab2530f751a4b490eb1d05897c988a2f83f58352cdcd109fe051cdeb9528e5ec291f4735e5bd712ef3fc826bad494f139d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa987261736d1349c2c1ead183279cfa0442a9c2d464621715d15d131d24aa36ee262b56789003ca8e448c55271171aa4e43cbc831d1463cbd3f2b0d6f586952d892807c5d84a19083b9169b7e4ce8f272389131cf12408525bec6b3dba1125377d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52db1a2065da69c63274fd05a5c18e2318e5a72a2d8b003c67ec001e2b54beded6dd02decfa082c5d3761b628f607b8ca4a7def22e07b23595b4ccf5519ee9c321f5628680807359ac169fdd7dc0e84286ad32eede7f93f7621bf2cd9f4a21d0dcf7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h239a9072b7bbd1a1741ca5cdd3891862991457459396cb4288b49de7c4aa16f6828df31dbd1db907e5a7c93b25d7909be5bb9d90f9e93ccae78de8aa58daccdd14f35e39aea3ab03dab5a44a39cc5ab04ccb0a3cbe748aab3cb403465f8411cbd7b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he34e3a5f93042e6eed59496b49fa1e2902ea0a791caa4771f85b27c96d5db514168aa27d13c96564586c0789828a48f2853f24758e9294a27851725dc92eb16c78d8d5d083af52e56da03d9a4706f4b7f25ecceb61bf213bd5686ee2d10778a810f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8049f10b9d48fcd20287fb48ffea4175d3c959f231f6f13907ba86d97b3cac318d321ddce610d9f493346043ac3c84ec679cdbfe6cfa9dda80c8b08987f71fe9ec852fc70f82e2053c19e0f7ccd32a39547f95d88da0ebdebc284508168de4f304a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h934f0580d58859eb1a14f8a840ad3822177168bb5b36a5d05fc910d787d321aaa02b469b8b734e2160f8862872429717ef262f41a8309fc676031b213a7847225413d9169198c9708ae27fce3834389576378741f0965bf0b0cf162b6a6a20aa4b69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1f6a41737ebf6719eb9ac6ffdefab444fe075ef9ac4b94ca1a713da7f87ea433e56672599a15e8999c01640dfdf3829d9a851441a4dd4465821c673eb74189f344b4d4941581943f88855959c31254909b48384e5524254552be730985fd3103efa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7009ff9de1ed6f36ddca6df35cf0726a8ee12d6b150eb5fe140e40e5772ebe5ce4a69e31cbee946b0ebe1eb14bbf44349dc8ce47dd56284027a6f200a25ee3928c61ffdcc572f89e95e674c4abfd7cebf46b136e054488b1b4e2e6e04c368b90335;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h864952419db4d3d12b3e6ff8994fda82b659ebb2ffcd3bf590330de8c164e4cb6bdf64a99d3e28a42257448b7bb49ae4e9903570e66c97f66019e0f455e0fdadd37fb06905ffa14f8a1217091a694c9c3196f0814340fbd98b181cac50f4f8127ed6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2a4fab0a60e5b00039a71ef59a8e8b1b09af79091402d93571953d4647660e44f65ad7f2f5f9d7fb9dd3d65be6d91b1084c7f277eeb5c15dfc65619aa928b21ccc2a59d400265ad632f0a3c9e8ea42bdaa80728c27565d54423304dd2aa3d6e7d8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d478b98dd9d1a45368d1d49a36e66fb8947f4d4de426aacb5322ccc120b8ecdffa1ef8c660d3c591a5848b18556a1782eeabd136bd6a39005b99c1ea67a162320983f081e5232668d4838c397f21db7db3d4e8f192914fc159274e73075b4e4d305;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8816f89cdeacd59d0a08060d0a19323fef6ce7bdd777fbed503a36df833a89ef2466979281d90f65ae6165990cef530ef193047b33cc76e50d9cae5e6187f76d24167d5091fbc74785266f2a4d75e349cbb5bc79595cdd6fd93849f5cb0c94e95a6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heee411bbb0a1f04113a77f118ad9e3491cc2114d41b118d0097629245117237cb1e7f010f95af8563132831d659af412b9f633656dfe32ae3bec4838eeb42526e66f29c59db5c6363f907b845f213abf0ba353cac4a79a4952cb708a7b58dafe59c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ae8b26c409ddc98fd8bb55a7dfe855fdefc240c5424cd142def699841e108ce08e46a867e5d7c2a292a18258ee33ed89b2da8fd0612e0d188b252ce3bb7efe0bafc14b28726c278f2e0779d8d9ffb6ce354082dbe687af8e3ef2e03cfcf3bd7b4ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfeeeee8fdd0de1e77b03dc96489ccd53ff0ab6abc16f7f77ef6d853612679ce82094e2cf187c4674daf7d7bb0fe61900b0707ea57baca3723cd766fd3611cf86eb0196ae90cb259ca51e2771dce38e4e5dd780cd93a404785476229d928f7e4bcf5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62fe70c71a3dd57fcf02279722cf74be02572e1c991cac913569262794296c4078ecae4286b942fc0c316927e0eef4be2225f20279cf72738e7828071341a3fedf3420c2151067d9f76fd7dbea503c2236aa7f7e9ab33566aa6d120e1885208fe2a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1980de45427010994c56622716d00b5e8b6b12ebab414d6c2dcf235bef493ba3e2c6fd3b68efbbda82d0093f7dd768a56314282a2b7a72c171d5fd2796c641d1cd16d20a7274ec07b11c2f43b1e8c632b51fecfdec09a2abdc0c3dceabd22fb692;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce8d720608fd7c6b4ecf185323bb57832a92677b8e1a54fc73d45e8e9fbdd2ea98aee5a7778a16b7c0a95ad7b4280c1da72bed3eb0746154f6e4cbfa52944986064bdaf28c29c7bbab08d21239a7da3d989d1acb420f471ed921ae96bbd9d463d9b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7f50b7d0f20191f15e5ee011b4bce37dcc401bcb67180f67df3d78217975938725823cc2cc7888f82e4e8728c39be0265addb8037cfe2544ed8205adfcf741aa3c7f819131e29f5c3f36233ac8927f595c485b4138520503473744daca7e16ec82a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf66d2bf69db3ce8d6170f663b5e539d1ade494af6a18b25428c4dc5da1088c20511a1f95ff6f3a9840ec93b869e7d699195301ffe0f786380504e6fe00fa86ca9a533ffb47b7be3b10e30d020af50743ecb233dbf5560bccac1addbd87d9acb6c024;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haab7e7632896c1d3cec6da2d3a51f98c204a261e2da79e50077daa0918977b2d5f136c9c821d78927996190670cc92bcd32851d09d5c7fb65fda9f0a6d7b2d43183430c756c0b9878e11d141b2dffc7c844f5a4d23fb7b8ab418f14f3ab1bcfa04e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc707eafa6a4aef1bb63c5da184d39bbeb8534e002747887db29bbd23df4545e5014d33bf9af7b310a174f643999cf8e15e062dde9526b701bd83ddf343f9ccf969a896cd51ae277fa84a60153af1c67cf11431964983bf392f6ac05e3204b76d22ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0905029f0050133541b211ace3b7217ce5ed0672e3b7b8a8fa537d295ec95c7487e3e5ea672d824b1f515363c952eb65988b8a5c863e406a64d7f346667950073429cab7bbf442166be1aa81a8aa548e8a30db636ee3903aafaf61eb633366e1381;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a4dad1326ffd4cbc8065fbf2c633dfb789c98ed9c1d2df533575a2aed27e4b9b247d16433ba29492500edf9fd5b89d688ce4bf055eea0dd4c6bcf9f27671daf95176176cff6fb83849a38abf170a34ff5d4b73c8e27980ccb6a5083b0a2a8b39d27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f6b3b788bcb3b5d3a472414d7de40774cc4510a98787ee13a29d23eb1066a1f58135a3df7cf9e82fd0db1a2016455cfc1bb38e7eebb8923e06a23a798897972129e3a308bc6bc1195a2be8446f78ffebebd14fb1bc77179508d7517103c6ac5b34e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haba5e38d92442fa8bc0bfa995a5365a516b147c4028289dcc4993d6f6c442f643e3fe319705591925c1a8907f6d31ebf97de47ecf80e1f9fe6653f3ba63161ffd00837ca9d1d3840fae2e2fd799b66d10c529c0313f3a9df70331ff789d075437135;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb314d810098088411ec13b423b071e074d6011f3805bf4b6f7fb39bb9a78e5582e23a66388893a439e7cd7ded00e64c77ca5436c8893bca33ccd6353cfc4a50d10a0b646ce159e97ba2496a9eb3b3a247f3bc6340d2540011b9bcc051f8d74a9cd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6c95dac5d5dea5032409714daa5993a6cd1dd09bdc8d6d266c182716cf5463acb1fe511302e507964bc2ea3a2d6c36e1b82daef409950bbe508a0368543e56e27e4c847423894830ef14e65ec9ddbbd1405ea2bbd3088b3eebb1b575218c84088b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b6a29a55e991b88ef9a51b150501e5bfc5fbff944bd8222939b625b1d88cdc9f56a6e8669e39db2fbe354e8175201051b4df9e4b65cc4f56306cd9525a4cde837fae2eb70777d69f4d0f9e04c1bc62598c1f946e36696a83d9ebe3450bd62f1567a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf85ecac7cde3e9402e0ea3f0b1d570a064c35f2a29d9a0566b40cc32d7319620222cc15984225139189a7e7f62ada59cec1ece3d9110663f6ddb0cc667fe862d6cc294a8e44d953a7172fbc8ccbc87578f44b1df4ba1ec0bc8deedc3201decba4cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38c62ba6d196fdc2415b89db2b93bdca5dc1476095d66a2dec7ff0a1ca464f7d3f64108661d5ce93afe65a2d05ef50c8e518795a5077a07a7b11ce2c09df55cd32c6f772f8b2c5a88b765835a31909cc2d0c1b0ad3557b9537f436f0910cbfd8251a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e92ebacb231fff9d2d989ffb159238d5af305575bdd190454d68a15287d921041ab8eda48ffe30169db579d77d65c35b0af6438b57211c1691f490694162c1e309f64736bec98a5ddad43d5f8dab6ea024ba6df7f7134c414ad13dcaa41151466a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90621cec385f6db97187bfe3749b76c58084f274a45287e3eba46ee3c082c7312fa269d314b6a48e1076e016518d3ce0b3df8e8766a165fcbf322b2b9c7c73648af793a163daec147c89973b162abf751488788c79a1527acb17a902d4a4aeca1184;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f82a01e7aa9a6f4759f831c8c78c29a095e1a6ba1f92237a02e880acf5d5fdc4c7b61476ca18ec0137823503700f0958b987bca930e6af8332d878cc2da097d8d745280fadd4084ba0b49b4611e5dbc844b1511e468bbca1b5851d6e840da9491c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h331ddeee0c8d37616ba44e68caf502cfaa49188bf6068610f02a9e0ca12e690f7d30ec56441c41f7f890b5853912f59fea7ac3690f7fa1db57fcade2d7c3a2bd9ee1346b0ad08a0b31b1ced925ad27a6b6cecba9a247db4617bed010cce86fe56421;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6615fb55426633f4b795c20c8a6eeb74f344dca9b75be92541fe214e9ad5075b4e03e2a0f8a09ac9762be6141494b0ccb2bb53ffb77f39646c43d7d9d9606df1624b6263b2a2f623effbe5c8fa13dbdeb342192917bb92e8d0982b1caee9bd4f4a8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba437a495ce09f63c7c33e54780bcab6e607ba453fbe08b231394949c3ee42c82d1a40bf795ab4550a2f0d3cc87728975387e62f54817b34452e6b149177a68b776bd17c17c590ec14df1a76b553afc34d9a37d2a6bc07653ac6f4877ea4502e8684;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e16a5a0679d898e034e4b6dd9517b9d1517e6f2d68d66259faf57f7b1eb561c73e4a229d9b251392a1e3c16de49bb63d00dc0c361768a33387c3f27412768568211fa60b019b3f877e6eb5f733a60b0a7427843b908e245beba1852a7582c81875b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34973b850570e32dfbb4c82d1b681fb9c4c2b3d4e3d87dbc5e1337480fb60d406f074cf1b74c4f8590e55b6f79312ac654d6fbd509650ae312c1887553f144384ca1bdac7f400dee46b7dc08cf36816c90d3d413076815347b15f14c9bb06d60343d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9a455c6d863813191340bfa67f8d9b41bf430d944eb71f87cd3757ee6780da4a8b6514334a143bf74dc027ab88250463e73b35c6299bfb5592067dadb71940663167eb04c89e7a54aa5a4d8d42cec6e852795dda70f1561a36c4387dc123cdc6165;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9b7802d3f9e55a707511cb12cf09c7a91c8ad70353eda7c0e4eaf29933fb4fe6d5a6ffdf8d930b148f468b62c242ea91dd98474ccc4e93919f4da84db0482147ce7c6270f2d7034990c14d751dbc2efd1bc45eb857e1aa2e8966fcc493b8578bbc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h964ae1cb60e1a877180ccbc80fb2bf26f54e4c8e3e87934b23676929eacbb93ff88798e2ce4ee225a5cb3a1bcd1c7a0fd87068875d9b3779b8c42f28a79aaa5030d65c513074d83c712df18d7736a04a31d9378d126f589422293f4e9479cdf04a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0352763562ce221a85ad04762bf303ea48641b34dfb114b126b03f42e75ab4b25d0b9d7627d9789afcad86c476604e5f4b4f0c397c47525681c75bc8bd35846cea4d9db754c396942613d7b0b7a0f9f033eda3f39c427e2eefd305598e6febdb630;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h164d30663bdfbe958c371fa51d5a2a946d48531698775cbb1b85b134234cbacba46eaf8547648a9ce54fdcda86decebb0bb3c27dfed04677daac5441ab8cd5f420b8df75077c8a3fe81b2d74734fc083c6a4584521c2a49f06d082baf83557bd294f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5abad06b48b46a159c4a361301e15ca1ea8c2be0bb6f58aaa0907b7d00edf6987f79d75d557a9921a365462d1db8cddb8cc48d3b303e6f3242cf02fb9bc3135750da8ffa5b879516acfe0104919ce2fa5af33b76fd303f458fc689e77b2a0ff4ad9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h217e6aadf2743ae186beb611e35827c418f975c8046aa38b62006cea4b1fb868774e206ff6a4e1030e5159ccc626bd2ebcfbe766d0a35876344b1a3b0dc98ae93808c9c3b42c7b3947557132ec72669b21f01da070ad030515d214ed7828f895b01f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bef3f76e867e4c14589299025506f4b74a1abfb8bb14d153edf5d67fd406e9008eb9e4466512660f3f4d400ce43fff819ced9335d28fd49f3c5943bf0699ca1e6ab65cd99fa518057ebb0e04efab032a34833f351d78d3017a6cd326dc08a860114;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a529491b4bd03a4083855ba1ff1c4ed3f5eb47946bb7ed7a5815c470cd1f76eba89efa435838fa2c4121ba465aca4e118ff98dc9aea6c5fed740c81797a5d1653b276cce1591111c55e35af25abaf4452e87ec454a97afdf82ffa638877f79d514c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h533ec91468ebf4516f3bd955808d48650bd28f308dd56d3a17d2dd60bd8ee6fdecbb8ab0e3d7d079329a27a4b0db0b08310df78db476255fc5fa39589090e9bad9f481b8c0270d859439c091b239ab3ad46d0df7bf5a72a79525325cd27bc6da6962;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaa79fbf77aea8dfe394cb1cfaa48d9662513ab6b0cb3841100360bd64d60650a2f0c345598c17be1c406e69a0b0f47a52230f8e68066154e05e4306bb008a0f264c74257d065d0e574fffe6ffa8ca862807377dbc597c6792c6f78ae39c5d90bc54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7bdb3a6f9208cd3f63b4135ec6bcfbc59d70b508768472ee4a7ab0e5740f0ecabfa91f881a8793949f26002c5b1ea4381b9e714b79306c99d029151178b4023a4090eec014e62c2eab567531bd50dbedbce8b3d511a5590a0304a4e612deed7d2d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bfaca382663f9069b31cde09a600f4529c1807aabfeb4921fd6296bec805b965c23c35de1e2dacce2e8d75497aa821bab3552597eaa94d1b9ce12f2dffa2e38fcf6fc95df52fc42c5ee374ba5f0b75da6b32db9b1e213b33bcd4edd50c5c2c1b64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc0cbf9b358ecf5c6c39c6e2445ffc175336160bbbe51bb12090ae9d0d875fa51120f5a47587aec3b4b90f7b3a083fbe8244cb56d82b455754709ce46d84f5dda547a81f62e97b5cef21509b243d0f11bff3da3ff1beda2a54b7956ad8287addae17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d97ce9338e2a2630d44213049a044c284b4aeb7f22c6f3ab7756822320073a673a2018b7c1ef254e2d993918fa153d4a477688d65553036d6e49e2467ee95a78aa56c2382f81bdcf67efbbb18f5762feb66c234c80f4f712600b5a40a33feacbd83;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h142ae336706b831c5fe8761e73dd1d6bfa637dde8177615aa920c3257eac9f90eaa6d277cdeac2bb7c42771f7bf5b8f21c21e70c849a116af132b32896433e0bc149a8c7e47d2b53bfb3eaac3361697317506e683f6b3160805a8a2faca4e4ba5a81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8f116163aa3ea29e21965552b6d6541761cf235b075ff8388986d99ab298e936b25f02270212a7e54cf76abb030ee177919b33880bbcc7b99a89afe27e92e4a504b1c0ea94d33f8d949ac991c7d42b267103c0796d86e54d4ab347d813d19d8201;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf608654788ebac9fc5bb7827d20e331af24f292db3167764e7a262589f8542ba2e5ebcbc6989a9ab642696f3ec0b2dd9c95c0d97c427a25d792b8a889d047fb29f3d3d083c3be696767f413a70c61fa95cf27a10c3a102fa68b34e4953c8ed2e6317;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddb08fc4efac1f05bea1a4adabc41dd96f9ecfa3e406ca74951cbba6f57a0041028da0457d8c185e4ab2694e15cb37fa48112c4f66b6e3d2c2f572903cf5e045ad2b00d051acab291d15b4cd27d2474644a05ce88e11a8f3b12fc3009156c6fcf2de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee33c6ded6eb437c2b79701054b8686c59f3c01a1cbb5abc5268d69e6e3a8c22ea5cabed062b850a35f92117ae509b093220b6754ef61bee3f729d91fe8d9b7323a226687ba997dcbcdce688c12b7e5e2f1e901b2a21ee4e6d4a641f31f098b49007;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecc98bd17faec4a6a70d4baad9aa72c0e0de3fcce965c9c5527bb5e5f4c5d9812873a42f6fcc5f85dd5800486dc38b9b5de53fecef7afde2e1deffc70536261507f8ba2382c0811225af8e0c2eaff5c1af3ba53757e2cf9df130d35c0ef2bc00ae95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h465ccef0017cac11a560f74097362d497fa75622898380e570b69a95975e9a94f7b847eb769a0fd148436eec547d93e8bb9314ebe2d92f9735bffe8ad9d3ee3a5f0b486aefb353ee6d676fbb3c785415a443ed4bc0e2aaaf15e6b571e46bfe2439fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h341c10b01cf9ceaa6f8a2c5f7d3013bfe847e047f54a61b3009cba5503cfb2f1a77ef5401047fe56cac657b2b691361a8ebafbf6b0edb2b3c9ec396545863369d110695a33943c346d7e62e5486f8064001e69e4ee15d64c2177a213d18de1fa2579;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcff1406ef888b3c72992363921f2ec10020024a87f0771772c2436ad6bd6fb729c866b16141fc6ca70fd47d4c1da5714303bbce9bb78a6038351933ee2f2e7eb5cc5f5bcdde18a0c0fe042cdcaed4e58f2cf35fc9293344eb63dbd4769b56807b9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6fc0303b003cd5d02e0286a0a44eff2eabb29492b1f76fced9c716efcb014dc4e325ad1eca954dd5bdf773a3f8f9ed5c9be61924ca08ca7438a642401710cc4f6fdd403586dd4fd19963ecb9d4db08c7734740579a0737e40ed9864187ace947877;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5834fc442201a26037e01d8b34721cbbc061e8af174d0dac927d048e7b2773a5e45be6e8cf8e299a046c8c576c14740b7edc37a5cb27fc9d83495f5b9d78615f814fac6ebfbdb51971049f40756957208f7c46b9a3db88f14f86e2f59547524dcec3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebb75c5ee4c9dc70ab7572a80731e3e0dcc22f081eaaeedf1b6bd63b5a349e99efc533766b173c08e070b5b2b72ed6c1ae3cc8a4db840c7c87353cc65cc8c0dd195005ef9ffa811f72785f96281f1c83bc9da3296d03a18b0975c10589d814067b1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8967ae0b54ad6aee13fc5e1b54c15e16aaf297fdbd692a8497621bccb30b22b41f328aa986e00fbeb3dacb2be9c473478a158a9abbd8341ad5ac6c9c0efc1edbf472dd56b18c6b05f670693208ad33afe7ff0bca8e9a68a8fd5772ef9e69fd767c41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66c8583382ef5f76b819b4bfe050b0c192c5bad7cf36ac19dc4d4f99505f8473ca898203270605a199d8660fc5709eb0e243064d5a352d835afe0457105ace6c75f413395bc56e60ec97b11f239a1ddc71d27b9a377b0281c169f1aa6156b27818f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a932dba29d3ac31274f275071feb2e694da599b4bc372b5ccbe804b3835350bcd33e7268854ff0026556bd5fd6ab95198d38c6467231bd28bfca955054c723e00f4d493c3c04e7b22b01a6ad312039c25ca5e0360b3de2a689d4dd63d100947c84a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8daf23a704f3aa315203d452f925133ffbd1fb7b9f3b7609bd827a164a5bed9a41e155be775fba0beadb9533dd2b40aa8b4c1196eb58d1db917dd3dc2a47572ad7c48c21bf647b2c982ae46b7d8efd2d86e2ac8db0aed87cc92e1f42c1d94ee8b055;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h867d07cdc31e219f4bff9e310b12c839947a61200e47c8503e84349cb83aee0aa5188ca39f1b56f818dd50d114c2e159c783807787fc0920cbcac4bb76af416fcb0f01c21ac2dbcc4f08adddb9f05626eac812484e940aae8effe5f83755ddd49b7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h649ca76202675f84b7be2fc1d072678a98084e5cd307915abd1a53a1e24b0da5dc35ec4f20ccc4c3d6f016ec7b46c74693cb02d39928eaa588ac3a0707f78aaf9b8c5fa933433b4d78aa2b47312e78d38f0c1f9ab4b38560bdbbd5f5c6cb0723e92b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6273c5fc6acdba86e264236428fc75b30cc86397c0ea58c0a10558bb905182cf1f1a7546c75c39b4f63fac9a6ae86ba8238b67d102cba498b24755b484f1b79dcbb38262b6033c6bf2e37fd83abde7f39b21a8b69e6c7f85f5cc8971fc03ebec777;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf430dddc20160fb9cb7f774c89bd613b9f097057c5869f83a0adc4bd6d07537f7419dd4d0da71446f119ee984703a7687a9c455c40c8e041dbc934fcf43f8ca6bdbcd98291617c4f16e5da8be18c57ea6aa3a35fb1bb41452419b179455983a89981;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37ce391b77b3ad7d935b3c8df06e5395569e2f0daad16a31382f21fa01e8c80c7d94f0c52249faf8dcff542be13bf18bef90f9b2b67fd008d476a79ab581ab9f81cce75d9dd9c8c5b6d995f6274c53dcc97b9a3f34aabb92b7575928a847859d5cb5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9875d7c88e07afbf4f3ae21796e58b1d750bae873de413ab2e2f3eab9a8e256f138b71d75fc29e1746ebd0a6e8afb11a73fb73d64252ce646a7bf0c3f98d41b138844a2d72f417448a5d058c04c3052b114bc23753cc8cda18155d2bd4f3855ea8ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bbf4054d1c14b059eb8ea378b1cf3a61a1b24054c658cc7bb63397c2953e2ac6f5f12073781d95327ed67b332f2287a63d43d402c88fc0209ae4c36aa7879723063805ee66203fb2675d6d78095520a41eca3bf382b06708d2c1cc277342f6f2df0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72f6a2eda25044d6fbbb775a7d0bcf9197038ddb09760764ea04eb15ef62838b11617fb03be2c79bf6e78b27cb2a46b4eaa23c6bfa6da0c7c4b0c978c81c7a5e6cf8f43cca0103852f797085427039ea113b0b6f03b64ff1d61cf75ef56e1e0fcc55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he236e52e9261b00c3cdcd178a17f90d80717a6ec453ac13cded644e1b57e778d32b7a8310fec9448170f29a53addf79ad26df2c99d82e3eee0123cd9e474fe6534d7b076673cee1c3e4cc601913220acf89da0a80439d4bfb5bcc37cda7e1a0b0fa4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b4cddb31b7f2b7819a1ee1a3b4e1e99487214ed4b89f877e464975bf3a9d573b7607c7e5d5aed99c60e1a6281569bdbe16fea5cd6b500b25ebccf7dd3b6474b424d52afc8cc08cb3adb1232e6a5be6a5b27265190f986526875e5e088d450eb6eda;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e34d5f510d49b7e9d7368d85ed75c56ce38dc9985bec4f4cec4d3842a6a8d4020af16d0ef1080da82685df0959418cbb398793e62c944b61f4594c0e29f912bd493f4c50d40ee753e3194cf6b04358a60dc0ea135ce937fda93b623eeb0b6ec2dc9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b6c1ebd74b1a14b26cca7f723a688e9be1ea55188e5d6719ef4003671618cb65bc33dcfa36f8fa47565bcc06c193a5ccbb685eb8781a9c70d5332d4971eaa0fa38b50a7370cf1e21e84926050e2eab905d3e596f018921603e3ced8e59fe0b82ff7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31ce849217fda373d33b443cfe6791bf51f60763d8d7fbe0b0e5b543424e04a3e015fb1a10428eb748ecc8fface09d67791a3197712ca813f5d983b0e2f7ca59608468bd7b76c1ccdd9a5df9b6d991667c380d9a7c9dd7ea6ccc1d690124ffd9c3cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb990cc26e2dcfd2fe108078c401d8bc8dcee958e32ea51b4f5032567d3378dc1e66ca741f3e3124980d4bf6e7c320b5771049ccc718ab9de8f936d5a0e8ecfc6327bc2e4738b2aac42b7dd20efcb082fe2a5ee4cccf883b2262a330c7aa7158209e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb91fecb0ee1056361db0500566511ae27246203522816040a4e831a9d853f6185df27753b6ca5881dc9fc4844edc90a5b06d55f8eb531dc68c51f8315039cb691754b959dbc7e05bcfe4b7c6af8e873cb0dd55a63c92467060842ae765dd84245a1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89bf4fd774eadfee6b1da9b63177e91eab65814f4d917637c1ca187f9336be69c130d382ec087ab7add9a34b68234fdb0b2f37eb1c14a8599855602559f720eeecd4c6fe05af143fad798e00169bb1ca0d7a941b665e8c6a401164af95fccd867c75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0e7196db7e1e492f8706ea4021e7436893e56c065e84c2d24ca76d8492896c420a592c66a63f56bc7742aa30a28238caa61cf98403022a059133b339c80194386f1256baad3efec861f820b73e3eef1e59cc0c75253a07cbcd88714205ac57b7034;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce71c672b997e7fef1ef64e5157f4e23adf84d7f3aa9a60530721d756a1efd96b0bf0703907393e00844957045da0f215dfa2adb7f39e71497e81fa7b76dea725ca97ca561615d81b2f11d3cad05f84ca577ee40a9f8e63276cb6ccb111c01bbebe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76f72fec42751d49aba47421f47532f4f96f7d2e348bc11eca91b046e943ad239f1c90cb1d8fbe14161da9e4b94e1f8f29dd99ae625bc2125042814688f24a8f5e98b3faec1bd5518dd4277d23a7ac4e326ed31975ad072381c67102dc6ce0108e09;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b6f8f6c312c9e17b6dbd015c8c30e24e8b203bc37d83ef3099a2cb2135eb69e7f30a950176edd495b9ba90648e0250b24389df206de746a8edec9835ff7945eee8454a17c81f7e900c49120895f97b67f7a3672b46cd938fa5576cc1d73fe53ee15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9f0f8eef3bf5b5d5a8d0d9c3128cfed2ba663acb87a2f3f5709794babec2b217f1992f38275a7a44e09d5e9c782f6a870fce929a09cfd92437e7f0bfd9e24623a26604a6c4ade6ce4c1ded3cad2c1f21a19cb467d84fd3b1c74fa7de8b4079e3012;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had3b97755a61203863398624bdf85ea2ce75f1f56b3e45b572b748f57904c97bcca430537a0ec5f3eb3f8e497bf6447c7195c0d9deaa742a08e787f2ff97f022a13df94990ac7c42413082a87335d2569f4b30131597b4fa4cd32a12119ce631be72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e3a984cf4869e2b6a16cc87243eee411f3a2d9cd422a9e05e9c133d8106d353ff10ea726281c3462703f4262d915af6c0ed8c5b06caf30a0a449de5d7553253c39e56d0a921f2f9f1be854fa084d2cb9f76c1db481e688126f62f738952845ccb7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he42cb0f45b73dd89bbba1ffe37fd74df8336f94d7156083539f9c1275b718147da0b5d86c9ca1b8a3da729e9efd15f4d79c7ec750a467e0b85ec639d0760e8da79738b0692a267092dd99a8da31907e6ccaa8763bebcf8f4ac1d920f3793efe93da4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h385c367d773877aa4062b1ce76d9c17bc76e280ebb22cebb797c5c0ea499dbe4236ec564e14f9cc29478e65c7001dbce90cd04330b68005f3c297805e3571a6ef5b08c5b14436c694e8ec6c9ca93b0aabac2da3ea16e9a38c28592262ced62915b16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bbeb7de9cfacc619ecb48b742d677e75241093be17783036c9967af05050caa2c57d83525d56f956b77f0b893a2dd9849dd514f11da302d07b088cf9a16239b9d20d27bb2dc0a0f40844ce55951b3caffcb0dcb20d37952b7ab97b182be5200e6f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd55996f2ba48672e309f097e6947e11c7909ac9f3abc14237d5cbe998ede5070c86e5827095e580e5290e541da2c8744e3c026938c81465a7a14ade60ece00d5a92813775d2ce2758e0082791c3b03f3ce91ea69bcadf21e31fd4fb1d6273495fc73;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74446965c107fbcdaadf84ac1c2bf70d55c64cab06b6cb883914304ee75904f047c9c7ced6880b6bcada617cee0d9a0cc3a3502856674699a58c0c173228b52ab252c6437c70f42411a327d3376ad8c3a269ae43ee9146ff437b7f29263eaf7a07ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a47c95e273fdd05b67dda38aea81483b73b699466201322d7b0691df78f9ab126ce5c7572208e0f6c1b632e7c86c2ffb1fc1aa6455c09689c3cc7615e4df81d294f945029dc5b4337ecd8851d041154d870e3641a511d59321102babe4dbf78e7ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h171a079929323e685e57ed1066d47c4c68aa9928a1c4c3e24ffbca36ae0bc171d8d03e54832e71f70fa484ec500927b575afdcc2b7d11a5e41f7353ae10e75ca22c744ddbfe890bf387ac444b4c0ed621d9c043b1a32821ff55fca92011f903e8c92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he580bdf16de9136cf7dcca251f9a66a8a206006150026b79093050d8f27475ad2c6d6aaddfb4c72e214faf9a7cf348d6ed4b6d6fa700e6b214bb71aa81b0a6bdbc29e95e4a7fcfe83e89f6249532491feb40f52e1832a76e5aef4b0326899846c20e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9e45e7b5a83a061b19732958d30a7476f3770a634af3c4edd08940a5fb57e4613e96c091b1e557018670651552fe4662a574a691376fe4ad959483465e4fd025d7708186232f17278ecd59a1f2a2d3b2f3dcb017e37a1b27d8d3b8c2de731a67ce3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52b72916efaafe69f30a2205029340e65a815739136e91e33b531dfa73d54617d3e58fa141e3fd9e0016bb86ef3f2fbdca833b1ddab36a15334f81d420832f2f776c9595119303a2bfdf2c26cdfcd7fc29bc8c9690e99db6d048007c478e1f2c6fa6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36176b7ed325144ebe177588174fb7274c66d1359ed4cfbdb6a84d1a0f1d6fc0716596a4075ba2d4d7f01a28f54c77ebe24e16367c172230671b7531c28cbacd19f0028e9d76a20058eeaf8c2cdff8300dd563e92fb4031c79a4bad88f380ff32f64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bce9a03487513e2c59e65cdf02a40c3c0106cd1c67049fd99ac0440daedc3ff2309dc04f2b02263b64d224e68cf6ee549c7259a6db9fce500de4ac68577140be7fb8e70af78f0c4623353416aa3b928fbfe9ef65396a827bfbdedfa811226ae8a94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5a051b04439c288c3a24d44eb62ccf212fffe65ada3386ebdae44663fc14b42d3dca5defc7ebd08fac7d5d543603f2fd86833d51862e46faf903347286076ffc71cd1cc27e543f141350eb8bf04f57778b3bfa674fac5d2e32a39569fc9911a90a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6eccd8d91a988f077e2978de35dfe89ccba3aacd41b0edf062fbc859d7615b883d20c59ad0e100fec60382902a8332fcc2d8c6ee105e3430419a82e3553f05ed0c56656746f9038baebd783a17387bf610dfb211836684d7d11e48058b9beac206cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65313279d46f0b86688bf1d711d8a097a1491aca01793d4c3899d6f08017af8d361d5c8d9b939d8d8068518ca63ff404d71116967bd4837f9f7229bf5c745994d59487f7c7d79cef390ea0824a9e95c828eb5b11d8fb361ea71327e27e32624873b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32921575071dc7d1edd9f2a0065f6472062ce96190290920609978af17978372e26ada2eda6bc9ab12ada556b7e191163d2b23cce6c2d48d92920117f23a1694dbaf16c8f193f8e28f0bedf3bfefeb8fa41063ed3585936bacda0f495c03c6128ed5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57adab2d381a6551908114a4d190035d4123bbc62363e4475bebea525e9d978dc68fc70f7a3de9bc325cda436e8cf5179318a8392c0484168a068eb47772e5ccaef6d18e820247f922fbbab513e5b73ba473dbf548dcbe5110067ed37be8bfd7d343;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2461ad8af5c891672badf626bacedf333ba773001423b320bc86bb1d2267c856c209a3e687d550bf8099367a2f79ef720c12ac8cd4609817bb06a9fd6a9d477cff7121f9c464c8a0cac32e0a9fb0ab1935f7a5505aac5d34e8b21de99944461a36b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h409c0c502e8f2b624294a880b1392b9c528c12708160f7b581ef07b249157367a0125607c14ad74ca40bc5fde22e741e8b3a81f79b69b065a749eec87320e24f002e68a066d7d55653e0841617aab446cba66e3ca54444102b015078fcda0e4beb62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e3f0ce0198c0e78a3b726c2682d070ce32f6ac91aab8c2b5b4d3b859da92e902071a4d53d80c1a515851d204835f505e1dc54560c1edcda87d302f5f8f9d84c4c5f1a15fcbb39dd9fbab6cbe075941a7c858c30dc9ad389cd65641709a8273f1cb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2c5c15ce083af5be22eee1d64bf7277037ef6849ac4ac95f36543d9e5237c076e838f045c2ce05e771cccc3f54f81d9c091eb9e2f22592584843edc3bac94d4731deff5d5262924e46f4194e65717913acfd4757b6ae34183f0f145c492f63eea2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he62c7c0df60359e92f62c2439f3609d37eaae97c2eb8ad5aaa792c399998ae74bbe9a392a2c9ac57bde9cba014368a535daac156c459d202f354f77a38211b1de356e21824f2cee0eafd45bfbbe186b1e718825f7e33f80c34d949e78bd299cb30a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ed96774aa610235e9682e33a86c8662cbafa6b0e0dc679f3e7cbfa7e6cd83995be2f1b73df3741a50e0d45cda179edf3ed8643e06d7f01337dff2308de768160d51dea8e4d13cf2f993c7c223cd137640fbfe6517502ae90399a3005301b78e65f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9fe85485d1216d32a9255b9a44c6f362f6167ae332b20d57e5ff70d5dd563194d10bac18b3b44840583350405aceab071f1d9bf97451069f6399d8b4fd0e71a55eb2bc310bc286730de8d06dedeeaa41d0897c0dcda056b84ee339ef47791b88e89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc748aa2b5b1630071a22f5f594eafd84c8675610be9d54def72fb59e897c05e8e6ddac5b70c25dd4158624bea8e5dda46b592050617957105af89faab25c3e9121660c530f7090a1262656428a20eedfa331a36028ef9985dc9828963c7ee7f9005;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dbe11f9d5332fb3eeda03c859c7347596909bf498669a4365f9e6d3e66abeb868c005097d1071af11ca2878fc9b13c3dc18913bc80d109824de6ff39921e89dae34f071395a588fb96b854dcd774ec81d889594e3c358392ba8067a0b717f594f6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h368109425a717da4c71b7585ab6deb0b916aedd30f5fb25c3794d9cbecab48af54978f0aa64a874d11cba60a2a14b5508b28d6033540876a42170ee0fe4652b77466b91ada8f008695ac747c9a3d10edba2b5efd952879c339c174c1833ff75140fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h169fbffba40897fbf064a6a512f41f1d1778116661812537a950d1e123aaf5d61092e3f26666fb4d4f205081b6cca095baab650d640bb79e3f291ac6014b4b1ea1a648925b0e6844ac20dd8420da68f0416c33e3ada138c55067c6858e28c7a2e8f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haef7bf8d83f0a228b33f5ed99d9df15d2407fc8fa0a37120c642758d63b0aec0b027c8187d8ddd47233a20b52fc39775f304e58471f56bf230e925ae811123310f0e8a78599baa63230a358b506e20a4534461a9486f94769394f3f56ca8f573970d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bd2941afeebdf37d62b9861b789d07413e9e015f158b4adec1f95f0146c0b16318bf698f151f4d425e72f92b59015c7cf1812a106a1836b526980aaa176ba87ec7e9e95f424e71864763dbf1ce1a55cad672d63a36afd7244098834fcca68535a16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6122659cd1f6ca9c92340ab1e10e4f49b1a7e91a4cc079463d143abd2b5e360bc84e91a14fd0c322f4e83dd57fb07905000dbf65fc7c02e31c1347ab8020db71b287622dc452e3d0ed5af6d41c60f7e812bae23fccc9ff1f2d15e06b38bb4a47da43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha969b0f5ce7e23c38a920c02e7b749f161614356c614a4502ddd91e018e493c028c65d1eba097258b24166ed8a26381ed31744992d956c484b0bf4cf7c97a71942f2640369fc6e169aded1567b00a9b6cf07f1ad15224d1dbea7ca132f1df430fb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb473a3f66580ac3057e3b436fbd158d2a7e9e2d176e1bac75c71adafd899e12bcc418258dddaee91ff2bb903478e0f5e2f0ffd5bdb747c8ad431b5fc6d240be770f4e7894a066401433a1953eb318bf0e36ab3ab8aa8680a2a94b1682e81cfa89327;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf342e0534c790f3ac277b69b81b9497bf8d3e052eea1d42b6394a08b42451e7624df8c00923286ddbcd71341170091530af2aefc89e881f4aae6c877e7de7c2501fa8144e719e2682a3d4d1c1165b33300b152fe72fdd7054ec13d3659e66348d935;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ff818a4caf140ccf0999a5272e52cbbb347829da36d0a2b3697511969024d23c9a4543ba55f8c310b2b4982471a294bfa208ade9f470d4e56f25c856eafe8c1b6f697e1bbcb6fde9e271a393d128e938fc0a05e7f7b4648c6a4015e374b12396494;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb359a95fd43befbdab50ceac76e2c353983c1f9870d444cdce2edb0f91fab4ce1959727df0500323881e1bae543c9a2bf7daa47bf6f61b2878e8a95e2053c4228a0010975025eccaaedd2c03a57e991101bc7663a79d33134628c6714d053a8c1a22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e48a3ed66d3c306196a8ef134d93d29a248d20c9e2bbab8f0c69c08777a9d9b44daef0903432475ce9241212701f9a65f50278e34ba17fd98d79ff686890352e40859472a0cf3af5c716cd62b9b55916e9cb48b53e9de285406eff8ef6e5de25fd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbcde9fdcf2100af4dd6701b7f93da6455067d9ae86fe0369061ca3a209d686d5972cf0b47fd288391c90921bfd28bedcd3d5acb0c9225d869deb57ab9fd3de5c6bbe40543e776fde65409782bfdc387e44d75975dc68256aa51d353d363e9ddfec3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cfbb5c51b674ff96a9caf16c9547a7c231190217aa995f2164857ad9d450d85672911ad1ab510bdecfc2c337a966f40550e088bac39b91d0c29478718f7f78c90f386e972ab76ed7846b3bad08cdea0bc9d877470b2b83c39f7de60e5ddab1d8ba8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba97c9d5025cf7beda9d64b2c0ed6ea60ded97c3abfe92995a2793b5945280b9cb94f0542b78e422c5141c08f0a7895af6b634206a7cfad51775e69305c68b913d9e6825364a9ceab6b300864bd261d94a44f06508357ea32592a131dec882f376e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1c6b9d00bcaf4e50ae1ce45b3e55d731bf69bf1278d331a80a48395c24e2f0c4af5b9c2fdde570c41c12abb4171480ff81ffa3f2ccd412d20522547e736a97017c52b36fb08ea56c324414d35f0fd33a2056c8149e5a485eb9e09a32e983e5df1c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0402dfaa853c48d55b7a1204df7ca4de5d29163e3541c0a25129ff1ba4c4ec4efdd6f7724870b1d3d84a46cd931703453f0528e1256b2f56613fd2e5e25e44f6f2b01233e197edbcf3607d0a83fbfb8b43cbd138d37f63b5d40c147c6b9ec89cd84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec49b237152a58eff8f78144520d4e77cc9c4b99a6daee744aa399ed50f2b414d5e293e2edbce4a5c7114a2bb8190ccadc66343551336b3649b0c3a3a4c39d44428307a49fb63b84e399ce73de9be7ef9dc7ff76c126db40d2b0d9629fc9bf9972c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcec01e81454904ca22f599114f5b3a1adfb0246184c098af5560c50f0022f58d28aa02442e707279c4f568b4795a3f48089e8292fdcdf2bf74003c3ad8c58907fe76e1d139a651b9efd8e349e45266df86e0b5a55a7d8cfcd917046424ba6768a7c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc078e69e611dc07c7efefcd5b7154b21a1b6219993486f7c264bf52a6634336d0b92b5f635285cfe4c15cae4cfd21ee5a29e1a79856a7d9f5f6ffc4932eeb023793f6a47dfadac8b12a41d3d037f8e1312a1011e7c5506246db655c4b1f9cf91964f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafd132d0afe84140cc51400c361179225842bcc991540334d0edb0d428ae21c5e43105ee04a20c383091f744e63efb9cfab4dbcbbeb204b4b0438d08531e1acd43e8153baca7e4fb5a1bd7d7df27080a49d43d723631c9cb32cb2c10c40c46fd9a5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ef0951dfc63fd2b7059f53f4cc79062a2c83cc31c1aa708c8dbbdc338eb6b2d4fab3dd8e2b27164456efce1d08c7d3ff87083db47232320f16e082328af525a8b465ef255ef301ac6057adf2fa300deff471a37bfce3f4a4d4b2a9db53c8a69e63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e52ec5a7681a2f4825c4c956546155982b56ac0ef8cc5ac09a6e5f562b24a482652ff666817ddbf1b6374a62304a5f5166ceebe649feaafb6fbcce219c2116c2f8d0a9257f684c3c98a4f5e66795d1a0348e6cc9d1c056a3df22749e6906747a86a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h429ecca2b4286ac0ef417befd47ac17c4dc5bd842a234c01db575cde4c19a9e7fc15bdcb1c6a9ac0bea7b5334c8a1cf69707aff1282b53cfc01bbd497b67b9205fbe892c4037cbadcc973789c48af92c200fa01979484f608b3476a4ec48075f9492;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd73edb3671b7cfd48274317538678b8a962a0e43aa1c38044a0001ea657be50fc014ddfcfe28c51a9df64a40d82da1631f1e81561304cae3ee1ada1e9957d0578b071df4dbbe983f504402b5029889880fd92b5e9f88877f458864356f44eb8fb23e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e99dfdc77fa825ee6eb0380130ac9008566a9824a67f41741219acdf3d156c2685fc276f5f9eb0a30a899fa4fe8c3aabaab1f32639c2cdfa0e52d18bf183d8d12382511d9e2a663dedbae57d92dc1cc6e5c9b370d3c332fbd54990f904191b1ddfd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6371eea9cd967a0d8c297ee818f75d361225623bc66232b08543b89f1e43c1b106c626cfb4ecb56a4796dfe2c52067b467dcdcc93eea3c5e1ab22dc94aa5499b9bc11b7b0f8d45d01d3937f406fbd965d3c37fa5f7452d4927b6088eea108de1d13c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d97543bba28956151e81ebaf8d740b291c271d398752bc4f89ecb7e26ed4b612a60a9b2a509ae59be81071a4818cdf345dc36bac0db0ba89d1d41321f703d93cc441bcf1fca18bc3a0d722993f650881d47b6fc2bb8e2ad202e3d5c6463b09f15ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcea1d8c57bb98036d2ed3f08a02050addbebdea01bd609a86e88cd306a3575cb8080e2bd070732f81fef917db9a5830afbc8988019c023cecff0629a715580c760e70cd7ddff46deed403b4698a72be1af017f959442d2092292f84f29613e47bde;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f4e9c70f3bc40a607d38f0f14c9d8ccf9d62fd36c5d569c6530e3d0e0d55a4e217040f167f61d3750eab726db25f944bd1923cf4ffb6703e1111dc582bf1ac1b9cbfecc14b8cc80211656fb409255b45c445e480aa532233f9c117a2ffad5d0f6bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c58d95c864e82a0f090610f8919edf83d7c7c07051fad0149f7ca6b8c02079bb85e9c399a22073251bc032bf8b6ef37080e3ccf053f7fe50f1c2f1ec93e28b125f908fb693c01ac5f856a5124a3ac9a8731879753890f05b275b0836debb7c87a1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d3508035945189ce7fb4ec7e1eca1e4c07ddc5e86385d95281bd89e1b48a78b83f3ef988bc77e68c2b2fd9c442dfc8630a7f46a79ae675ffb4a5c6e3ace7e82a414dd433199ae87da6aa5786ff51ea120e2c2f8b403c94b11e2136d368affd2283;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8ac0f6822fe5ad2d8ec9e618592d1eb14512b5f76d461c359dcde8245d403e32fe3b98c63867ed71ebe28eb1cf99131532a5a281bca98ce47ba61e333a703506f17d5e02e115ec4868e44085c531a70dc9014d8d2868c0c69d3a729b33e4edbecc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda9bc84fb8a406de0ea9e175a6581af20bd75f36057fa0a9364d8980c3661bdba3b429b88661581a79c8d4f2a509c4e53131bf55d4ba5a5e4159887b2d834264e25fcaba032dff302d7a3b174c4a46501bc8fc98a7d49d5cb78ec10774c908375788;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5f2cb701637abbcac48a1ad01cc2e91b77a07af93df39fd2a707e4c015a918342669d12314a658c065e54a241c1dff4ca8ba33752830afdee3e5f2373c652c071670d1fd39523d616b124581cc1a3b69259231a77788171e7ca33783dd0291fcca7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bfdd1ea30b0802b312f197a612aea9075038b9836d718b3b5f048c934a63a29f7ae0ff350669eea5716df349ce6aaa6b76de7426f22aec22f98dde5a08860dfaa05fc77448601ff5b44f5415ab05d9dd930d8e09384c0d7d761febba93bc3d17bf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd860847013d40b404b71ea37c4ab3847688dc5081afdf8b43c364198b2d7aca838d0ea1e6c85389be69ae3c7469d6a445d6cbfbd912c9ffa1f528bf02934452c01a364f4ab444e824eb68ac796fe9868d3462f85dc3051ef1c11fde7be5cd4f6d890;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4524454f20b5936addd71e740d63ab5a3803d77d39488849e0450b1db09a65ec1efca850dc3ab90997b4c459af80bb6718edd8d3f2c6694826ca336d3ddb145c5a6c8d64c3d516a0f53d4e09da641ca13eb41605a396e1e988b137c8c743d7437907;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94df41b336e03232c4094521af63702e4f82f4fc9f00f5e7bda6ea576ca4ea56e94801a6a13425aee1104bba2e65584baf1aad04ee1217737ffffe8d3cb7db73a099838a11f2e8451110c444a0302de1a3075293a46295514d1144b529d3913fb676;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2312183d00452d0f8f6376f93fd88f1eb8504049cd6d67f5c1e745ca86c5c4ecb6006b655469128be3c99a0aac00bef4002dcd1d222aba6044b981f7a9acca5478d498244427ada7c33674ca4ec5f8dd0fa38213c5aa062854c2c75b6e9b001363fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef820b358821205cb726ecef11c209b9ab0203bf0662a44128f9188194a8209c82c07f4606c531d62cbf4ba842d2582ae65a40759fd76f4b7e5abdf9bb2f42ac399d9f26dc2929f0054d03d3c3bfa036ab06b440796949cc2c40ce54fb6e76b8846b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fa73b88f9dac91080d0a648a79e1ddbf101b76270a07c591d8e58dcbbad3befc5563a0bd86008049621da6b6e687c3d05eb60092987d33d305937e62b6ff4271c48a0615141216135119c70fe95c1dc70b8b2e1e7a36b3f184dad0a711817bd1301;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf2f1a073bb0d90044098995cb0025731fdb51a441a44f412c3329ff49627425b585015eef0c095ade4b566eee3ab22af9e215e75702a52a2c5fe3781234aa49c6e1becd21458190218bd07db14cadda80eb2d117c4d5468fad1eabd71889aad4f06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf349e1710c281bbcd1b478d55863daa4bedb31750976f508bdd58b88f81d82033a7ceafe580c888e5f17db84e633cf06b2c0a83d8dd1f24238bf6c56e80dcaba95a148a0158312a3d532e6c5b4c8663883fbf4d7924fa4760de57165d8e0e9a1e0a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b9a75730cbf395196e17262b0553c4e6f6bd497e944e7bffd6d3bbc62ff352a7dbbb454c06e6b081af62fe28335f6f45f6e4d4d2323721b17c2808ffec73b678247bbffd5d111701608b97a2b4414f3cf9a49b2df98af36c87f637cc46d3cff7748;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1073626bf3bb02aca0d463a0882c68713b480b58f15b35c5dba741ab92b743bb53a8a789e4ba88ae48e767aa0ae613d812f66fd3bbb0fa0826a6534d94385143060115ba277ff7f91c4efcc2174ac51b930414371c716b0d567626b6026717a510d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5aeae3da3cc11007b566d5db5491aaacf0de5f6eb278931b7ebf5da8f6b79d00fcc182384dbda1483c5d3feed7d7d6c46baa385e323706c235109e040341ceac35f4aa7a1cccc392051be3ca78926af5f16089d04693e5f5d21e33cd7c753176dad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h275901e265f6b24f4a2570c901833e7480c895573e1b3296417dc388eabf2d7528a736c24161ac1a6253a4917a11f1fe970a934e8b877e0ab8862f4bd6f00a9a0989994a00868ee63c6ffb28ff18a2ab91f13c423e875cd9076fb3bcbba350afaa5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec56a05fddd424b42ce734481873de97296f5e1456e79191df6c3ae2f2012556e7baad7e017b7b0afec4740246c6bcc5981dbbc795f62a4a1977a9b416ed45e6e9f30ef4be69fa1c49630a42321c71a2f9f33cfe753e78a406100c1f15ec1b54e30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haed80400045028862f508cb5dcd08a71bc4aa451695d3d027d230e6b4f4076ba82d66f5f55aa375876ae96e101c18e833be7b2ebc5968d955770964cd905ef2138537c1c80581f528d9083163b5b8466bf6429b45cccf5555f732efd901e6cf2a046;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25fce93d438f46342633167832506d1baf4a9b3747c1eaa79b0f15b194ce4fd51766b3d54a6d53bef5359a284c19229e1ddeacb6e560e172a0b1e5e5292b6cd515f29dace8e3712486ec33125ab3bfd81f1abded20329f082fe9b3fb3e9b6696ad4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6287657e047137101ae14d39471a324639a3bc0e0df0230849808c9e4388ef24bd2d8aa073634d0476970d435f8fc990efe207b1c64dd2956c58db278e0156d60847b40b2e211f8d7665683d0d809d9bca1e87e681e7f37a5e94143f69c6251e9ce8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb0beb1acf287dc021b017018d2b21b18fa4122a832d62a2e61084162be25e96b67ddc26b76e21f48c554c4de2563c30f6343594b586c1499dfcaf4229bbe24bef5d1155552fb51c5435ee09328259e5c7cf0bbb34d083f46346a50db381cf63589a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30b26490f759b0ab7e39a0c5dbd1dcfdbc600e4d440e4c4b52dabc949ae1a69c160bc479c867ba02cb7024619d00d9e4eadc7ac036c87127f7c64b7327580abe17726d36594ea1baeed6df79702d575878b640485e8168fd9ee1b94e8e5dd80fe89a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc874e9de0c5c08a14a0a5927872a75c9a845cf5be289dc12d7e04a5585838c6d78ae5b3841539469dedab78b1c2c94fb53185ecf1c47a8759e04c1164b4b2def2efc54139c5269384bf2cf3ec85001e148b86663b2cbc75c5782921bbc755f47617;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h640bd7cb49793dfd6a0f9cf632522502e1014d9935cf652459563b8f2d94321ccc1d32ecb76061f4696d2eebcaa317bf1f021563f820b2f3853c7c26c5a819f105783c3b2e4abc8ff7f2094fbfe8ab4f733468155a4821167904d873741681fb4943;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19dfc1adceb02fe802233777aa198b107b065cb8e27ba42b3462cf3b6de02257ed73695031a8f525bd35b6ec3cb59cae5976361082cb1ba4a43dff8bbe07f6ec7c727be80f06bf21c1b4f695dac106da41d364e2dbe6b07369a06254c723f918044d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfe268d34fbf5b871e7d01e6f113bed5df97f34c28991f7387a668cfaa14692ac500a8218ecd562541776a8a56211cb7e4556c67c59e4db9fc9ceafec13a010b403c88add7ee2ab0b90dd55e9dd59d190fb939826387c94c4c823d4821d378884c54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf3899bb177374aafb773e385366b4894bea7bd3e17e2f89d5f84ed37f8317132026f77c7041b2cc9ec1ed81c86489c9fb8f06405abfc6f0870bfa8062be7405f86ea8851eee62dc07c46dfa9f2adf6cff9cc15c04c8a78ccae0320031d0fd9de4f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h465322d717cb831d22c5fa9d23573eb108a129958f39b2cd1bf34ccd9c2b2692d1571e8b4ab4cb2051986ce90b49de2aa3497e7a010d1e438e7f50bcd7ae7bcd80746881cdea74c47a42550e97cf69e66f926038e031f8f00772f64fe037607a63e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb2a27cd47c7e21fb4cd42758ae31317c4fdc47605bedf11254cf3c480cae05401566cf74e2b36f58ea3660b4dc699b8b00c9dcf92519c0a64618e26873956d158b8977c3fdef734430de1bf23ae28be12efce9042e39e45771242a0e5d1352931b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6afacd7381325110b7f40fbf5b8953a0589a7dc810b591a466106bf78cb8e108f7814770cbe49471ec8ba1d633bf4b2b30e030329ed4f1a11ee1040fc31c03e197894045c85b5b2b09a90f777857a48b173bcc124e42c1c79f8fbf709c06b47f0a18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4f6ad23b44944c8cfffb48158ce63eec63fe2c5d95e69863d58078c661fd711163851008d372579feced5b4fa3d9971de3622f4c38fa926d4fe453332a2e923f01bb91835ec4ad12704e0055e26f005e262f73cbee5f658fcc6ea104d373fed40f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ea014101dcc604441dd2b6f39b14c796e12e4963f75ac3fd5eb0676bd8586d1ffdc6d9e9d7b13d08ec94586dd0231746bcec47589c333414a0a277d6b761aee4cfeb8dbe382e16566bd2c883879f1824e388fd3dd16e140c2b474823a18e305419f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12208c50871c8c6a0f0cd661055e4f2b6e801241b9981dd6c30a282275d6ded16b03f3cc793fbd7eae332e9ee41ed650f7df656a508d0d2e8c05aded39162a8a35f40574a8a79a02d9e8ee56e595dd355ba88473867b2093dd71c0b54a6a54ae00e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he04e1ed319537912c6872c24988663841622b8998b1966055544c246dab056f071eb0df4bc7d5b6ebc15d7b8fadd48b90648b3ed7f07ef071f310330e8cbd1773431c3ddac33807bcebcfe9f6b4175b45a3a24eb69c5da0ffe805b86dad258f2e81d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9909c173bbe28e74d7c3193b1613ecffa58cf3b5f804b67dc55baf244b2158bb123e38de8ee47b8720bc63f4ab8ae2b80aba82bcf54bd2e60b2aacbf611f7391077fe41a10de9d8959deb8a32924e1dc6d75645dd44795b6cd5744a04e10e625d21b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf9809d4bf32a9e539291f7cc5705826e0eace855c9f10abaa3a500374ff8db371cccd8d9d3ad93d1db4d9ead6667082ba02cfff1fb050a7f5452128fb15bec2d47ef7795bb2b62bc3a3d7c046ba2799da742e8dc990c9801c816d0bf66b030f2409;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6295ac793e45e782d01b0e1634542acbd7a268d17434804e654268dc89539aa6826573c31a5a3a310743bd8148e8d56354b2823c8a83739a33604d079913f8b96180ac7c74cd426ea1966f55b98b261f7da784894758a45ae3433d6da7e082622aa2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b5d0ebb24d06bdc41c8d17ab9f02bdca29fd66380c94b65f7b946422970ec56ce7c791c715c5a76ee050c170349ce8b158e00e0532eb709b37257c63bcdf23ab03263fbb4b460bc6d72d4f8a778f25553c1325aebf18077ddac6bceb533cbcb63e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf77605c94ad6e11b29845f96a44d21babb4af003bd6c84dbce1071ab6d21faf4277169003b29358fbd5960cf9553aea6d7164b1e0bcad75607ba3c4bbcd641ca2ff63fb2cec9798e492e364a6bb24bd6c0dc25336cffd5abeca6fc0c70f33ba739a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cc9fcc1a028a33385b768af1e25a22f83c6a452ae3ef22a75b4632ec348c5cd1f3aebec2530e7040dbae78ac8e2d531356260a3f8a136a743bdebe916e8be27c7828c24757ee36504a2c56cd0ae6fb871a0cafc945936db0d988c840ee7eede8684;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78d6bf6dd9cf6a2defe29792743eef79c5622e29c997675117156f6b6f205f353fcb123b974c566038c9a5f7b885a61015d6f4885233231af966000a500916735a965484ffd95c40616f7a44a95cf8b02fbaa1786fc5c8eb0f8261389ffe2cef4f5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42361696bb3d0589ceb1d1df653b7e3afb9132406a88b623ac9ce8baf368d6fb3585961fb3dc67939262c22d59a52c72662c452768d30656f3870c94b27487f41b89e2b1a6703d47c6cea1c6e5a94d0ac887678710d2e01e6ecb5a61f2b3bb44b8be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34dbcfe4bbca1b457f12d732a25827d887e290aca801733ffc6aee23594e0c25f62a06acfb5a483448d37344ff575a83a1dc45969d5f08d77e749b86737daf587cc9f3ac2ff1ccef2fc2d3241c746227bde5f2850b48f13479965c693633c5e081d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he58802c2f8aa8901aa988e427bf88f1c016b085083d3a1edcef336c1ddb0845856e21579605d2e8da78e02497ab227dd662f5e5c59b7e7546235097c6a338b3eec2c09c844e44528480023e0a66a9f929b61fe5cf1b2575265b59989d753d1a235ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24896f9576cfe807eea0bfac1095880e82c9797acee9f09f24703a02da7a1bfacd0cc585ca5f1d756e872a84ca214d89e7bfdde8a2f30e8d3a39d74cddb3cb0b959aae2ea3f30b27181472df0684803929f27dbc3080b405b2d7880be1fcb8978798;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d345ad46d0a20c791ecb9395b57d1cf0e80149b6848d9c0bace8131b43cb9e23f6f5de9cd73e9396179b4488b1c9f5c876782a885218867fd18c2a9ed06ac94a82b8d729058d9de8ec6813f1974249f7a47f29a9953477282615ac1d2e0f0ca511a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63294e6e1546919dbe4dd2262e103af347f14a70785d9f1a100d8f02b327099a3ad3e25a5309f7be8d78f946adeb1c24cae683347e08814de4ff9277e379d04753d98fdf5e89ee82d2b3e5ef24b952545bd6965842057ae82d3447a4d480a9416b25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61fa858c2068a9737ba3879cc1bfda38847c51635405ad1beb48dcbda9a5f46d9e3126e23ab415975e13a4eb36444664913c2dec2a3bc6db641a41809a15ecaaa9694336f21773ee929c1f64e15de09758c9c01c598838b1953480756882e6561c72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dfd8837b004f2316dfe5d74c5a73e78c7e7cb9b578bcf9674a20a2cd509f9d64bf29d689fde0eb9b1994fadb0eb5a36138443e896bd3886394396240e452d3f5fed1c67eff5638f4a7fa73cc7fa328ba2a537119e251bc491c87166853d980c4618;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880b5f3728b0a2de948803ec1422e75962b39941d05bb36b29e7904ab82c6eb3d7b129c6f555747aa139ba8270a0e0c349b9d02d8243d9ee138761690ff1dd99926c955bd1e54ad8ead3198a847a2936c9e6c9826bc3251bc0feebd05476ee73cd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb54b5b98d84432e31e2806c7fc50461fdff4ee90074e17587d3f0b1292dd0c68d5f3f012cfd15ba588ac5c4ab5908873af93d0742c3eee229c527b9e7807b61fcab71ef43fd719ffec6b25434c72ba58ae3b332ccbe0ada650c3a12484d442f48dd3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he36eda31dab3792adb50dc1d2ef99a1006b7d647ff0720de2c88d2dc1c384416f63f97255c81f372e181a02a11fb4ca02aafdeb31dbaf86311878786e5254bfd41afc4cd5c35e9c9bc51327d8bbcf3226575c43273a78331b0f4e0f2dcbf535975de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he207ae0a61beaf3e1dce5622c8190b331b46f9fc0e2751b9b9c5b8b9098d4e4aa0af2c9da09aa70668c32eb6123560dd969546f2346198634185e0c4ef5b726e9eeb6155183d29a9e93ebf4d7e9c2e36fdd8ab9cfc062f938a2e73321226320fba73;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e099d23e539baac46ac16ae92c6aeacdc974a4c8e7337b6983b33f4c6f3782a581d46a819f72bd5d24ac6a093fd5f444c64858129906cc14266301c999ac075f6d4206612d840aaff6f96e3099290bf42a6a62d0a82d853ca53b42fb1d081f3d9c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ae77ea6cd8cc94e3423258b50143946909b6c0a1e29dc3da2f44701de7f0215c0ecf2c1d3615c6f1cccb43eab9675bca0e4dd42cdcc4ccd88b21965433a1bcca1fc70c3df319e8eca815f05b83c479d9388fd8da0f9cdc701e52ffc914f4fdd2fb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a084829971f2bca4dbf34f569f82ec9fd98b4b654ed8099c9e630b5fe24b07c4e6635fc0106faa32b3ac4686797c1ced17a481cc5667794bc9c6dc224d4d39b60c63727540afc2abeb8ed39c7170d6b36845adbdd8c91ad2816a3f14e781233f3c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17235fb6c19f69f550ee845db386b85c7dcce96556bca88472192cad41c1bc5f8f209d9e50ce4cb53db13001b948c339df13f1ac69d64bf6587c2221470957a830874e8178b2d06b9f778802271443d6f1f5b71c728e934953e57a00aacc0846d1f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7fface2a1fc297686abbfabed83281f402e372d61869a04eca1aae8402b50f57514f0ecb45249bf2e94ec179ab5878968fced1e70da0d11084696a4f2595947679abba65cb3123e9374f0778474a48de711224628ae429e930af5a08f80fbf295e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13f0aed6026a411a5f8dfc7c25ff7286f53a579ff75bc49bb78c48a7f4856cd37424291a8414ec09132e9d61ecea0e6b22c31cc3825a746f709d727ed4f49b03c60dec4689309596f4989fd44d955074945dcdc94d9738df5554ca8b36b29eeaed2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd744f56c8ec019bf8785d4948c330202ba6e4908be34ee280bf5bff3b31b7d18bdedc9221052688d6fa22adc41e8ebe3001e3c9ca253867b3d67168a2d525bae9263387a72a4d0a4ecf7780cbd9d27c9354278395e4393918c809fca393042d9ee77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2408b93f3cf81d89ea9edf7f8c23452adbe491fc49433034322c53c96e7ce814d2b2609cacddd7246f0f54aa8bc03436db21eb551e0009f67ea80845c945a14e0c63da204c65bb0af4096b9a5cb2803a9a3a49b694954e46125b0e24d6f6f8066a58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab47379761ed4b7fbb8385e3024cf549c8229f5ccb8d01b67ba3feac6ef7d52b3fe28ea32fe5a0826180e9384359ac179fe686dc1ff7f75a9fbccc7ea995ea3163c5cafae993a7657741692441b59709a2fff4eeb62feefc74099665df77b718fd86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7ace5cccc2df9a5f4461420490c6ae4224dc76695ed90c4e634aa012171d9e26c5b2b8b959ee472687a2d16ba4dbabc829d85803d8ca47ba16d2a0c6f9aeada107f3f2178feab1105e8132d8d509b60bc2a72185f165a5114ef1545bb8766a5ff54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6afe1e17cc9c6cd1840da7c1de398d15c57f09a8d8d25aec7df92f4453d20c9c1ec49e2edd27a7eb054661a6007c5158f9cf5c28d3a431b0452648fd4e6044a4fcaeb78ba048d03f7354ce1fdab976468c57f4766f791cf1bf93921e4f47c6cf0f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56d1a173109ba69b600c7acb11d01f8f5d791d1fa39d55384f70900f1416c3f1519aa58e6f1b58a3de6d1cb2ec896d1d6d29e9078ad7d1ca76bd18ee2fbc563932a0d24a140301e65098fba8de69b59262e9ebd07ed86fd60e7030eb0cf5fb06fdb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88bb94d3fa83e1810a2cacc7da2712b8470927f6754c92edcc5ff1c5ed1dcd2be979728c834cf607777b1720aee704cda3d0daddc2f050d53ff5e019ce2fe53af991b2bcfe0f37e859d5dbad0ac7d587bf7da3634e93c0673f1c1975a3d4bdfc8af9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb116b39e15cdfa9fd03458a5d0fe10f35af23f808b7a6c695b804f300436ddd98243a1bd3cececcd6e4f1604237689d286845ed301fe725cf6b4e4216e3bf8c2f87032b3acaa1c31986c6187cd9531203422638fa1afe9bd348828dbb87117ea1a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h541573ae7b07fc8064950e372979fe239e213ed16475e9e88c6ba1b2ffe8ddefa49eb63cff2a607b9e60bcf7dadcb928e9224ba0a3e4e4b18bdf6bbcbc46d5b69e54abc9734728919a28bb4fb6fbf977267cfac4e64c706dfc41e7f92b3268448d32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42a35ee1c67656f1a47466e61c5001aeb03a5dba66dbc3ca99409f551e4f8c684a5ed1c37d09a709c1135e5a70c5f05f77ad5aa93e318cf123458770e8ddaa97495c0c3a29a041d0e1b0943540654825b36da358e9c424b4f171d608dedc7f4d93cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb08f36df015d1a59f19f287d4105e8bc45404b93729aea8f9f529ac3906775037e2e69fe98d70921c307006688e02885bb5cb86a8876ed14250ab5fe2f02efa389105f67ac40e550dc403f62f1fb8cff796199f811af0019337be7ca8626b3a1487;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87ad6bc7289472c2afc239c0db77e01ac164e6bc1acce87be06e5529dfaec8995c6b8c33046de036029fd0251f647dc38252fe30f789ced89090b3dedbc7112322a164f3fd2fc0aacdf7f9853e9d776dc726890ada9cd9f905e73ef73aea4241846f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58b16ce8b58325f3fcea779bf44c575937432448fc0c64cd69ac9bc60602245dd5d06a68cee36570b68294ab72c5520def68aa829b85d8393d9d7e0d4024718cc5cc7c57f9482218b0dd7faaf8618d4dc70e3d6ff5252cd4830dcf267efc75499694;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb1147a6b979ac6edd47994e549998a2c8c7b1275b5dcb56975a82eab112ad8a4ad54d85610332a7339a7e92d1f59417e8a7c3d0cac875c30dd02692f51dc4aaf969a3d5c631e8478f87adc6f18dccc526cf623749c5b03e66980bce0f7e971a410f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h793831d578f85f30319720f985b1dc9a6870c069b8f9d64813ab976c9c9ca09b978e30edf87774e9f8bf75f0cac2685c53a0877bae432212431b4740577252b54e5f760a5aaad219c9e3994c6b88f87ef4abdbf14f2a594a06a91f048b8bced01e7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbbf8d691920ff32c36f1cf494e72aff40d2e40ed747a4070ec6da3c78b56e1331c4db9b4f61158db5d8162c0b878d7565870853c927f5caed9ede7fd9c44a842a02c60831ea65df536f346e49dbcb28211dbefcd053bd761b9271a28847fc257813;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34f4e333bc534b4c0b25e7656e99a0b7010c3a86ae9bcbf835c433431f2f0b49053ab40eb37010550773055a8b4b89e11a5d69c71982d0a9ba06f0ca9d693eef8fcfaaa6c8886e83014a56a7f5c52275a1ace3e325d629b57e6feb66ff610d604bcd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77e894da733aad1bdd58bc681c0fa829c905dae6021a8890215acc4ca2f495260a2c05c507a807675d6c2d47c4d07fb44c40af304d72809df3e081486df270243ab3db688a5eb2a60bd5ec5398ae14bdec826c7332e1ecbc2890ecb5978791f26f3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6254e3d026d60f63e08a48d1f913e2eb8ff66d931dc2594b1ce8514fadc068e0d01c8617dd5b5e07d3361565d8d117ae5c4d71606e4e5bb641bee20502614f317c2de17610d972b5715d7346239b78ec744d443bc55fe20ccb6da41ab3ee7b12d5d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf69bec6460dd56465a2572395b8b24c14cf03481d94dbb51766436c1b5a832f719dc21e30274c2fc7bc902eba3199eaf734a5c4514179c862400a68a58532bbd3d6437cf1888e6aa06700c679d517191616f58f27521956b3423bb81d026d2123b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19015efa1d54cc2d28a8d4310761cef8f2d61dc414db3e8d4f787c5105abc7766a4d8112a8491de7248d67e011c411226b06b4ce39c841e65cef3957366e34b8717a7734c1ea86bbdfd3baebd8f5c88316ae2fde3f96a260d31f8aab285bb6cc0dae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bf0c9b63ea2ccfc73834a0206a20fb6e8fd7fa8a39ba7c1f7835f1ae412dccec7ca049503d89ed9b1f4cfa6bf2d11bd70f92654ff4ae7238ebb98fb1120528b730aa3fbefbbf8e728ca1b390f39bc6a100a33edcd90c054d3bf5f2b88b1c1a9f91a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3837ab0efcff407c808ba25a29c5d65e251ebfd883a83e7e3fd2b48677ff32f60772f27dc7eeacb1007acc95fdb14a14248ec2374ca911463a53dc5cad0e6a7026d933d89944fe60eab4f0dc63875092fc3c0aefecea0727918100655a55d316433;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21fd07a8dd2066a3191843b6391e0cfc678259710f406e2d0b4876dbc23c22df0144d4f220c374d67fd8f66b2fc63d7ba27cea8f35c233957168cb9b82756c08b12efab5476d94be866dda5fd6f44a1f4d3bd7525e25ff1b81f607c717536308ae4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha98980d8e3f3e8ac576d63caa62d51a296ead058ea93a5d198bff00751762c7f14fbc3fe0984775a71db47e307b2ddef85022a010619248026c3f0447aae0833144474e20c5554ce5a748aa0925f27f78c7602b525eeef555737b7b75fa386c1f85a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5db538ab742c8597dc539ea876d1bd19149b1f5859110e43341ba806ecfa044b814030ea594f7ff5c6c6743ba0f2bdfb1a5f90a8184bb200ff932f7f5738beea7459c7760920456683c9f7c39ace5ea114bcac804e1eb72b6a1efbfef79eaaeb31f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f3a1818809f9d5821046c3491c0ebf107801c55558620fb95f1b8ef7d0ab251dc2dfb625640232639c4bffe7f341cf08303e8d52b65f4b9100b6192c5a8a049238b071872d41fbb078944d60fec7f93a95a3b88dac4bc668df0ac767a718e8b6be8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29407ca5469e2e08f43cc83d00dc6c1727d0888a01b49984d7ae5eca7231e5db5d508eed3a68cddc3f5e6dac57e9431c931d2da501b6baaabb7b3c8318eccf8ad4ecbac4115d7ba27a70b6c92da8d2307d9cdd306f5b2ca88845432df722f9b8b57f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97d98d4bc47aee978c20fd0f0c3b8f334310096e529bd54420d23504699d0d29ebdc2c1e813adcb52024d28a532ac79ea29a4b47043f7e71b3b5886dd3506a8256845f4bd48d76beeef66aa2cc791703f5c8159946a206c82ee6b571378ac2edfd03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h359786e20ec966399d3b60c34895297015c123a471092bec79b92514172db75c0840f3014f0f57b74d37cf0605c297428c41cc9f48a2f4f7d8053720dc1c62e65934731855659b29b94b6d984ecc4e6e82e0a5d99efd552812f51c450b68c224543;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72786f4fa450dd38beff7b48bc856091dcacb48747d39edae78df3677fab9067b0184a63020fbd46a0a451bdefba2f30268c565629213abec1f5e9d9f72caf353a8bc83355ad5f5efd1b62a9d78f577d0ba07b1717e69306c355e42cc2f3a1f242db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec0b9ae25d803ca00e132772aeacab993decf4c609ec6e1076c1ef4185536dce77e8fca7b6faeb5123cda642fbe6378bcddcbd77b86a02a5c96871541ee67bdb6b3018d935afabd196d6aaae5088c3bbd43a858ea1a983a2767febe21e0a367bb704;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd64026a4d1fa870e1de6960ecf5ef6b98259d770df35a6e2a5b9bb100635b4a1a0c5a4a014fbf6677bfe2841c63dc70c3da09fd4abfc6da5658bc4bfcfd0b254572924d5a8800f6d96e2139c0647a8d99a8f884799a0b3e6e9a361f3015ef6c4725f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79ae5c92ecd296092952b74110026968fa713c61c5bd06ea9daf2e9e75a05194209076104c1af363f1ed4ade42079437556cd42667151016dda3bfd331d0847f36887db3635261d6a71fd9a78340746386629874edfc4107c76aec612638383a26a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3d72b952c89a16b060ffd1a93b8223fa7d29faa9b327fd9bafa75dff2b09d2e1011384ce609e807089d85c67ee984048d5f14468413112cb8e782b483cc978a71a174566a965335f4556f9d84b39142ff02350885f36addc5279ad07afe861d45b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c1a5c0aa4636bf642816ed22d6dce9425057b5f7b31afbfed4fdceb79aa50d515f137eb20276ad844a95d71eeb89c9d1940ac924ac2b4a8699b432f82156e0de787c197d900e75d3c041caf9429637c9326972c3c246682a4bef5ec1d1567efdb76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47026a719dfb34f2c83adc4ccd04e35f540ebfcc9fd26c0cc9b723e16ddb359cfcf21b5136840cb2da1c771ef8b27933cb28b4afe53bcb9bae53f1371cf1f34e2a8296dc9ee0c50b947b2d0867b7da19924908120dbc16981a1d7af9813bd6872a19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24691049582c3d020196c37093b34449eb552219f7b503a029faa0cf470ea13deb3656013a8db0615d9960d61dd3721590377559a08ca012cd43f6f567f336256ae3d4e337a250ecfa707868d4c5e62883e910f2524a7167f07b8f3c96422cbbcaf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h854cc63558c13d43e4ed5ded46cf50fcc0c0eb99f9df4cee4c9cb1cca0ac84435628767b4332983676b04182a9afbdcb90def393a8fb09401e70f2b5902e408c0b5843c0ac5d3f40b62ed5ea9f2a2e687581855350fe43766791e23c86962a2fc1d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha640c2d48791739b66e16191d771e2e68784f0bc0f3d911ccf7081cacbe9f5eaf696f73093e2eec8852d39bc56785e9696d568d834b49bf5e4d377462aac6e34de5c0948a6d5c0470c1220103f8837b97566ca184dfecb8f668599aa01d4efeb9cf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc24c87aade282f0d24bc19049a0f0ae2697d9640d294bbe03837c469c332791edc0f3b5840df419864787e45ff391de024d2a62aa15969b4a4dfd5f98db003f24b2977f5f6cd266c48e0dda15efa21f4c79e9ad0ef124e763647fb0a637c058ff32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85ff53f7245685f6b149e30a0001d944375ef8cb8f7618617de1ad53f6da4cfa14de6d110ae5073cee7544cda2944a52dd9ee6962d050fcf7cdfcba96cb17ad2909832944da790cbe52a5e8c1c234306e64f017b5456de1af427ee7983440bda89e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had832d9434c751c81e1ca50b1bfd23e9ee9955d94ce19e830e7263e6eff54fcf547317bd4fccfeb862ee0336a2a83dc6188cb23a018406676d080c84198574b2ddfc19b2b84c7f5acd43dd89e3585afead5926e0cc9566ef4bcb08a9a749cdbdc965;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90e3938113fa9958e9489ef44fdfcbab5a67a7a6376ab63c8208f668167c23573b3232443013cd97849d10a9583ed02e5e7f6c45dc01cc1777b49a850d721533c8c248ccad607655076631f7b9224bc30d20b216bffb0040ebdbfb303ded07a56c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6942b9ca5efc81596916f4bb8ed76374e633e296e4fa2974177eb3b96d451fa9e54b671ab2f0e86244a0f23af77a1cbb15b63c1dca234b55ab589ac030e1c99234faf5c8515316a62ee1383a91a1c7466ed30e07a90b76c744e4c2e4fe49a5a636b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b33887b0295e37e49fc7358eec7fa53b0469a06fa843d9dd8a1d4d820c8bedfab93e7bb4f2fef15c5bf179e576829b3c643096c10282a7e88fad7cc72676c777240699b40e8f3de91466af6c6af450876bb46fed906604d3448ef7eaf2a71f75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha77c690fcdefcd3be433410b7103d30aa10ec5988cb18396fdd945666f6756513f9a9e0f36db5ef14f8c82a17564cf62e8ffd0a0543e6f9af42e0032772f31e64c63c52c165040a263c325318c18a40cd33e4acc1c6bc92482e609812bf77ac48e5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6badacd9bcc1fcd740c8e6e0128a4651786a863f3df8cc11f2a118dae2789e0a3874e382385d479ae035630e63fac52bcf7cf7ce80ab4cf0f0570e8c1b7567bc98272ee49a628d26dc70d2c7f1121415a515133774689ac0c6e936b5080d032a2bd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc803c11d0bff3e472244ef34d0dd7b499b33aeade70347737633c71585eccfa03ec7f38d4b48015de42a7433bc9d8e6bd6e8893a5042275537181cdf3f4d61db57981acaa57ace7539db65eb9dfe08f871b8bd4576fb485d907517d5aad86833b9de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3104b3d5ab11ab15b25c75abbc614d3cf9b33df4e9bb7c18483494d2cc04795985c69e0072590f47e359344fc6d2fa78ddde3088b9c6208e573d7da783a65e328950a980ef9abec31cdf7a7a0e7fbe0db832558ed8fa599da5e4c3cf8a2aa6e2585e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecae52dd4497eefe71bd34ec762a76a954528562bb0a44961751911c27042867041e39273e0faffb46e8b0abb7221216b170724f08fefb0a262fdaa3c7a63ba9477ec07e470d84740388aa739f5cccddd29f36a38f7d6071df1d5cfdbe82693122df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h154f326ad07341495a1def9a56987257f7f38ca5b65a4138c22f8ec1cc5eb671ea38028b4a4d0dafa5fb3ffad2405331672d4a4191c4b5ae603a711947fb58d6fe81369273987f3530c30c91ee20c0c26add410c5c5086951987a1920732e2adedf8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b64a5f937ed7c435c46d6a39608b3e19cf18201f13f6b690b83ab319ec46fc9e3ac12da8c679dbdf8853ebe11c62f763d2a79143bccdcce3da676efe425df40f96647fdb9f56a6d29fc1d836c8f82be6e6a8cd1f761270b62ad7be39ca916313d51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2baa32fa0fe849a4b5a0bd15bb1f822612bde480139db9590222c361750393fd9008b6299d74c285fcdb009578cd2bd909902bc2fe104c2c7a4a9fcb8190e4961e7f8403eab82541d1cff6e06ac1a3bc4819d1909fc7f16228c652ef968aeaac824a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ce6e9cfdd43b19f7fc30691bb89f0a2c633ed0a8860c5c9d805a78b7d8df36a84f079dafc11f19201728ebb0459132a6990aec5e44c480d3ee0b418e97b13413272a63f9eb6dd3512d7eab0644adeff5cde56904ea61574ee99689a5613b581c559;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd22b210ffcb56dc2644f70e0f5928158e81a0a0a9302c4a85a690c27a0f2afc68b9b3fcde8244759483c8ef76234c02bee9800aef185366cf7d53e1074ee895c882749928bba99c069b4cff88d91a925d9162268b08470d7b051810ffc79b23aa262;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba7bc5653dfa3fc327410410962e7f1af64e41810b7372e548ac97ec29ac3a81e2ad28d2a3243a705e2a3e2261d831714bb1ef9852111e6fba82e8c49c531c81f3ff37393bb6954df3a12dd401d7517e40f16cba5d6d991d4b2f688e97f37ba6426a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50a42ad3a3979fb62e86f3e30f0e6bfe47346c737dd1a32eb8c11101fac8f1c4dc4dbc0cbafb96401c7f1310168d512388521a3835337bad196043c69209b0afeec869d1a9049c8fce2e2dba6f243ba763a9db2f353d59c8a28d3710f3b1e1210127;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3128e7d2abf30486077cd1815b7f87df253f610819f59abd4284e32e1861663933b09b6498e51db4c7a59b7515e7b7bee270d6ae9e34aaec2ebe7501bd599db29b5387276fb7b86bbf7445d79642c630b7bb1e534971eff12286a9be79f0696ea5f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa73d7ff5eb52cd1bf8725ead1eb503163c1b7c0ed7e0847c62db75cb89e3598ccea62c94e0be989e649e6d5df18500c8bafbefd1f91197d3846e815683f0226c8ddae52e64b11a57a01156b91c0c505742b3ba024333ea4341c3f78652f2d32353a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1807207246dee665e232ca966f4f51a409554e2891e9d4422083cbb3ee2857e611d55b39c7b829a9b79a41a4f4e454a505774328611da46290d8a7ce77dd86484eb9c02bfc8ea08dd89f4ca3216c1f6d62de9d651a2bb7c88b695ffb411fcb67817;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2054ec614f5768c5c576fedde3ff66a707f13212f2c9263cae5d598ec46144e6dce382f8b1d540033a4c020a8133374c877af77bc7f9a37a9832f5b09bf022edc69dde2fc5978fd1b2bef62e8ad579c0e5ee3928d472bc2a0d2dace1f058c34bec83;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d112f40a5b71b0abf7948df29660d55aec9f530d9dae4176af15408ee74c376d5f7668244cd3c8e92e6f6a1fa06662df3d91383abce950d257d1bff1522bd414e57801d3bc59d0d87cb3854dd955138336b26a7b19bc0b37ee47df8e5946e9b1619;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h471808b29ba63488c0c4bfd5213dda2cd3a78a445391d73f8c25740ffab9c01334ed99c60ff05b2e9c867aff2dba2f133e031ba16e50030e31bbb074d8a4af61ab5ca98e5e247121ed95c5359a2a8eacd6ab9917a0824b554031bbac1ec3dc809a03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83b43dabc967f4a856a4be713f0bcebd0fb784dc8a95e872266a8c0dbbce03173a1b9757ad122d9a31f50d1c8037e98ba8a0802f9eede9dd0ad442884e2e5e86f821cf6698bf7602178c449f1e888e541fe79e8085804465464c3c8ad73680805f02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ddf721132e8b7982ff680d7738b89addbef3470847a177da3fa8c9bab22a3e6a7bc119088e79157ec40df422e590678cb02e7a788e523ff6c974a2d599a6224770a7277740b69527633d60b937e5927be234418b7ed673c67f4a3ef5f69f6f443c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbcc317b0df7476df7ef013b7a32725cc5eed8e6c67cd409bcf02d7a1f0467d9a2c4050adf77b121cf65d8c978b00656efc80ca8e4b027bd35523e9834c248aad3044ae48ccdf68302a438bbefc1941cfec5b27283144338a920a95afde1f2543793;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa3d3304c6130733bae46ad75ad97a0e43887feb250ab6d470c45a1c8173dd2974a9668d2f32389b110bef9b6b15b264946b0b12acf2c75415480aa93207e624901d6aab6b21dbb58f9d918733516c37e23d3192af0fa9cf370603e899c707e8f521;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e2fbfc80fec13ea03d91553f64fc2d0a216ef90e088a567e1e949c7c811bcb81744ade448b2a4fe382c38f524beb7b32f93200fb85662372e7690174d7d3b8f6e0114c8ad63acc7b697387e21127329249862f58c1415e60aea1d30d93dfc87ed82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha526fc7a4f6f5ae59d35b9f6c9dbe74c4281a87b2a1d25c0bf8ea194fe772945044915ce844a75bc5c285b07fe339b62b96572414e8f7dc04324c90d6dc980a13c5ca1cf777c38898e89167f921c1fa109ccfcdc05554bf685b140208d9aec02c8e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha79a1a755432906292e909eb054ec34fc8978b8a7b2e1fc3af2a8e77692c9b0528b57543756bc22a8f9f28800b66e6da2acf25d92bd922c16984481c27a35778b6ebe719a77604d77826665e78076313496e3a485c71a45ab003ba40f41f5adff908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he889f87dd5c425b37fe2314d6f4c3fd18d62d1d83fab526f83178d5acf043e52dbc2e29e7841697f819768ba78eca04338cabef816b4ef05b0e732d7d42e0d275cd3786035b9a2144edc2476b30a81d4c4c66aeff6ea17a51e8c2dc1c0baebf46f00;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77e2d2f6f84b4517f3ac877a11f1607a508a0500adba73285aaeaebe4bccea6e3a0917ca442ff14fa77981e02b3949137b586071b58d5f020e752a04f4de5831d69e71a7ddefe799baca9084e8c7e5c99c9fdda48dc67a89bd778c75ca0597f99054;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h469a234d780f4ce88af9fcbc731ef325aef9e102399e655258041441dd00582daa495ef6e90422c4d6aae3fcb5cc3f32c76c30c57896b1b3b690b487e7661b76502e9999e662d92a9c16475e59385279d3b09a0c6b05f877dc17644cbcb85500fa6c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46a925d86e6f152d78e2224a07ff8e9223b626a96b2684710512beab74b7e171d91e72cc0f472fc85478086580cec7c340b9a43586cd5f56faf73b9ba68dfdaaee4405727db2c622b541aeffce68f8369cd35a4625d61fe1c966e031259e86b88c96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74bad7e60af713545dc8edb032e0f8f726049c8d842f0982bd92a8582c5801f1edba509323ca3ae3824c295f068d561fd1546b91c79f181587556f01f288519228cfacf2fdabcea7f3bd4937d4868a7247450393a76e0e210443cc0b8ff7b2f01506;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aa3f415974a1a5c988f274f52e28e03a99946775d337a4f755e76a86f4450e20d65ca8c0336e08bb19d03f5260841735db50168b7385bdd673a058dd08dd74f651e1d9d8ccd69100ea005516075bcc9a575a3eee469bab78f27cdc4d5cb7aa53fc5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b240b2e2e01f488e6cc991d1afaadd50580448848bcf5a5a032e20232529ad297fcb5500d617f6481b2711d604a73abc2f5ef2ead4799acc9b67ebeb7216e0da5568686d309da42ba065cf947b26992f4d5b74ab4a90994f081cc49952142bf075a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc19c1c6ce0fc383915ee2298b163c73715db8d9e64f1019ab8b33ea139b2076ca94e1cc6ce449dfeab93f37330f6b22c5cbafe82e83659e380c6d9edcc647385f1222374048912771f8e2a15fe9c0c140e1c135518607a20feb6172a952c2202d4bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd86079a93977276833c09a4943f02cc5680b16f9cc1c2a23431e5a1184e9f1089b1c971c5e988497cc855ca35c2f392bb2951d64a53a8dd7f36932270e1d2e0ae3935b2454a66911e717e79c18f4bbf31a2985509cdfc625aae75504840a7c061c7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74efe98b72310958383424b36ae6b0aff8884b1d89c4a4c9a525a5ffff6e024191758506d8abf09e2908b78444f6b9bec3763b11720d3d015a5d41dffec369505dfd0a35f9b328c23251e65e2b3c460e645291303b36f2b558f7e8b9c8fe09c52661;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd86fad3b6ce11b01f74b49e8eac9d60ae75712e9da27c76f6458359b7dfd72ca281f72460235dee84347a91f7071ba16a9f572946083f7d83fce61b0b6c1713cc9831444bd104aef3747a058ecfdb00d0cc23c1204b5219eb4429c62aaad07e5c4bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cc9fae5e98e2605b154f1a3ed2d831e3021bd39382129573f8b548d1821f2c73c37803e3ee2161cf10fce5cc08b3c86aa8afecb917b511069d24e321a58912af4250ae80f5aabb30bba6d2cae8b939ab9eb0e9868b6ce7a96399ac6bd3909d27279;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6871f02d1bdcbcce5df2f003b68231f9469fcf4bdd367d633889e1d34525c2202435f0afa6f523ed4acbcf98782ede9db4de6dcf2104cbdc25793b5c4fb7a25219f204a0c8717a18049b6ca86c1336ff32e00cdacba439e66b6536e5ee30e8af8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b53ca97bab039c4df69c0d7c189d6649e96124f125503e09748908c121bd160d86450bb259d8f5e5557e9328892ef1b7d2e06193ae16a96d859a185a577e42a8b28e36dbac7cb6931a4532fc0e5088be379c8f7e3ba9276464f11d8ee66de5938e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbae392694b7e7f52973afaeb64055647b443c39ded30e2505b17e286e29fe3af4ea34878ca90c4f2e0071da727f2f133333b9917043d25113d41edf1758fa207a1a7eb435f5c1f0d6f0dbdab44e2659724ccc3db6a93dc35430853d278b6a31db17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h577228ec6e4644b2360af515bfd6fa943949dd62b0b60e88afef1b5cbef9f8f792dff7ab1b5f03b03eb91a91d8c9ff6e6cd6cb96b2db6cbd76166a2759b64a786c251977d84e923852f2b4137f258cf8c0bd51bc2d83fa049635a02315c00240b93e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde21bc3a5b5fd43ac32706d9411576640b9a83a48654b34228df66d44257f3fa8eb8638e233196d9f575ea98e095cc09d4987bda16c0954b3dd9ece091386eea04fd30135531deb68bb76255a13b74ebeab902f3e9569d8be6c9341794ac6f96e48e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc435a9abdcd6b1132a628bff10d6a44fdb334f0a873934b0516d95971739863cd2f47a3573e8a5f2ed55b942e1d4eabac98adefd121a55799c06fda2315c125c9465a241d7cad9820e4398377f0750df3e58097d0d5978fa0e6c08e2eea284952537;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c78b8552788b2abdda9d5a0f71861561b4d51ec810d825062d1d46418bf2b5fc628437d625219448a2db35e438b4124118540291f25aef81910b116bca6d5836fa6962241f8ec586633e8525945c7f848c954775df856542383912fb59aae47ed2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2562a66ae8de763a152627df946f62b23cb2c929513223c4e7b24b05a478efc39f418c120f3a195c0d1f20e793aa4d4b505a8d46e1be45a73477c258b8ca8cafc5d381602c34919f2fc14247246f5bb39e63ce28d55c4c3070b13662f26851538602;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1eb27a00a0a9d1c672523dcb17d0f63f2848f7398ccf4fffc99513ab9e4c87cd49f11adbcfa2cfa2c79d2200045e0e12dc60e7f01fb8711467969b079b08fff082ac0253d39070821cf3a0acd4883bb6dcf3c9423adf22cf7972ff45ecc26a0c4a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a3b5f8d0515ec64a35a2092c90635e4127d8b1105c99bb3784ffc9ffd65876e4b6ec113bc83d04b89e39b42fbd7570221a9c2f787433258ef7476c95ec089020809cc8712b69d88ec4cd8f59334796f08e83ba18a8442e7bb1335124069334f631;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d566b9e6810fbbbc5feeb9ceff8def56e9e8ad49e5a44aef810812c6218e753b8adf0b1a4d335932d2e115e29e6ad01826e85b0ceb8af1bc4eda752c0e1a289eb22a99c9f1efc38e1255400cc0469845b8ef4ce4a51e272df8acf5c9a163aafdc31;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b93893255483449c7992c567c515f86213501e4cd15b2917e220f5145db5b135a417746b5d18aaa0b43f6297c698b2a0b1ca242ea7922a7d91fe73266b0e8dd5a17f428b8eb951453581b6a87a5aa917bca00498259ac948559311c3ab967e4b6ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf94e10b6e36b2a57a767a571743e0c923627cc9d2cbb569372de209fb44799cedd8469ee425fc45c6b9059d776cd50762bfb4af76698625fe171564f28f577da7969e5a835bcc0ed758ad568d6aa4d62d31f660b1023ee8aa73011c8a27caf980485;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5503a03547c0b0e377bc82d0aee1996114d40d94dd8ccde290e8da740284f848508445843263749675db436ff3586bbc01fa4b80e42c6c19fde062a91a7b6fb3e14ce85dba65838a601e4bbbeb1a121463c38971c41c20996eba394d0dca12be376f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ff4756478e8774a7191262bc7f128d1d221503ee354781b76dacd07cdfc0bf03575bc6fe2d6c2cfc9512d5b064d77fe861db08fa0d42731597ecce0b8028386c6505aa348846ae33f2f311725234d8f89ce344a02a0e4c7ef9ba35860eec7e7c311;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h837ba702b372ca98f031ba952b2b2152f8c11bbc1fd0ffed07db3cc1f023f35018b6fb3dfcb40080561a5b6bf3d783b7735b00ea4b07bc52e837e580b2a9c79bc8afed431a5736824fc2ee369213920d18e881801389f53907576168a01579a39377;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78ee6baa4e6a2a7e2e8cb2a0c6f8e69e2831287c7b6a797810af82b2ccd53bd975cfddb61631d9681bc7d3d70d1ae8c61d5a650d0007b2fd672605a463b82d2cba2ddb5f88a17c851e811a4327b4d981ef06463004f48dfaaa48da7a58ad45d5724b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d684019e7dce75b219fd5f4cda24f47078ede862df580a66e9692386d458333769ece2e2054224a220494906d661b4fa720bf40feac944b4ac35af3efa385ff6eb5910b9f3d7bae80c73352cfa4d77634706b73c74840601c5721c0e060fc110ee0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f2783c7eedcf03a45f55a92ab4cfd18fd812837b81f52e157cb6be6149a2b49cb128384ddb3cb2f88bd5a696e9db8667ea7c9cc093c808c0e4e3c9a1b20646a127d7e7276be740916fece1995b75d319215a72a44ff33fdeee411e6cf9b26e1200d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23506d1ac5f2a3e113f5d0e596e95382eea9be63cf5be3209d88e60d21d64a30e3f630fa7d54799156dedde525b322cbc6f874f6005fa341fff5ae492785e88869dcd73083f15bf800800c8964e0b8f69acf322fc6e4763bda4dc8da84429037a2fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27e4118453bbbafa1901145ee2c30ee3c0a7225b779e7984be784bedd1d9516d5a8f309302236ef2351409e30c3e424b8dfc94c77decdc12350f8945d23be0440478cb20730aa1b43071a2642bb38fc94da294df6af422ed3a74a176730529ba494f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564ec77336eac0bc37f5b1d21151fbfe28476660a62242ee8c07493829d5bda7327869cb851e91a85e605a4bb4f669f175426ce5ed35a40d4687b6a862ab0f99a57a8d9dfb1af8dade3e75fdee76102f132f85e08f7416f2a253170f518c393271f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h528d5139cf6dbc0d55ba93ed7b7f1727d340a6a0f40e3098feaaceba6f1a0277dca7ebb1ba4ee2318ece9e4710b8fa168cf502544447a76f28911def2ae2448b32b9d793ace19385b4503c0e4c2ba258bc2bd4a4199e294059902207a5178d195a1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9699e2bdc65bb67fd5cfe4bd7fde14188b224a95a0a0d9bfe581c9d4a774b81b85450289d860cf34c3b7668e8fcfb015b3ddf55cae1008eab8d7ff4f3c779baba89fdb9cc0790cd4a90f30aee65be95630c9eb6a6f3740bd0198ee1f62ae0f16fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h144b14fd1b129b247172bdf33a331452f452e647325119c2d38bce3e7a24300c6b1ec2d7b6c34c0fe03182353fdcdb0e5a8b3df74bf5449d3600e2bd4522488ba26caf8e2818ccdd9f73619546bce38857aa3865de62a4186be0e428d47709c1f72c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1df7e67bf43fa141f7a91ad1c8c5a173cc4c745e4d6792dae6fbf04b931af4a8c31bdffc9099b488b7690c0d073ca800d668267cd169329c3d919fd42f412f53dc62bdae029a75876f6aa6697f29ab78c116fbd1771f302de2b1837cf00f31e0e60d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79ce96267ef4f7e3f4c79ff17ad732eed392f40708128763c00421e2ecb1b46fec8ee59924593a73b3c9e6a344672e4f251b39026276d213bbd7e3d2ea64d8c77e17bf88ebfb134e8845bb7452f54f301ad2fdce69d303e2123aa9981bb28d81971d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3803953f695e69aedae81daa4bd58b6c1d7c34fedc9508fd7fc825230c090f29f3ab21d2a6674e468fcf42166e1ccbf9feec55d305cdd9a9b103fd1e5e25bc9160bb5e39d55f228112a294040184f7a4d71728716a9e8f3cd4977bb33fd5017882c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h954227d10b58b63352f9a00475f0412a6e932814fd91ac2c4014f2152c24f1486e848bc280db8b645a382c3bbd869ca758b0f9c11e76dc1d1901fcd455403ff43299fb79f0e76427a15910dda2073503cfd1416a987a0c4b6003c50fb357ff4167bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64e1690c624747f2060d77fe03c03024faa7b10075d21aa3aefbf90bf95078f2e981e9d6ee31a11e4688e32e743fac60ea71acb6f7acb2973f0fe638a4d06d5c76c714069d9dd807641583511325539b148371e3635d7bdb4bc0ae4a7d4e0ab5d006;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h523d9a99623a0ed146b7e1a734aed6bedccf5ba8812701823c88d25ff70e5e9d41029168e34d1f21d91bf3d439151798ca0829f592e2828536f3a9fc9e0f389d1ddb01b58205ad5d41497205f1824eef6611bcec043f83a88b20834540187abd71b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4be4fe44335c359b27670a0c80d760beec79e8985e84ac3f0208e26594b2a300bd479f7c7bd99bcdda90538e192799e3081022d0a5a911e1873dd0e08d29c43a80e099f7d91551f2e070d05904f736fee472aeefe655dc59d40e8b120b926a4f8018;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h128923673e412a8a630e61b9b4eaf471389ae4354d95402464fa0d15d518a1a90cc50b4874450754cb291ea1b3657ed1732fb4f96102374e93e50c8a7a971e4d0e5ab854b0452db7c1af83e1cfc60e170b467d2782c9b8296c4460c8619cbca3a3a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb47e936a4a101457a775b852cac66a64416c337f342188da88f9346eeaa5d28309070faebf578d0c6f2aebeca996197ea51480f06fa43817ee940fee03d75cdd523314f7c2f12f4bb7dfd1c74248b7ed4113c42e3fa7c7f4ec0b9a123ef67b3befe3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b4168c4f70947627dcc96988a47660f3d965f458bd3c99efcc8cacc3bc8fea2de5e462c119af12f137c0ab090d12289267ac30a1660b249ae82843eb756683b38c253d1e3c9d70c20cf078fcf4cb220c5ca498d22b1438cb4f974200c089b8eaf9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefc3dcb97ae410c0d0b983a05e17a405772d1ca998ea3821ae9a18722bc3f7a55c4f14b6e841841c06be418d3fcbe8dbc7dcb10df9d338f4de4aa74b660eacd376c6cb2490efd2d958ae5429e73d14784efb1e41842da05133c0b1b8612ccb7cd4c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb9c847d57fa246bb7b9ba03c89ff8045a70ecdc9dfc61873dc77a6dfe1902216c7623f3ba83004d89b3596b93993ae743c6344c4ca38398842d9fc05f2b260a47ae7c9173960bb9635b2afd50425700522768d95f097447dee85b45471b09266354;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0928923f66a09b6cc0329c3a14b46b8f59735b52d439ce56c349907f74461b1ff075c9757d9346cbd0f5a3655fc0f22a342b4c60c98e79f2f2cb3e91083ec31008d477becb98738d910092c1ccee2d18480294341eea319873c6053824e0818ceb5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23fd0af38358c7fe9570454a49ee8c327a6244e02e7e8d582acc80a7398930c25b4dd94a8aa8cf1537022cb302920c348b1f46d3fa3f32802659bf9887482713ccd9de4b4ec3f42ef9e1674efae63d0b275c75385ed3d6d3cf7a714811e222d84f02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8df377d3d7e063a2f0764e40459cbf55eeaad69a2c4f0ca47f784725f9ffd18be33d80d380a772bb635cdb9fa365bb3457109789c52109dd6613ac437f2de5078f3982e323d386bb3a0e2d9af794f99c075cbaba6e1c8db3484340653b6152fbcfa1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8bdfdd998ff69c9ca132dbbc56beeb63743d8637d895bd80ef9d6f12f0be5543016e994d8ddcefebf75afd30b1d0e10af74d6ecd9128fb41f56c66c0f299b02ac653cc252eeecccf3c64777f83bdc7d238a31408b1106195aac637cb612a3dc621e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f328ed44c3c1f6b78c39d818ad25cba34e36bf393ed08d11b5aa474458d0d505fadbafb03d2fa682212a99f7b37adfe512597cfe581f40c0569089ea4e5d7bfeb954de14fc53dfff2297d081cf1ad01d77680e2582dffc738a0d51725f760be9d90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71648ee608230e668f3451e9c37eec80b09dd08394ae14a33bcc3883aaefeb31906ea5c37538915f65371a20b2a91fcb7189e6f6a59c1ff93643539878f920496b878f22a01bc9031c83fcb272ec9fa165fa0bbf4d9913bfe08f658a602c58103e0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcec4b4f4d1672651a374e193b43488f5bbb1efafc09b479bc99c1e013177d2dd3fe34b259c89e7822ab11b8d3cfd173f6dbc6a115af1f664f4b55a9dbde730db3a737b2402bce0f457b55675564e0f712a0a680f7475b10693bfade52beb39f2185c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c4b976fff36965c9eb8c9bfcab9b63445260d41b5b2d8d2540de7a902b1edc3239d2a1e226992cf0aa1d098cea15ff523e78f4bb230a79f70fe769461fe5970fc1f3ee26336ddff5685e5f87589e04827ba55275379a6936d32b0878aba9c7e7b14;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he28f61b1740ee53bd97d269748fee7f2d211a8ab39a175fcbd2ecbc1d3767821f18edc69f9acfcf22589105bd69ab17d3fc005828def67538aebb7d55190e1baef46894775d707da559fe60b3742fbce98a17476f7db4bf6f93a4353a1662bf1ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95f38129311ebd1bfdca939671617c719e555bd477cd52abe3ecef4221eac3450f7ecd8823e95734e84e1af21689b8050ecc12473b19647f1ca7fd8cf5d7368a32bb83d2a7ead93e0c05bf61d3b0776f099da5c9e432235465bc6b61dedd31c29889;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd06792a07f0cdf341621c2a8d318bb6e459b27b4d6635d6b647bc6fae4d5cf69817667ac546be1c0152cad4c60ed967c205edf70ff283634f196b8b74daf88249851227168960886e376fe87af832e5af61b9b3eb2ee3f648690f407769756b226a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h869359e0b78263e7a94de2d9f92fc52d84e31fd23f29be52ec4860afa629e76a39d232ee26fdde828845094f774e7d3c3fcf8e7618aed35bd0a313e024aecf7b10813e6e6bc15949f2a5e601e5698d729a50b8ce38961d872159b9cc3c9b71092f79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6836a6d78f61442feb3e751303fa427d93f87f07cb4401b7b9ed669dd0f4343e1ee4a735cffeca794821a57b687b89852649e1d3202f0a63a063f0e84b993df4b7c1d124fdc925253fb1ef3148ca409edd87aefde3d241569ae548410ad648b4cf4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c5c82ca52196503ddb67d268f11baf27220e7741c84132f7be6ed71b6fb68a241521733036a12c7bc00e0d34d978adca9990ab3811ea3c50f95f2bce2ed88afdb83539cc4bc0a02ac14a2a63592694de5b7feb72e6572bd3fa00f68400155463015;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7be6aa6ef3cc2656f184fb7c668ba37371da82ca8756075feb6cf4e67273e880858464a989e8d93ead031bbb4b17e0caf856897379d1dfecfd58da838aa83f152ca7bea54131a06b5668e056605d2c3317558560a471394e71c5b47c13c7bc2becce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2751da62f47e72155c72a2e618fc75c6919032afcd9480fdc013978b2175fb7bd90c47002bc47f5eadd26fb1e8ae9782dc16c4d9b31cea211977cd1daa8e72a4f164ca479b976bc37cb33cc2bf04437a5ecf8dab2f8343e703951ad1da4fc04bf261;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd438a96e85594c115ca3adbe7289fb9237eabb526ce5ad8152e515bbf906fd43a61e50fc04a2ad6f00e025c3a0ebd5de4a84561a399c6ffc51074ed35f8312424090a31c8d222664fe4f965eed5733aa5df55ac1060f1af8e5d420b93e562f5f6f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2f5f87981e284e6e5728c2b35766a72af2b0ff138f30102cfccdaaa9ff3023ffb6dfc570caf45f1d71cc009cb3b44fa85f284d0b3a46da34560ecab00daa75b8e3fc2e0e7127a5b9bbacd7c55031ff6dc4207a03848860b3860fd90383b4156f6e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecc2103f13cff2415951c9c0aea9bee2a37292f5e5749fb2fa33bde121b0456008cfc0cf868997fef8aed605b096c8f3fbb0ec5fbc580552a5f62338df8dc107d461138acbc49ff4bf32c19333e89273504cae376f85e885ac93c31c4babe54dcad9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc37f4650c1cf0315e8c1e00b862a2b128b7da76de7e96dc070145acb84700bd55dbe781ed9999ce4f3bb76fc078defa131b20cfe395a64ad296e46be901c39241527dec2145f886a45d81d78fc493691059922903002d6ecdcf81b0ebe59b6bcae2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h399a26b55d28be287fbe93bcba37ccac78f6262413ec40ebc0c7c78228650be38b8de863a5b4cea56535a6dd1d0371068c33d6d5f3c957f52b4278b66575a50ff7d5e452710808529612fadca745f2bdf4bb2e64f7b8f6e86aaaf858bb9f1812520d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8c3e8fb7108940efbdb73894cb1a00cbd4ecc3f029d5dbf1cb2d86183b062bde111921a6e6a1df447d02cd4b7f5f93fae08106cc7491d0c3fe1abc59ebb4072e281af974a6a89ed2524e0ae2e39c8ad4ae80be65447438f16ec63b2d0a22edf7e75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h307568d62ada3ed9c038d695e1472d2d0f0cb07bf0abd0442d91cca9283346a946c901544168962db11860ac576c0b032c8592126b23acc5c3905fe9a5fa19060ca3122c197a70abe0e19a74f8c3b6f4c41cadf52738aedd36e8d38772c18cab6bed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f633e46123cb6273d052485f312979b712b3dab72af21edca3205c1bdb5431f942b428d2c2e62f67a719ae8d46166f50f0f11582747b3bece39e0de5d2483b8e148a2882b8ef7822f5fc35d725db7e4e82308c775163a94bc3fbfb1dc0765cc6ff3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h548dc801c25066019a23c35e5a9227df8b57e22e46b955099456a41ac0ad6bcc482a40c3504834260966814f40c79be3d97cf85d14f6bcd422867f0b10edba37f302ef8b062050d8503d5fa45e9d4b71b30b552325516be95553d39a10581183a6fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7b0176887b16c9f0658520f1697d8b9c75996027091dc0a6b9d7a5fba0a42a1f612401e97d3e85cba7b3f88efa72812dd6f63662bc3b8b7c785d2d8a3e90f43c8a27b97b77eea37656a3583d731b5856b1198236d1219bf839bb31f1ceb89fe8f71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a8c589e876e1f5ae23cab91d97d7d78ea1c522f2625f0f6cf119d4427e1e1792af215a9b0deeb3944408ec2646bd8bb3bbf5ca5021c0f4c3049d9cccc0bc7788303ff6f69f6f8a8d15ac0a1b6d019142d43e7cebf57ea97d2f2a2ba7782a2c3278a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he38b019b97c3745e60fb65accaf54f59840c8cf3c9b5a872f20545850a7e884c6aff099286f55dbfaef2b022cdc4b00748181bff9ed10aebf031eb9aa04168fe0c9e4358344d2b01ccfc5570a700f5821e3fd1e985b952f5e33a6f4fb103e6ba65af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bfe2fd18d07eac5f79fda941738c78c5f33694841aa7cffd02c8cbf1be1b2c12c38bb46439d10adc8d5575adfb63d14ee261f5c25645568858fdaf5d23cfdaf7c51b825d3277d6bd9ff40d178613c21f44e03ec38a9c025f21f5b17b6885ce8f2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d9c7e581d00589410ac1d327cf46b857197d6b9cb1f2b954ff34fe3f1c131c5627b17dd879fabc5b4914bd5d632a7790fd7e030dd51e126a3b4b341372ce6461ca7e2e82cc3cabe8ecf1e8ab7e2190ede1058f8139d106b277cadcd1f88d188f6a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd03ec97f9b80503bb39a5b6d0c99d447f32a38a93d87b8d11ff23cfbbf8c3b8ece85b8114df078be0fbfa481775b8a24aa560718337486466e724e5de2ee0f9b7c13e55a9e72f8e9fa5c64ba2a1ccf3f40606461d232ea20853feb23e964eb4a79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57076bf962ac6338373c8ad30eeecfa3ce634c7f0bfcc7fc1ce4cd1358004ec80e3c60bd9621312f49b96b470c1b39319f3a7bf6d26309702d7c2d7970dfb8610e212ac7a4f97f2b522964d548c060369f8b7d6c31afc797e797a6c5815d86da1ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dc20a8f2e376cd6830c53dccc330152939ee09780ef723f63741688f23e4c7efbee389e5db70cbd2a559377e70a8ea10d2ddc5a1bd28070e4652f79b70933ef399f244e4894421065e33b49577568a9f7abe2c63261d4f919a0d8e607b1e21e345d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59dd29889ce25b9e2e62bac6e39f7a3f8d2670e12ad02b77420e0f4acca63c409bcead0500b15fc8788c90c116418694bb53f275caabc48911f76e26e77c91e171254ddab907f00b79522590fc469f738489821513a5a3ffa351f8c98c80fb611550;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a331b2eb2b31cc9576d930ab88c2099bce2fe03b281439d88e724f3e09c3a479801243216c0ad8d753d5eac82d00569747de70d8d4c572d9328bc4aea7a50451233383fb2a96a34da6015a543c203302fa04be99402eeecfd68e6972d7dcdc0154d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdad50b250abd556de962782889848b26e92edee0176e168ce9a5abd8438e55d96a64adaa4602b29a9e33a287aa2477874757c318db6501f51291479259081737ce36fc0613a15ec9af83b49c0bf9d10440ad218a53b850d2d3ca5341d8b13f7c583e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he064d642e13314422bf4a0255f44900887fd2ea9cb222b63c1b20c1ad03f44ff2aa7ffee78a9f8090a72f2a87cc62cd49ef33c531806ae1d2d1ac388d5df7e8816f6152fa4318ab6272fabc3d4caf0fa2bedfba66855c5835eb3cab835372cf6278d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f8a60f4ebbb45b0af22b110d5fc349471508d353fc9c0c4efb091bf6bd4e5a2abe114f2eb1ade809626bf9f505ce858e3b9a84336305ec0444e9cd392592fca23f4ff835d32657aa763cb92f27ed0f324e59961ca381cc75e145e8a494a15c0be81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2cbad07bc7e94ad80fdb2ccfffc79c0d4c7c88794fb418e9c09825288d07bfe88f62d191a358d3ea4b498408762e01b50af14f30428fc333f0d28fd71717d9e56a4083b458292d6f9d0eb37bef624d9bf6cf25f0c4cc0a169b80f9791812d99c7d99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha84634b5299f88dc049450c939179106e55eb4c6438420a4ccd9f6971f69125cd538bd3643799b591346f40d488213ea9ca0c18a773bd9ec28eea2ffbb56636460168613be822edc85038290f44ef476ac3f896b0ff636a0a05290b1e3e749a7c8d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32979969158b9593a799a47f4c28cb591b5ac4f1ea700b4722912c0a9af05bab55dc1428655d95844652e315e16ced62a460b05f7904bd689784dc045aece96fbd98029485f1ab81d2e835cff5d1285164212e6c52cf9bb718865cebef696c7b6fbe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7125255490440e43a73d7dbfb45ca504be3bdfc082f5b2b743f097dee0255eabbb8150fb1e980565d337a25a1f65e1ddeb01aa272b2b985cf799f5d15d6417b0c88a95369e14f56e362cd7d5f8d80fabe42251e7030c31dcaacc129f6703342d2aa0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64c8b67a000b388e3b05f32875abe483fc868117f5d444ea8cd00944b33c317d94e7aa5da0e7900d991a626145a6cefb249089f330749141cb2d3a1ea4e49cec74997a7bf895fde250830d98f8aa137c0ea3f29c52cb4ffd00e881b646ecea1355b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1049ca06ac4e64e0f20ce8326770f7eb41b2e7dd32536d07a90a9cdad81c794f0e5c3736d6d3e77c9cc94f9eecb6d7c1d136c82d129182b7cfb4c3a98c277bf1fa7356b839634bdc98e7ab06f79d810436bfe0b07d182ac1a83f304bb3da49f99dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1fc577ab3ae18625132454fc8a278369f061e36d3378dff0553b56b0f1a7132c8ec6643e1ffd36fae3e5ee78687e8df18ad99b49cc7dff062dbcd29b3b8936d6af9367fa3830b9e9f50a034e27a9c3cc2962def4a31d12704562ecb9d52fde3f505;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a4fa53e462771b27bd246ddfc316847a61309957e68c9ffc7b8dd29f868f332dc8582fbc93ef76283f91e72f416ff7de1bf366556fdfd0d3ef7ad29fe8d81cca21f5decb3c1b27d37eb49193831877cfb5f8e0aa641c140a751b785841b0dda1883;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7eae10b2a5a800bcf65feb82041920c0d9b1d16054e8e88f11676a21666c0075717d415bf80f36455916f3c4c638035ab5464fb56f7f77f5f3487adafef5ee67658d48232802d82184c185dd062766eaaf401fad74bf9d389bca436370df22bae915;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha19f9ee7831375d076d8abf05459e4b1331c1e31907ad870c741ab9d927d7b5c92222fe2e769b78ecb3ed7884760f2e6d565dd80b4d5bf30d93162690d77da887286240f7103660c28ca3dc52e64ec13c3988930c0875c456cbd0f697c76ad824bd8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfdfb86d4cce81250d020a4a2c6a814adf1f4d9bd86c1e899110c2b7bc18c2ef0f2b2c74196653f3db2e1e1b4bc5b971b1a4103d1de8997fd1c174a6ffae7b5995e668df9cb237b732cac9345dbc2987d26622cace8ed769f3bfb437e2527153bb2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e123d2a9b9c0b3cafb92c0bec4e2ded27d15b54a0355d87596c3fe2d8d92500b3483c0653d0225063cb2d5f17b9b282c4abf8f1f3e72e58edf7a6370ad6970d96132a2fac00d8e85a26d99785ee83eb13e4a564528ec9a0b2b85d4237d1f012f212;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h834c7cfa82c9c98826eb7b38265850d9447d7761345e8f498a2780a857c90b8a2bfab712098848714a25c4ecea4bf36df69faaf7665a52195f473cd6112f89a4f546c43999ac993d25202f4e0e24488652b93f55357a2a8b6437312500d1ecc6b5af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48db618444c851161de1d42e60a958586bb0d0182e9fa77dd1a14f6c592a4127095289c19f234c7df1056f25eac0630cf395e2b7dba154d63d43e1b1e178c98eaba44242fccfba870f074208db76cab1c331b23bec00996a59776ec43793df545f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h687fe38e2bd3a1a6566efca548161a02979dde8de2a003c320c3ea2fbe6d741afd6afb6bf5be7a7c6fc8a9696105a3e145ac4111912907afacc6237016f028acaf7a8062640978e47ad31738ec891747040c07b30456baf66b57139bddcdd54bf46b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88b22c8c5b6816f3ded7b682738420ea24da07f03410a27ea974f7a677ff434dfe085a2977954528c38d1499f4e27f19f0ff1d54efef6daa06ed95aa3265dd4ebcb6a07da940044e71652f220f27765d44968aa54fef2eea3f1ea2ede9d8b80cc31f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6868aa88095382692513f1f250a9be35af393853cc4081c1755b65d391f62993cf7719afa30a60c8f3dad029e59410a2bc0bfe770d6ba233029a4258ec33681408421db511506bf7f9255a8d4414f5989fe3d6646d7596e94ccf10658ba630945e1f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d43a9c33d325f49b6f20b2e14ebc2fc758da68d701c04799cb2c999f12dd5003520e995cf4af57a88d8e50c9619d35da4603ec95afe27ea9123093e8a9c428a9cbdb078abcb8cfc596ea9bc8022b238da30a5c89c106acbda02f838c1ca90eedc34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a475dbcb266f16c24daf7914a42d968d4e9fcea7db553c2b05318b45d11abc621b198da93aa7688c2f2fce14a595bfe2036d3b94a1d19607962da2eab04b10d49b66c0055c815b45f5933e08ca3aec5052c5660385cd652682a1baea10bcf44c8bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h463950727c30be466e0f30efbfcc1c3718a41e99c0fd29f6d669c45286cc28981d40f64eb28a75eb4027a7a275b1f125a3ba1fdf49bb313f6ead95b9f8195284549dad1107030562ee5139cde6d2a5149182fd586b350ac4baa38efe1898dc55ab30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca439f550dddaecb2e78694294b7f404ec2f86fd27bf0080f3384d4859290cf50875641647ec56c5bc77158ad648f9c862037710a5984d4d74fad76baa84f89eb2557987ac495092352a95106c1965a0a3add0b5453afafcd61eb86b0492ae6a9dad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37c67075c529abcfcc1054d224bc92a963a1b7d77f66a8fd379a8bfff5c3d62f55371d5acb7b785446b85b8d82ab7563cebf8d805068839dbb7eefd6e52ddb09a83268bdb38920e3a3ef57ff5889c1e6bcb71eeecc7163e2be3c38e7d0a7c8eeffe5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dba8269ca7a6fd48b4368206a96af9451b6dac81a12a2d2f74776bbc90c41819a4851a2d3cf62cd5b453668516782c731cd00d0254f305c73bb40b2a197c819ab010ea35f353ac83d07928d47010ea032ea4240530a923b5fb9736d8507db40fc47;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ef88304fe8c8958a879c51f332bb0c57f12a57d96991790ea2851db60f71b01b2b9f95d4d0e2ab5b6856e70ab5fc69a3eacade1a7674c872de174ff43da74d0e3e50f645725bfa579a7c1d8d5605cf6ec39862d791a776f901e71f43b19831e02a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he42113f1bfaa99c2c14baaccbd8d92051c4009c983952414eff2483cbcc6a3e5ec31ff0bc13fc461cdcbb752d68f764af99d82b575f3260a6c8772d135afdfc980fae1ae8ff881b5a383513c81fc20b839920407afd1b5bc6694ed4e0e84d003f792;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e8d965e17a9ea97ad832ad85fb7700ce73d3595e97dce19bbf17ca9009095438cf48f1233a817faa8551f5812a23bf24e76d81260e890cad2aba93b955759b5856fbbac742a971fee2820ee127275eba13dd396b23359b67689a48d43cdb21431e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50392befc8f2756a676e1a614038c38ba4395ce03ea8a21c6fd7b4044a1865bc5162dca0be9f194945f60e01a63d11944b130321bbd534333b5e96b231b8b215dc375583f28b80b2cac0e36a7582b6d8577ba849a0cc734fd34fdc4efc89deaa755c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haef3c17a8e100a5bd1e0d9639409c12e4b17cbaddf7d2ff136c92e6f880e8b29ef6eacaff52df2ad5716c0242a81cdafef111b20048298d0de85801d3c058e0f06e0d9eb5aeba2c287c4350f60d508466cdc9d371231f8cb07caf6755fa18f03e322;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1777f70a77fde69639dd1e2fd218f86c5936cb8dd4935a5f671ef0bd31a7c7150995289932e9123ed9a032fa8c850b1970a768d154300cd47c1d23413c2ba1a5b3687e3ad6d49f8a1770b8d7200d205b78470b168851282ce5af6f71a5adeb10506;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58858617a67862b9e859cd2b0b686fb707009eaeabdc7784fb1908d7b4ce72f685422c06a6e096d7780a1fe5c426605b0a9e9f5d645af244a8e76069c1b3e7a288456f06749c424d68f35cb423a1cf3e72bbabd7538fffc3e4db7adb1e0aeec71e27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fd07e0562757eccb48d4a95a9d428f18ab10cc14271f074a6ca5df458f1e9ad890fc61a5cf2ada8d9983ba37d18a8205cc64d91aa39250016332deb9507b0fe9f7d3dfe17e4e9bbbf56c00bbbdf540a1135ff8d085577abbf7079e29a95107b5fbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbae411a93411461ae6273e4a1b140bd200eb73212aa3e49a63f61017cf96cd051bef09bc883e6f9106a1732f51535ede2f4219ed0803ce5e855515f754b0a3529e80d0d9ea158f877432bb9203d9a3cb25e3d8ba01a4a4f4f32107058334433ed71c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha53cd925a597b3831f40abb65fde044b5e0e60c1ab43c8374115caf62dbc934cda130af6963ca076cc6d97fe9994e995ddce882d89fb65f3b909bbe935d8d572c9bca7199282104225eb3d037253210aa7b0ec0968c6ec5e7fb2479c89208e839db9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h188c3ae2abafce97a5a5be46b16231a3a36806dec229de00ca5c7164adc2273fa2e1511fe9497ff7858fa911bb30ccdcb06bf192e7ba1b5e6ae75d2344bf36c70ad7b484f475a1abdd0e64e23250f2ef2e20568a1a1fab8fb43f13f5f283932b3495;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfe139b6c478733e452608c235c3ac02b6a1dfcbf1f8752586b65498bd1fecaa6121006edc4356fbfb1cbd6a7891f0bc5e3ca7dadd16ed1b20e1576475a17665afad690c6a0277282c4963fc884ece5db3b7f0a9f332e4b2ff7dba555f8eb2752a13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he04a032d547deedc2767feabf53db8f6cb5aae4bcc05ae1e02e4ee30927920f3627685bfbbb710fb329229196f302dca2d0794052192debe007ef520bcf67155674e37a2af2a9506c11dcf9ab172f74e27d5f45a8b604789b852d8d24624dfa0a149;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c3b21f21470f55def76482ef2d290103028618deefdd6e02dbcd53c825db38520559be1490ae186473a338de5099626f58c9a5445f40ecc7a9dfd0fce0ac022e5e7ee0aabe1f7c4a8f85343b2b798a48792e5415cfaf4bba75da90b8ec82c015e92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacbab1adfaf0be7917785d1e5e72423684d5e9f96ffc34edcc74f7946b38f7f2473c3e834b91b514032734b2afa480934e68213f2f3a50ef22b426eed73f2a4c373d089de913a5bc6c74decdcb2c1823d063b85dc1045c315cb94bb5dcbfeb913c8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf81098b861ade5b2fe87ab5618c25ce818c8ac5029e2a5bd53c5fc5eb5ed439dd32948f59bbcafb0995642547bb38858574699354e6ffae7925dc106a08c6abb254bd636be1506f4b79d55b4b030a07b85430a300eefc64b6832a3e2ffafebfbae9f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19b2b21c828c102f2ea31a15afb5fd597747503d5892c964e5f40c2e0a980283109f213c3cfa89558bf2a83e155676400796c6009d7af4e361d7f77a8eb98278b4dab549f40eef0e1efd8111243a6347bbdb6eb2b8f70a38b209596f47147b383c0c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39a635fffc400c51ea2e1a0b6ea2a3e1d547c2f4c677636256139e49339b64d7fc5b8bb5d9f34492d01e4042a888725086a532379ca271bf60c4690abfeeeb1c2d3c116d06a816fcb592a5450e1553872aa267f75378b40b052adc52d239421b187d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heae80d3d906e2dea6e2d993f539f9a006390ca2058243f21ab16b62e4f6fea56208d7b20a2dd618554b7ad0525d1f32fdfd0b09e1313a6d1067771236bcb684ceae0372417880cca193157d0283a588c071b8dbf77ae3932c7062d14ea6394abdf3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had054e246f904f4a60062ff5a457efd5f4e1f85b7763837e72d14f4b9a675e128533cbceedac8fece4d43a2c1b630a52c2b58053d9c2456987710067947f00ed558ab436d69720e6220ab1cc2897c98d6bb2a1d9bcf5a85ef728442c2012402e770c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73ab79cea509cc65f0a03328c0f38f2f1627c87ec9c33f991a366045254c8c0a8f71ab63222bd2d8842e3724b5154c80e9f0eb9170e9e9c309279dd6c1f35576342fe90604bcd91520d79f83eceb5055a708350531d99ac48c5a2efa7efa1cccf62e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf29366dc1931651c127eb7709355ef566e00363ed1e9c1ac8004384e29bcfb1f11513addbc4764d2e000f5993c28679c1d5814772a07b370841b0972e1b96fbd72e7158b442c91a3c4c71d7d8dc74e522889313628553a79b1a1d3c711c98c057d68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha008e94d1caa72d2b87ede03372ace0b49c0df9ae482a4d08cdfb9c199a456af4be479ec55a29fbefe4d30670565487e9b4191bf147398edd731f1a76b2209144dd6050d7982a90c6b71c361eeb1568e0699ec1711c9c4672ccffbae8d6b7baf15ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h601383b85a36b43e51c761d9c2fd919ecca123544cdc0df266d813cfb7cf755507ff47e6e03012c4ccc2d4192d50c0e720f56a04c2fd72324da8634e072f8f88f0aafd12cce8b8b4a47c1f5ce7407c5879eb6acbe7fab46c565203810cb2df5f26d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha241102de8b1a1f2e519edb80460dee1a6b335b56a59430d65362fac41e379ae930fde9bb4d081c041fe55154330f5a9152b3dd8bb7fe2d9d4e83e95d30467af246dbf096eae27016f67ea6efbc7f63f93c2b072eff18bac323d9628efa3033ed9e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e83de56c58c6fc292d89e0727092f1a592261b98e5e53186188477f2e6fdfb2353f1909543fb41f6a0645d3e25b01f90d389901cdfcc40bf529ea0bf4c9c5086fae03bde9d6b866f79c662abfe8ade49864564dd5f0f0e1877e06d51caf92fee07e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec1379073bfdb0d3a1bc4bbd055047fb127b1e53f10b2d82d9b3cd4f838755906977586e6ebb4219efc8234d130436e252f48f059c99ba9c0470e358cacef7bf9dbc828c466c8038739c8fdee572109f9a03ef091761c4b2a146d7cf2452bddb40f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h177b23b6042e71a7dbf54b4e30e7d62ba51450919f7a95e9445ffecc479267d5dc3e9670a5e62f0f2534b47b53a7cf9701823ab418d8645e284a7ef2ab27c66300325dc23869c4160602b79049dc883499608dcacf1c57d215a96b5e173362bc315d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0005c3d5bf6d6ec6ad5a8b419c6277cc90a6046766412a07512fa49462394c54d6246662ef9b158f0c0652d6d40d52f4774302c4be301f81a1918167cf8cba29d89a01e39944a988ba531d845bd227c24a467fec7486363400df8e8f0bba5eed421;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h881ed28ab40d32b8163bbd7bc5e374b6ec996eafd98c96bd4d0025431ab6e123bdfc19570302d60db72514ddda8b0b7250a0317438a64295d4de706047ca257d55488c9d40cdadd867d21d6c5d0799527cfcda858d205713306927eb66366a1a2699;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac1e3a713324f05561ed17ab70a99a28a1af39c8ef695e4e54c25fa55a9db7dfdb1e32e3290b4df58fb4ca9384b6388f99edb30adeae027d12644676b10b1a4c53e1c14de00ad5cc841b560e3e9f8ea9a172bcc7ed7c2387a07bb2450cd98653cbd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab78ec979f9e40c39c319ef509184517508529a81f5a9a80b2fad6dab905512573d5fde55235de91429b5e1e12550ec23c94d2c969f183b164b527d24170ce497d7ee77b15bb08f69c0a617b30c3692dee39e479fb4512550e07a641d71a9b102b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c2b92fae3242136aa6ff2dcf099ef5d2caf81774a71410c1ec6c5e4dd492c3e6d2077a4e39082cb26f6e7603e6de0e6a95d1104de49e5a9eefe884e802b102fe7fdc5ec46c49ef4f0afe8e7ed7e39959233f25514b9cd7d0b83d5416499111f68a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53c263b478f2c165be9950b3cc4747bd35aae374412730f62b03f06235fcadfc541790f7721bf2be2a48c5ebcaa7e102f66ce9d9c61922fc1cf847e42e31181ca9767e29432cd2875dd86d58b99a6121d175723c48319a7d3761cead6c52317d0075;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h536c9fbaa80ab7a534b8b18733fb72b78c04495be30c93a5c41b7b9943913d9c1c0c138e4ac1f44db8839368c44fd03b6c6d02ed46ea3f84d78804d6e48d026fff325514e89395a1b391a180ab85ed649f2859ebd7658ac162732d3ed9a0ec87fd57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h744113041797afc0eda3d1c5472db636028ac1055e279592a305a49292eca69d7fd62b18c8c76b192907c5dd0c690f1b2de57e6ef5317da238328ea521feca5ae38b35f42673cc434e3912ab51786243e29dc039dffadd6f3eac2638a7c072eb9aa9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3515bcf11d65d27ecdc6ab277f78999db19d5853fc8035ecad2e7a61e153b8cec5ad17e85ab6d7e6ea77adcfb2cab85cbf5b03c398a109faccbcf08c2eaff1f32fc2b1bfe982bfe269875adcc0299800dc41a409ec0c852584c197a1bd497e9c886;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbceb99b202a67770011cf4d8556e0caa753b4cf05318fabeff61776efc7f8c6c4f291eb5d3dada5868969ff01fcb990c5fa13a27e899f8c51fbc4ed8568014f38bbaf8e3176e1f9173768ab84769b74b9ded27a69a6f475e842748eaf1bc24eac03d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82fa2e5f1684bccbe6916ad4b6a3d6eed9dddeb51fd71e2fd1dbe37eb1e56c98f591a2feeebbe506748b2dfb0c18ec94f5c50bd6771a39d026fef59b586e18db8f534e674799c1c38277e3136107a069455b9ac3bfee0640fb28cbaf903feca7d715;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha17fde11ea888c259a1ffe49eb601868d75ccccea6d1f6f854f32a166eff9d082973c69a5d698106e25a889448fdfe5b03a7a1e8d09a6727f1e8e35f8d232e46e498ca43837d5bf30ee403c37a08ab5dd9b5fe4dfc3dca02c7e5b9c716333003d351;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h988612ed1f9ebb3cb85a33b4a7354b7445fb7f4f3fbf9a856fd95b6a516ac82baf396df7da99e49cad49fc13064d0b70edc353fbc4be37ebec7af2a33e1f9dc72ded53abceb7f0eab6b51beede95f5c1fc126fa131362302324dfc1b45dab011316a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17b4015326f4d0d00d448fe1ffb95c9aaddde8e5278f2ac71828e3026f18fd3ddd74296c85334ec4a01f8a72163300f872d5e050d32a4ecac0952ef1afbd2afe569e366221e4481efcbc87950820b400c02745d2e50365e2cbb1acd442bb6ae9620e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde99ecf3e7c74a0505e74c4c9812127dfd0ff3d3c6a340e2e994cf0f635721c955ee4b79e0f6f60fe6fd78e7e22ac28dd900e677d1ff1a0a1cdae6fba18b5ef2bd1d66312e79ba5b019d59c82b01f1b416b32af586fb38a83edcb8c029c834a77394;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd53592ee5948ab447c4f6d09587cf7b22aaaa784f603d0cd161989578e3b95cc3855448c04cb951ebec04742f33ed457a0634afeb400cfacdfa70b5a257ce8471dc2ca6c6fd277ee68ddc6f1b5d0750aad0198d30390b57d103eb63ab72dbe557a8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19f11b97c441316bf2a2c56956eb872de7b032e4f2359bdeb55e2f35cbf798f32dd4f2a22a6caee46426312de10b153dfae6a37db2604afaf31672d755d52c5c3f71225e189b2da61826492c5da1e10f784e74f57b7c443df82d676a760215daf29e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf93283a06743661c38455421f1c3c3d1d8e771eec0e262bd2f9e990fd109f366027a66cb060c8c7c47785d20b25ac189c2d32093e590f34ea34dc6f780898b304dcd5ffdc5ea7497f0a7acce0a557b8ac6d6d73d42e3341f3c9c6cc3d6c7fdb21f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6450cebacb167b7c34dbd7ff211255185303c09f88d60a26c5efbb4b902895c54e76af57589b3c9d8f653aaf860358f102b0917b196a744a1a16f5f4899a1e85c49a2c5ea0de17eb8cabf32cdc8bbbd21bb43d130fb6b3408b66c72378f84f5963a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ef015cbf11c29c461e1b58da9e2761f7d6d4972d128a0cf0c13544c9b56ba04a608dc77e4497aeea9edd0242aa5e3117a280feb12f27a344f23f0891179cf9a1a4e8232ed0efe4d468cd9e509db971bf8882e8e7e506879bfcd554dc9584d70f56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7419adb3670b858d6f1c40aad054281a614742083bf5b120e7b48b644d79dced6114f5ae03509f3c7c5ac4f7515ad5c07210dde9de59df8b97752e248cedef467cea37cb5cc41baaf1737e3072a691e91a64c9ab4500b654b405278a2255b1693441;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ffa7cfe3d92dcb8c617d9a8147baf9271dbf0c86fe8fe0b962a2ae88b762145f765011ef518cdf3290f3aa51cce9813ff85ceb56f52e489984d9d72dabe5c3e628c54bca1913090018ec2b8c58375dc59dbea31057ac629bac90aedefdbf07a3c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fdcd6ea031aee2f026ccdbb41ae908e87bfbf2abdaab52c108cb38b2e4a11fc44ae6217e870f8f871c720a6fe8b00a85fa36c4bb892fa121b854ab7746eb0d60fad7092a688cc5ce3d4e788923d2016a2d77ec0c3ee7226a7554d278114788ec130;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2089f6934a521a70dc6eba6505207489a744e4e14346e3fa67c4373cda5138282c4dc415af90e53387aeee3b463317ddb3b1aa665890c41f83d6319be5a891eec6e79c938648d9693c8c5be42c632172300da0d480293315d0e50c34ec8f99639f07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3222405606078043ed5efe94ec1cab0a2ac82c6e4c1e991061e71623c1fcf4a42e996a73d1e13f8e61c6c3031c8c358625a922d4f06fe81355d3d7b615cd8e5bf8179d81183ae53139ed150f707ce6693434491e730c957b0d279dcc9a3e3b692;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f5dc98f94e5ab7d7590b3f3de4aa9ca0986f407929feb45aad41cb019f4c8fba1acc423c948a5dbbf0e04f7b96a44fc26d0a6d439f612008153b0dfdafc15322aa17ec22944ac9f9ad1d042adf39d79f978dbc885bd16e296e5a5ba70ff16c5d98b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f59250552d73501150c1d6e132c1a97614864612533f7690446a5254a860b9fa65ac6a659d31244ec2375b8430684ead7c83e8787bf13061c8ab84ec95bf5a72b7c7b6d81751aa8500fd39f3cc4cc4c524083662206bcc02482468caea5e50600d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h124339a98e869c0b1da457cee8546948f33f915984b0428050d502161c53ba7021b04a1e7744ca1d7f05cfcd090cc753359aae3555c08baee1f5b0088c2e0cb4de0d38baf2538ef5b1a3f4a0f231a16b245494822e0d85462ff5356358c546848b7d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h115e6bb1baffa49616288c0d9996311d997f4b8f9b48d8f5552ea50c22ec3765168a4f5609e8227243710d2d3d5719cec0e68c99698c60f33ae4492d884c22940d230c49fcfadb6cec43047102dd9913b9de4ec2d4462c6a82f1d3ea28418514bb88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbe9ec82e4e16219f32a110b8bbf442ebeb89ba8af554ed704279616afacd4aa86948f2cdb56f06e115a7c7b8348c62d684be9551e8c3389bc19145c768e89d4e3e2328c00b5ea9e4fa7f1e736e29a70db44d4bfd307e7091a00b69c1bc0a4a06d67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5a54e223cc4eeb1411c4d283b159e9904a3eaf3ba26b9e83c1b8cd5d7c70235eadc719650c58a0097a3fabf082b20dcb5fe0ecbd194e215eb86a3bece5b062853ac3b355bf6681117ca4f1463cd4770b6e68461cf58e5caba2bf0b3d42c2d75404;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1fa4c310a949ee40edc0bab79119cc7e7a95f0460d070cd2a08159a0cc27362271f3cf406b1a5c91feefe906eeb413c731e8fe139655cb6fd7e6faa7511a9bfadf6ba83f9ee9415b1ad9352921ea0e643d651d98b322d87490e2919d6ea577d8503;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19bc2065a62d3f0e85c5c02dc3d42a66d10b9707522844a13c9599b966b078bf67e47d457f839f0e5f0dc0f7a81e0e032421d7ae2682b244dc98f50d2f4042b3bbfc63f906ddea3e23edbba465aff440a9ceb59de8ea8d0fd39bc544ed16ecee448d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab18f42c88bbd002b28aa13a0e48c46049d0ccdb132c66c60423c3d4b1650f2bbfa9b1aa36b435865c6cb5e975cb0ca045dbaea41deaac4d442b9d1670505810c174cac6d8283f1755cf3337a20af70091197e3a6f4fab332edc73b079855f92aa87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc46555a1e869c6b735e455cd80e7178d62fb4534166a42b38054b4771be747fd4810038a28a677fdb3131bf1447a2131c556bb8f223e9bb5fb27901deebc5d0f67b52a14df42674fefae66d6c46f35f3c9dd8da652c50d66102860e49194df45b491;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he958a176da240ea042061eefc4cfec3d32f3fdc036a2a10fbb3c8ea8e3ba8aa75b2e0e856a99de1ef26fee665a631d0fab100010e26f8515572420a4d7f48ae7edb608a2728878af55d106d13df502c1f7269928a99fd9654d98f7f34ebd87e1bb2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedb081fe1a9429a5923cb7b5861732170f5c876d2f2bd7a432acc1420ce1a83f2da3feac4a5ada3a5385d7e583069d1fd7b44b816d788a05255a3eba23e59581f8371cc27282471060ea2de93dcc2c1dbcbe04d6b8e9d06cca254ef97a0ead210908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ca563e342d81e2bf448ba15d968cabced83f7975b9ed13b3c568b81699cf23be7430bd83b86ec120a8dcd5b83c2150e8e708df818274408cec75b35d1c9452180a330fff9c2291611c757b4e56924965a9f06068a3c8aa00e0264bcce0f6fd29721;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he55a5aef6ca4f804ebc9ab373b3897ee2a0ef3968c426f21b6c3dc861b6e76273d1c7a177d1fed5652a008b2f4d9ee1659a3f3a8feaa96025022745f9341fb1f6e4f831bf998736ce062df5cf24740c5b8873b5c49ef76b27f54dec960b2030b862b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h308e3ebc0662f71cb5e500b5208044d18ae2374beff335a5387cc65eab9c556652f789975b8fa39048b7f4b308986a6bc5253806f818e387df69a626c4af540bf556d0f6d70b335e5389b0727bca9063475ba10fb5df9282417396df16a2a6e7694a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e25d4d28e88f4e1dafbf3e3c17386fb4dbe195761084d7adff3b5fb83259595dd00bd9eea14d51331545dd95889dfe206b5435f5c255368ad62ffe5e0dac64c07efa518d370bb6e8250f042d6867712f93e3a94b7834e33182637c8ef0122d4fec4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h786dc9e8e1eec71bb3b93180cadbb9b0614656281ec087c5ccebea592cfb312e45c721065e99c65d1e7a839ba28ae1feb23420ebc60cc338aa603af96fca01494d99e9e9fa2129ccc6c920a4c2eb5b09caee67ecdc9aea4b5cbb0565a64164f75754;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc16100d3a1bef3dcb6d2f6a47a5268eb6ce4a91f6c784a994ff7e54a597eaf2ccf0bd0211dc20c75a40e875bef98ef8a9891e83bb24d62cc3a1b32d1749cdedb8958f75921917e32fa3c4cb7ca2dce8f830cb43bfec7538d337bf3d146d84e1e0a44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b8537b0859746933753c878566a9a5dc2c42269344e50b374df7f36c516a7c2996d94234240acf1b42237a5e5729d6d055dad405398c988cb5d94a274faae7b4df3349b515b9ea858022548586ea2bbb520a9954380b80e95bf044a916b218c4654;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7ec3e44a60e16a6b324b719d4d8a8456b76e4f81bc4d7a2f7755875a937521ae8566af3b8601b07d024281ecdd0eb90458057b52536d41bd8de6c74b8943d3fd96fffe2b9d534977a4582c150a6ebe2718bdb9a678055c9b110d80f3a1c8297679;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d5e5e1df1a4dab086190699b559d3f69f28eb2f5f89a4728f2af0878e7cd60373cb9d57981bbb29a4eaa85ec883a1c6ccd97b04a61665a126a5954afdfe7e03dde1b73333b7962439c0dc063af72ef460e4db94a96db5c33a33d46595cdc56d14d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19592999543742352b1f17560fd23340b05e4df4f02b334f283b8003e1529d8ca3d07455f8323195a4a85627d675270d683539ac2a47ec2a67277ae09e206d99e842dbdae6f669f68930df4646a986596341e75c744382bcf3c4857c005029a06e16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc14b9ab925bc32082b655f89ca938b9cc66521cc841e81c93e1e947dad7e427549f5a4e2dff83e23e684e1109a273fa8c3680fe720bfb6fc98f72d66fcebafe20139599e8e274b296eaf97a65f26a5dce8e263b83bff532eda4f257780ceb0739af4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha084bcda7244ec1dc294e591df4a7495fc592e79e4cc66a441b3094eb2aef2f7a899f14af3f986deb04b403e25514d938f89163bbeb48cafc97dabb1dab51ba80ae907fa285f891c07a4f7921a5dc80c8482be8ef195547785f5f0556353f9f4ea0f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8bc9ee0c2ec58f129d9f07645b58a1dde6a256bba726ae353db7f22dda06a1ce4afa4cda5a0c85a385aad837e7db4901ba6d3752972a002ac84d964f698b7bd047ea692977f78bcd0af9ffb8b022bbf682eeaafd1fbdca9e7565588f0f344312bf7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d888f0d887cd263541a50f133b3a26d598dc580e2c91ef28b2768a9a238a84c46adfdd8dcf303d99e886ef05595fb37fa72de689cc1984ba2f45f782c97d17a05bfb3453f37a9c35f0cb7744a229dc1f68fc65dd1912d4495897e374ec3039c6caa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fbd7af7f968c4811d1edf2eadf255ac1b162d48791f6c7e2466348e2adb33877bd7754b3b3af0a39477bb13daf65de576e7bbe62b7c19afeef23346984c7c9823da951699e1d4f5d54bf2dba5d7b4b3273a341d5577b39584ccc2ec81f71841fd56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbea5af9207840347bf2ded3ef49b528b5cfc6d783e6cd3423d98c8f9904cf2eb8e8481f0705ceb644802cd3c0d5934796b3b649cfd03b592a42b5755fe2a76360afc2e71972ccfdcca867c408c8584eed2759259660180db95e9c9816587adf3ad18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3df077102e510a07821e9b02707f5a54299ef801426de2fb70960aeb48c73a746bc71d1f64fe2e79f86e08c1d4afc80f308f89ff18816fdd5b80e74cc8b807892af77ef4e159660ba834dfc379724edc954e88f1422f40ebb175dff4c96ee9398a69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h256550889a2ff69439b0d8ba857ebf6b63c96217e4fa7c82757abcb304edaea3cfd201894b7740e161011eefe20696916f24699a58f65d441f82c2807262bf9d04e6d8c69c0ec09281554731b7fc3b0e4146d4b96eda17d9cd4d7e802e3622457691;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32508f462b4644dc8512d4a9e68b623cd6f876ebdd1484895245e9b28ff11256d6644ced9bf0cf8aa0620eba9a197cae721f5cf98d3c37d08d62bc02081b60dff381205b8361b3e4a16d0358c7784e9a2c5d0cc28656fcb9364fa85b0097959ae036;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5600fcf1c998e39238cceccc27f38dc60dd126529260ac7f39f837be80fee63d8625ef8db6474619232ae0bef97e8294bf6f226ef738eab0575d139d5b3de848adf7612a3ee01673a406cca9aad2e49fe76efb4d026dfa990bd05334bbbeca022e3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf775174554c39b03b82bcbfd205272e0e154c91844d9c16c91768fdc9c2b1da76899fdc41fc098794fc831766f947532954d1f21358470b0127b81c154e6592d7f810dffcbd2cb43357cab077b44e6e0e069dfd441cad7607fc579a22361cb798b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3f0d65ead8faabf9cd85bca1b30174def3d1e4bd4e169b83861ef96315493d5ac9e5a5c91aaaeb61c355a148f73f3fb4b71bb0712f4b586ec0a8192483fbd5ebb5284d3438dd12de1ee9e1bf35deb13401fe3383573995255c4e574a8aa4fd753c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha24f1756698b21196738f5b3542d8d4014c5c7965fe037f0ae396326893c74bc0e889f20779549f84d5f82482d61a86ce11fd201e918e06a136a0adc2c15a883114873fb69aa4ce457e87c311545987b49678cf865239b8b2737ac216f6f1cbdc316;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d4a99b0563de32279a69ffb225929e4332dbb5009b1e2476de8fba71c1d956520efe2298804f086a5a11c00d6626eedfbe2346596ba3c49a26568f6842026255bf02e2fdb7c58c12ceb123008834e269d9a9ee4f4d6ccfe06ac96251d2011485141;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8a24f32282e1a6746684993ce4774f293893a04f488e9cb127f578859d8501568e62258f7bf8f2ad75f4328a0c2bf827a831f794b9b0ba55e8e4cc450057458d1b3e4ebe15e58acd586ad4a0296d665372449be372ccf239c44ec0fb13a69ede298;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3abaa1f2c5f3dff042598e03a72397b2effcfcda6a5f2c3533a209342e3fcc29fbad0d0359615017289a2e49dc4cd9b4e4f5962dc9b490776953797ec4ac083bd135f768229c850f2c871ebebdc635fd497dcf4e9d842230950f12f3f392d177be75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb412fe8eb7ba41790c0fe9428f2cef5befa4bd3eac503bb979afa947f15c18db0db34ecf06b0b66be7486c7633dcbf3bfc5a9c92c644beb68e97588418677ede6e0122c4aac7b66be0522649789ee6dcedd3cc93ae80c0a4097ef63679288f61e1a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7d7e1aeb6d834a5e5e2b494d040535e615fa2d65d99230efbcdd6199a56d64bd8dfa2945d8d4e82187e4708bf7805c21407f04eb7e7339e1b2bf619614bd62dd4f202f20d098e074006d26db94fb557f71b12ff0b538a074e2d6b76c96693a9c93a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h539609e9fac3db3835436e95b1ce36b25c0a3fed6c16783af28c623ffeda4072598a407ce2e379b66b71498eb906b009b7b8438a1db1f8f992e033c28d712d269aeadd36265b78cba1f18392bb963605c3182d4143db66a6d0a025675fc0acf1606d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5116ab8ccb9854a83974b1542c349715a06b673c27a0ed2922ca894153623d89975c52b415751e7decaee75835c31d7f0e00259daede0555a8bb80b6725c55b77255393b6cb6e1e997bf1273e36ed2ae6c66334f5248f23998c566df23d5cbe8daa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19dfac63873e53ba2b1a7c0c8b963d676f6e4d8b8f8a30eb6fe76fd7b4497041bdbc6abc9f0acba87a6b3e131fd1e44a5d967e0fdfc89d014912fe8b4be1d9903b76a766a317c5de6e05c6eaff8378e301a6839971c4d2aea37ffa405daf70577dc4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcad8728a45870c3d2744cfcc8a6a71ae7b321622be9e4772cb406e08d0aae6ebc5cb8d9502523eba4ef831a8a7de15f5e7e52c4f22d8dd36c90c9ff254fd1ae1d932d5c00fb495721f66cdff28cb85a9404801ebf0a9e3a6dc85e5d75bd42ca5e401;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h112a9ab4b00ecf2537324493c435fc80b3526071311a7c92660b812ab38d9c604170ab4a7295dba1eb655f0630a141974d4551a5f80060a4a978e84fe7e299f90bf1c154986c877adeb66c4bdd0616e364c5b9cdaf7f91c9cdba1495aecbda6fb164;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84c0d4b6851cc49a401784af86555547ee4b92d2604d648d1e77a0bdb8b4edc37554b869a2684d8eb141779339c2b5345f9e8175bd31ec35e511e91700e120f6d44bf0c56a8811e519ccc50dd033eae2e25931346f0af8440ca5104f26c6238747c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36a83be5c941faa2e612402c0fdaeba3b63fed11d275974e1251ac4a73eeadeb0f2f714f6fd1e6c959b5003eef4b1a8d8c7f8a82943d985f4872658bf45e09d9b6ca4c3442774498cb1353e35e30bd7ea6c535e6196db10e82ab5d3614ad32a9c4ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb85bb7eb6612885548b04272ba6aa235c35c4e762ca6450cc9271e7097615e5102e43b9511af2d1c8fbab0338e30fe31b337524c285e2645b9b8d2dd960b84692a25a136d65f9ef3c7d5a584940c34235f3a8449b760e4bb4d1d4b96afa719037fcc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha817d19fad8bcbdcd515c535fac06be42824473ad01e7ae3dabfa80a8136a2cdcc72b03e90d5de11bd9d838958fc455ac108aaf2460df29d5cb3dd63360f47861ceb30fa8599c16f727bb64781976a2df0b25d9a2557502f3afb7e4764520746f974;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf95ce4cba48d8ba70e716a8bf38dec17edc3600cf48186a1aee0e31b153e73c5f6aaf42f065a857581830497beb86bb46a06bf5015090a87703b84c75172147b0a3504655b908b58dd9b55772ac040a5a8a377655effabf1fa177cd5c8a99382d0b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h828c28705780d7289fb28dd4f191fe31ebfecadb3180bb94e93fb977c4bb05ebf94e0b8cad52c033f29402ebbf7dd1e4e58825e55c3a61027e234f690ca22c5ee494e67cf22ddd0fac3e246deee27f7393e5b146d3d0f562941304ff02899ddda0a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52b3a1d11847f526701762efb94eb75c35a7640c3884467c163863bd6611373599b371f134ec77b570bfd71d128360b00b5642a4bd999d1d95fbd21fbea7762ddf5b7a6c4a7325dde86d35fe9cae1dcbbdc6f5d798bfcc63a7b4d07a6f9cd75f6365;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70f92d73a9d8b72b6c1239bd92e05189ebef97bcb86ba9aaa0c6632a087e4b6cd730c4a6bdd2054a7e972200c84dbc8f97064b173f471453244244275743dec52b216779adedac3b1f8ac57b3617d82eeeae4067627a2d036a7830780da91d30f52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbed0c558cc44f0445f5c51fd95f7d8c6c0a266206a4195e1be2c935065105b65f924f4472a0e6e1ef3ea73e9457d8bce51833e3ca507d4596b42c0a9a536cd78eccaea6439621ef9bf3138623983b0b88932c6fe3dc00925e84686d26faf7345f07f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b5b6aa832b42feea782708743564031a74963eb5af01f973165bb68c096ba57b4c139a4f5da91ff6c4684fbf7b2de2983036044be8d87e6734519c7d0d3ad44d7257f126143b6a12ac13ad90136ff93087acf3ca2425bcbc90576a6cb359aecc050;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h414073807a76f5716fff63055363e381bcd74c4d5f24301ac168e03c4c57d34c0117e0879e8ca4f6a91384d81092700d778ad262f090fe8a0cd17a8b57a269c194c8d6815aa7e80d0e7708420cec63b2640ef8354e9fef8d988dc676e237b94bfaec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h567c2e0beb3c29298cd65a9c4cf5c458607adad93401882b7666625bff76fce499ec7b951db24a611f8e29752eeb0eb88a232853c76387f2d7fc03278dda2b28dc259b8947b746446451053d1ee0032a870df4962f50d558c23553d8cc00cbc1cad2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h247ff4e9c8226b61fdd9f1da2248e396c2ca90021a7f1345da85e56c4bc61086f482b7396e25e6e77f49519c81da1d4eb1c3f71c2cb712b68fda1124f58970d575913448eb47a0d69f405a39a852fffe1c535c3afb5d8c8072c078ed91cf53be3ab4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9aabe890f0da0aee3277acee1d20ab38c6365bb04fa4eda94632ac26f15467bf6c854e48b2c8878a45a32b3c885537d926892762a41e99862cb91fa9c03422c8ff5d1d13691f311df35791b2d1389d52dcc67e0564094dc907cd2b319ea2f1b54973;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1430e593e229e6afd610173de8e9144449ee008efa44101188cdcec57e69fbbd686bc6c2cc99817fe5c455380bff51ad7e894b83c073762fbe9aab18d27771b7175e6072a2b2b9362114a8f428fac15850a297c45ae3d5a095e622e90761ddbf2b2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h853a10ab9bbb059e90708bc7a2af068822013582dde04377f0d2c42dcd2481fd49347bb0c200e4e518f00d6f43eca8aa38df98482361c22f0bc55c1e6ed92bf0dd67485bf466397c6f2b7b436736c734e3fcdfa012dbf6488d0da401d73bc4080d13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44f65ff7ca2fbac7409b0ed2b4f20220b78fd519dffca01ca693ad87beea85601e4cc10f01709e72f6f9214bd34f18b753e0e40f7f96c285ee10d422c55dc1fdb8d81c909c105d4b56552e6b0102406dce2262a8e52acbcd38a3d32c94e8d4d83ba8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1bfd64c00a20cd38739c1db4b504478d5081c82e2b11e31ea4bcd01f93c929c2b4df9ce9a43b5b9e4076b2ed5bb702c10427591cff47de88077636754b8c16ba658f9120504a3a3fe27b24c5dc4244fe242bf48315e6219a145ac8265cca4415fb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5da7ebe599a191c7d7c9160d9951d16ea55a5b5010dcea5b45c971253f12456efdce8e10d20f945e86dc04a70d83eea94b1169e52fa43ce2a99f4224137837156e8ffa09496e99c2306c173e14e41b8dbb6fa955304fc0d50793ada79c9fc2c2d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec319a0673d311bdcbd879738dd4c14e8022b1e160f67ebf14a8efcdeeb0d55b9cc3b7b3e07ae512b7e512ead135798e337da67cc2e8520ed895f9b02d25a36ef9bcf2ee56a4c442c9af316018bbe34289bc354c5941d21717c2ec64010993acda5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45ac71841be66bab2b09af0a65c51452796e5fc6bbaca499b6d4168fc01d29f4e990b988776fe7e0da175d17dce7df251c823ca0f8d5c28106caf5e10169a1a297a424f9a364ebc1dfc0a44fd030b5782d3ffab4ba63d5983662ad11c05504ccba94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c8a8ade4f0736dee6a98b776a78fbdc6ed0d4f2b6fcc3101d4d68ee1ab2a7e6a759c2e27a76fa6cf3909046433bd3979a4fe40b43fb89f99b0d9b3f39159a0bd367d74eb5e4376e1c409037f9a0d6458f8a51332809defb9d6718ae8e6bb7035107;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb65148bbaed7bc3fef68db06179660ef4ac94f8d0be42a227ac9757ccda39f5d80b7b0a9857cb1a8f809b98a18a2080ec01bb493ab03b77761db87256cc732fdde2eaf67995f30da845d31a5f92fecc6ac4f2c4b777758ea4b9ae6a96fb29fc6b618;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc96d6f5df9700ee7101136981de08bd1a881a99dc94196756a7507869fd11f5b3603e06b1a14b71f08ebfa3148b5a3941f633177ed4d59c1ec99de4ba838f9f4a41985f32cfee72b134f9aaa6f37ecb5e7fe1a454292bf1e928af369d07c5e38c7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3de359fe7beeba9d800eee8d873c260f5a7a0ae76c5a2d1d7ad6f0e603aafb8895906bfd00492086e3c5ae581d67c46ad081d76879266fc9109be60c18c149029d69142a3f5ddd59b61d8535983a0edb3baf39558b40391c8aa99d27811f8f359f4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a852720038d22f9433c52f352687f712176190a11fb46a09d0a68aae0f961e4f94659782a985c591f65424ba11e5b604e3298c16d9be72bdd9db942d7014646fbb89faf1a23e6ce912727d9c42858f486058cba500e3362bca43894f07401ad181c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c07c1c62330b8e6e34d16341a67d5b1fc7bbe35090ea1c4aa063b645367ababd17bb9951a14e4e423e3140648a551905eabe840dc6f58f157e99c5f0c92a3c0bb1ae1420cbf9796c4abf9f9b5f6e3262e30167b67d0ff86a6512dfdac055d20d45e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h919aada4cbec8b105194f19c3e916fc2100390f5bd668bbcb945e1d56a31ee6dacd9884c789287083b4de9bbc0f462fb92eceb80820eae5880988943bd2a6b6c63ac1c4df25fbea783316560ade7d50190e0012de75a5161a2cd531c2ae84eb6de1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfd435b905f2c9b6beedd7129064a4f022bc73a46e0d0f8e41961cdca5cc1a0d51f10008dc942057bd17e775dbc5455fa2c54ec5083b00997a6112510a7430d99b1cf3005f16432636ac90303ffc217b72f20446c6a808c08fee20bc285d722ade42;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ba7e6d179bd0c17ed9f07b5cbf8196a5202cb3b7bbb8340785a9d8a7e05900d742f6aeba8304a5f2330e7f16295893906390933b6410dcc656a63e1b1c569ffcb62855068bef75e3f311832ff439a635904872bb0eef0a1210ebf029d4862ddcd33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4883e490da63743d0c367a27e7bafd8d067b18e1b238e2c92e7d1ea5d07a62bc269de56adece0801a7454d6a23edf18b2c111a22d1cf8a682488575d400e55121c7fd3c3edff2a8ad7aabe5f2b537989235484fc8f79ef9ff3f1293ab52a648699f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2215de2e4c4739517ff9043f6b7ad48b930bfc9eab09f94aaa6556159bef158bf2a9c06683be33c9092a494d661ce469fc5e07aa1211573cf9453f1c9669ebb2c25acb0957e170d98d3bb044d496eb06bacc89bfff3036161039d600f66a517ebec2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3f90a09bec223183821b274f065ae167ee8957a5124adcc9f6d769cd2f847fd89f7eb862fad8ad68b5f587256e1d0d89aa4b3b75fea5d14400d803de550db10f3e299332144d2395bf787b2069cda32619c76ad9afb6442112a4852ef93d9c9aa76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf02e261694130bf18cb0f336e601478739f80f3cd9ac398d395400359db19bae58edac4efc9058e37efdbc3879fc929e7a3e7f4d6a88f8c8297fc12ca559faeb5c668e6adaef835483393fed10d2589c574c2bafe7e710285459f778f564f17c10d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd35e5ea6af950229ecbfbe0c212ac9dee1d6f054efeea3a3858e8c3c17517e68d012469733c37d9f7db0834477f7b43c28d930dfe6b68fda2a47ec30df5622ef501c114c903cd675efbcdd7c56680ef85efe9179945d9531f531b9213aaeb8c601b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0b7efcf40dc097706c879a8a4766ded056d16f6553af2cc6b5a1c6b51515e55b02d59e57db0a7f8ae995845dd6a66758364240f591747dff36dcd4e4199da68a63184e667ab3aaa83e5562fdae2c080d5094adc46560216dbdcf3d4d99186876662;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habc643e388c10787e996e21598c9e5c3bd4f61c10070d8dea360fd4fcb6807cb6afb0051c8bb78f6c62690f2cd6d98d1a70eb7a00d80e4f70037f11bb470ad36a8e2f7d418d33918065633da3f4d3379b561c734b401d1bf0fa7dc84e9bdd41b4636;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdee72c62bd502b19ac05b2e29c0e6ca146c370dc7996ee3308cbfd9da9478b67e04391c667127eb358c85637e1950470b9fd52eac2847877b47a587bff0198ae505f84841005b48b4e804130a65d2c83fffb29b12daec223e18a6eca71be390f99b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddf51c7ffde9037fdbf1e787496be4984ed7782b22d4a476351f9f5a9a2c8c9b6e129eb6f3edbb19bb63c06f34e91203538c0fbd1dc8ed0a93fd1d5a2a1392dce46d9fa941951524394f4213d506dd36b23153e2a619b9b0a331be5e6e95242a19db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habe92fd3f533feb2deba429f0715068d18610c688bceeadcf7fa9a39c8783ddb8cc65ddc0db9f30ecf0de1687b32c18b4baeb059f6f2b8adc57ae082bb3e934e69f1a21e4cc03535532b2ea1a30e9fd36de277d899e6646a8b4c8805b099c389f8d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c3e84d2a7649c3877c02f2fa1d053678205be5c6cbce3df763404edb0dcf008222e930ee5f374e0742f11969dd54a49f7870498aaae3cc3b6792409d392baa7d46bf9f88bcbb64041a5daa650542e03fada1958623d17f13d480a6c5e956f43a69e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b05f5c57b370fd586116a0c7ce508384909f699c99dc9aad738cddd6007a1d028cc2d4b0a835c42cbf61ac2ce49c97cde25d952b482787d70e9a61c6e18656a3e478636284967a0a073927cf260c5616ac9afe0d749f9c16db05cd188197148b55b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78177ee02b239719b84b188d2963f788f13436664ad3edadd23656da93f7498f806cf87fa91505bfd80bc9b6095cc7bb2e07dc5fed84b1d7d852da9b4e326a6468ce0f2a7b87a26b524c3fae6cfb9c6ceb699b68903508125fecf93abf6c8fb32a65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66901df3a235dcf74f45007bbd9b19ccf32bc4e8718ae9d97a25bbae2eeb99fffb7462ac65c4a0657d2ec7278a488c8ff15d0c2b84e62c6a1704076c26dcf935cdacc55ae1e79bca7106cd28fbd3b41d7f8cb24c184d79b59f8f1e0a56e6997594cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54b07efb98df30f04a685d638bbbacb61419d865b313cfcbb13f1130f492455342099efa0c8bbea60f454f617e4a9b4f8dd6a45ecfa0d6b3189363158c1d7f16397bc09e60869d8b77d084fc7ac1ab73777623ceca6aaea97bbf040ade8310c807e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12b4c366dc29326448cd4a49302dd18eb14ed50be5f2d346a4576c8bff730bf7361af41a72902d2695673b0826587454263597304d09f10a19f9174396b317263da5b5293c99927913b84cda2f60ad4bd7da276c73d109bc613f983c372c2df2b255;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdacfd7cbb83f3d392f6815ba696f747e2264a4c2f31725da2b356183da9b8ab3d8dafab3a6436c20ef2b453f3594c8156300f27c86bb1a028a9216c8b392a31628f5f854530c30b44431c36d52876ba96ff46b41a96f612a9cff75e585452ebb36b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4cda0de1dbfb92fc5f6aebffd9bdb75103aac61f03ef42c95448e335ffeaafcd0f048ad48688ff71687bac1ab032095d11dbb42c7f959df04b0786b44a1ace6b08153fc5191a2a1ff5d9fa764e4c12c719c66a01fe792ac0a6568c7488a55ca21de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25bfeb78783711de913555bda5705cef5c0d201339fca64f9511b91089712d3414ca3d2ab4050cb7a8a5362d06ab91b194d736554cecf88d41c9184e5e86143a89b94501566ccb29677719fa4abd0db486398e9c7c72253b9b831654dadc84966988;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he00f4fddb779ddac2a19bf226a681d18269717f571ffd0e7568d0de6cf47f902f560c6be36170031a389a1bd3a186362d1b5b3679e057d4d478d0b9a81aa3665eff28a1aa901d229f1ba3262c04697d8f33c60260a4393a957354feb279a573ce934;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fe2d4f734e7de0a5e13f22aa7e8515fcbf39b1554be562bc2f50493f2e77cd3a4e9c4f07f26523d558c6b53024cedca057a97da637431940ddef9ed9382f4f024472072088b959c247b2b4cc31b8c494e0d50e5bc9d68d991ad665abd2d2fae6bb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6931f935bbf5d25d842bef943c5a4aefeac724d4a2e41eef156e65fa40c29fd634a5b892d6e703268429cc26ce1016a94b1ece1fe3593991bc6fa1e89c77fe4a5a22f1bdb92dcc24ba1b57fa753d3f09051fc88247cffa9e68efff909a792adb9403;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6a144baa51500c1232d2cfa927263fa84a5f9630245d727a08f1405d87c5e05e1dec2002c4513edcb8b43eb81d9e20433c34a0b115e1e8eaf0d41cacdbb48bab7e5b8c9e41c3c834f5d831436f44cd58c49a0312f34d2eda4f60382693db5e97d03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf16e3b111eb07beccf9d1ea320da9297082e3788d22c093c4a7d2a91db874568643fa07618f13bdb982ed6256cd8f66d68c09f7a6f12dacd21e9151a0e5a47680398e373be38fc01e5de3bf282573f2a52d62b832a8cd6e22ea216e841862c725226;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h427d8cc6262c92f741177c61674de024a018e640dec67f1975b5cba2388455947d144ad646638601cee6d31866b172244f28c0fe401ab234f7feacae96ac7119a469612b3604021e8662a16cba5b84a1e99ef5f745d23d2f72d8fdf36c0cfd8fd5f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf2b1254d4c176e27800e03a40161857a48b94a94e2a106505ce80606e362c73686e221dd7d197de4421dd0e594efb334cf292a6788664eddbbd1fba27fb277e59216d90d8d1a21d5b6dbea0f67b0116d24cbdae869cefca17f385ffe68ecf2f5cec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96e11944e3c3a35fcb8bc906ac47ddbb2f791eafdcee34735eda99da59d9735f765ce179cb5533aca9a9edbc518aca5d86e8bc669a39e364f53f975cf9bc4ab8d4c735dcedb5ef04c80c0574436fa878461b71558e4f46596663c2d144a9b43395e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10179ed2c1be85cd80a633702a4adda12e0512abbeb0be124cc117dc643e1b3b53fae7eb693e27864768cc21f0d8f517a69499e9db2088e65d7f176f55cbff0d81d981a993503e71b2ae337b76878feb726eb827b6187e2ffd1f83e2ce0995a76a13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heed5f4711f456355e514605d8182670af65b2d20726fb05ea7b5db651dfef9cfb04a00adf4b98f2476f9119d054e23fba998ac8a841ef2fc9b4602d79dc1384266f5c80ea57d245b032df9600a54c79a68a6786686b7461cf86d7dce4a3f437a608f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5ecf335353ae9951013a77e0e5884860730d1f3fb057f270ba89202a295c78a07eddd86cc68d9cd721011f4f5646f6241f86fcbcd12d9eab09a51eb2616cf17a348af5857618e00f4f44e512585178c1be40078c59ef6cd106060d2ee71b33b195;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdac9130cb178e66bf268fcf34284c6d7306fa63e2cf61f1cf7222371089314bb48c158b890d31bf0831c7d3108152563574e5277e80cda2bb1361569559f47122b7137bd349709e4e85177b03f75dcf4ce7a59be04abe477af9bc1e128203d5e95cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44296c214675f4b78902996db3ea1621c1f5ce9594ce9da269b82fc4c6849c9fb1793b1e8e072f08de11de0ba8dd865f93f66c4f6cc3c6c10ed524ec584df2f9f374fa90815e834faa80d9c70f736ae4306ef75601a7f75dcdbde95d8823ceb3f322;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b50caac546890fce5bc69ceddb87f9f0f8bcdc6bb5627852f7f5ebdc2f1d2b9ced98007bca2502305d1a4a7c019ff95656969feee77909d1dae1216de58a89f7c2cc45382a850bcb94b0a11777cc230fe40894b0681cbeea45b18d06c4cb5861bc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd4dac1994a45c3baa9862b9e9baa3387dea8b11e2f3300812767de9c933f79ffb3199a898127b85c859b651f288bee2bd0c9ae90b7a697d3feeeab80017654abf67ec489337224554e2f1fdfe790ebcd0a7d1d2ed81a9aab6f655d17fc5df11d656;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec3dcba0a5c7b95b62b3edf4f26efcb704560b6ed14110a0a4390d994f6212ab403e9231aab7a6ea5b9ac5d93fc04c028fa268d84f36f342676a5b24946d477b8a57c16e9ec2cf10979c7463b0ac7220fe6b5445b73c07e3882bb45448cf37961995;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1f31129852fbba68886d19736f7a7fce420284271eeb070f7a2aff68043ff6c5873580008093b927dca2e1aa3360c181981917dfe67f5ff0bf95b3927c905c516411e3cb0703ee35f1bd7ecdf87868c983749676865ab243b1e3dd5b0ee1e45f352;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb61f6eb605b16992dc6746256ca7e0d66c61704393343d6d3e038f8e00f785b3256a4425969fec2d98c9e298d1f65e29ca316833f3523b94f147b164ad43dd750377eba7cb761bf8dc9bdd2a4e01171232d93da75ae9338bd226e42d1181d8b5a027;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42faa47da53223b954f7ade73fbe329cb54ae50da9308aef2167eb0178006aa8938f0efdc5e65ea62e3952115e9a494346b3d282518b44651aafbd8e7f4d9e86def6199f3cf5381318f91f6dceb6e84b0a8b80e6d2e5f73a468d149370d1360907d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae20aff48b421a04aa2a38f7d8437b857172651e54c49e9d48ba6e5c390d5f55190e004fa918dcb7101c8735954857cb3262e2c2fb72901165ce754c72af572b83834fae525188577f20dc7cae0bbc319b36aca8b94b7ab93d377ab6f71a2e7406b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h912a7454f111c2c1fa6896a425ad8547d2834f5963c555d36534bf9d4e557a4ad59cb8136ec6df1ce33e97fbf4d4fb3733d06992c0fd8e30f882b05d93a701e4d78b0ac95deb0255899eed1ac5cb166bb057b94269b08e6aa08a1af3f01160e0ca36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2c821c3c9dab83e26c7982f1ca0dfc567735303dce88d973e132cdada521d9212ccad12fe6478aa1568cd6e4e94282b9e0b8565638b57fe538413b2e24449de81a557d1bde5f6e52f69e6023a6c78336cfafd47ee2b4a01967affcb9cd27388fda9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha928a537e1ab8105b2e2cec495da7d8e3345cb5ce4176f3084b9e8d95327e0bf0d22ddca01905e30a223c07536761bc6954709ebd43726c421e103ade54451416f9d3de4ea15d4bef6d21a8700eed53d324a868f8a78a53c8a2ad4fe00d0df5cc308;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h714ab5e82d33712e75d3c7836a062668f27b0c88ae7fc5b269ae6a8a6b456c60b51e7b9e622fefd71beffcb483e81be8295cf1f9e830456f1926ec16124f31d8d0fa309ac79e5ae82c50c51af8752964fb056834b654d6d69c37d7cb37069e94a964;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf15c11da59cbe98c1a862d09953fd2a07d2b7d716e1733ff0813bbe2f9cfd9c00229866f5bad9769dce55e42717bedc1449334b6d8be47b466d40e2d8dd9e4b357a2ddc80e140590f772e3b689f1d9773164ac9f1e915d611adecc187cefe73c801e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haaac0baf70f79ee3b7743406b499fd57caaeffa4e0ebd0fd731df87081eabca23b9a3d61b7ad137d7f12404f2709f7a95a41af60a5e7fb9fb864221abe6ba423be373d9c9577afd8330b709982a2a44965c4cce8af7b6b3e7d716a54fb57b64c112a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43c6aaa231f9e3b27be3944cdebe6800544ea2aacea367feb4a5e13d8883eb293a0b099ed50d81f35d68846aec3ef8f459f43f40cf8ae338f2591b2500204b8aadb602e778a64db08dc98c56360a59cf1d9cb91428a470f27a8d158f77a9e571da91;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha13e5420ae0a47e649e5729ee091074d9ac908cbf812181862eaa5b69954275f212dd2ddd7fcd271377bb9b267cfa255ecfc79de7d76e35ed46d1ad9eab98131971a70b86f8294a212fecc36d69fc7ad7f8b71e48db9af8aabbddd4181c159571238;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h122bdd5d021738cd1b15c543f1e71260a89aa451c28e9dc6b1ce2205c05008cdbe86a88c27dc299608eb7c3e55e3f7f898995c070967a16f057a69846f6a5098f51253a89eac1e1acb83f02aa5dcdcefa60c3e7d709cb29917fc98c491e557cc77d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b84fd4eb716fd96cdda7aaaa97ef1998a45c9d67afd3144e0870c360592211a110410dd5136fb498f002b10040e4e3734de569a09e9cb3e8b6f8e598ba36feda2bc465a5ae42f1f963c64a593859c3c57395d327cde6184c8de9f0e73db6514e95d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81621ae620d3d7e458fc59a197a15ebfd6a127b6e68212ffd840e1ab63eab8ef02fab076f9000ce359ba20e4d6158e574e3f916f73a93f8d510577730041a008a69b0850fbee776f88fe5d1f6390b922376036d8f8a49044749ccb5e8c539edc3ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha82d76a1d9edcf2fff35857b020a8d5a5f7641a8017a673eb73422a76348cfbbd8f39d31b5bd5c4d5c1bb4f3bac97a8df24fcde36a7b2f95baa4fa151f153808a058f63e8eda2d8d51a0fb58877bf6d13ff63e666194477253ce67457a4d10e42d70;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd50598ac1198da959f9452f98225bda5f43be01ef8becdf628a84e8465dcc299e657bd018bf5e1cba7cfd3c478b407469d7c164291c7e8c954ae3d309dfc23ac85fe3764c441c8d46e84cab7a5521a9cf320f188e2cd240634a60acff494c65577ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h604a71317b68b756c6fbcab6a7779145918f697e512a94c8c8d9f06e3b6d0ea1a86dee9ed2a23a0d920545ba280bfbd5b0e759b1f55401ac9c272956a235490bcff9d5b169bb793c4a1fe2733e259b37310f959897cf745a05c2937b1062006e657b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69ad424b818a6ceaae2bec58b2bfdf81d083324b5181a7842fbd3474efc83120a2bff3228739dc5acf23f647bfab869bdf07df0d85c8ab7bf41f5c1243f1fcfffc3e96abd0bd742418b2ec07851875742e87cbbc53e0e4f29f3e6ba02d73207bd55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1b883e188b792c7805606985debafe5f6ba1aa10b2e5c8f43bfdd435917611a5a9cc0d445c0c759983efdf8115375f5287b75ae10ac76ea225e40cbc349a2d254c760198471587ddce76e4282a17001d7c8da03509f32fd70c6691b0faf270ca7e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7c3373c07d5994b11d4bba76a42ec6fb89d9466e8005c3c0bc8eb5b02d1de61cf007017fef47bfbebd2321fd42aafe8877030082155514aaa22dc472e1d1017e84517654c3937731f8b254c0a5a522fce71f3df8b1a517b795b53f37a369bfebe35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e9f22ca4b0516a0e5309fc37692cff1a869c062d8e5ecb3479b06f8ec58978683aae2fb85d6a8d5be83d5a889688dda7b231c40917c3cd2fae76f3d25d3aa2d031fea8d19486563693d46f782710dc3884dd64b5574b32cf99934c618d9c226c790;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha55b50905a7513d870a3e6fb57a6f96863f4c3f8acc713a7f77b9d249ad9d61f2719c2e418cf8c01386abe4e92cfefa6401b06852c26254092125f9ea599bb3c66a29badb93acab36fa303ac23c72c4009e2b465257e7b2b5f3152600e236178a745;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h694f086dd960a476e63c73301995b87ff44390c006beda6c7aa98dc491446eed37dfe74f3e323a90412c33cdbef0b482f7c36f8cdff91157f348dcbd8d5828b380261c9f6930c69e530e47621e9234328c7e3ebdd11f86126f962505cec766043ad8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb062d646d58a934bf59909253aa9dc855533f57c4e551248722ed217782e75d7a2c869f2f31bb92e2fd83ed8e2ac473136f3f174c75278df2aa9cadbee34d5934481e9059f23c20412aee41028d5ec982483729b37bc756cb5a7de3d638d8529141b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72e85876e3a4a3b189147c54aea2b68434a415a209eb64a4d8ca7a294f9ea1837edfe01ed422516e1b69b6b920fcfb7a987a15ccb0badf7804c15bc1b787a79dfb4cb6657159cda7d42faff1993620b9065f2a0c036a7d2f68e8259f1740a6ca7245;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3101349d35bcc6297f605d732b4e63b19fe168735c2f9a34128b8d32da373c7382d42eb8b07dec76c987afebccbdfeb00887166c800085645b14fc3b9f3891b64db2e528367591525e8cfc964e7b2ff50d72b329da27b633a70c53186c2377550131;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c1d6494da2eb7c5e43f2cfa236d279c70f3f34bbff4a8b2deae0703401e50f0b6f0453b1399909ab143b974d7c5e7e2590e236f32ece2f2c6d5b8dcd2a6f1ead15253cd51da181c0d94c6a81a57074711345f956cdaf784ac5e41709e4519e27bff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94bbf558de1266817a4a10433d0981482d3b7e033a4927f19e94655e883b3ce413ad8c1c0e3f7850fe6f5a62915cf836c1f2c406e2438a471e3f7654755c8b22c38c8058418cf27ecc316b89abd4d393206b09e7799cc47920d60b7c99b7f270c82b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6852cefef223641186d0c3c91f87e68d1df121957686d9d36ecbdb2433a649c2157b902a18db31116eaeff3535f6dbf07fdd838a6673687c7f29c734b48a85113f4a136949589d31792fc26c05d71572a3e37a614c8178cc8fa988556d865d7ee47;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ccc79893a6a50bc5c05277820831c4bbf6ce017c4e56a75fe4798b781668e1492dbb772b7e221396ceee33e97795a89af6bb90c0a808ec6770659be768ba3e27ca414756186e2975b90efe64b776dd49a997c70358821f96ae0b3e3fccad8863bc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac0c60a0d817f05d3057a08980e9f79fc109df4e7b08740a8b758165b0635fd4aa0918ac25c9b174302b352b7b2396b6f464bdbd625f149d5837c80b468d31ae259f653309ffc76c4dccc841b375379b9b69a001cda3c127d64e91f01b973fb9c45d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haed7ed8969bb80b3d3ccae4411e5d6794019dead530d560f3fc5759d768ed3a3c75ff5dc1ed5d646e3cba4b895adb5c534c3e5f54e240217218efa53fcc2cc36c3fe80a644932a6eebb49ab394a681bc30a2cc9205db912b245a0c5854ec5fa2f7c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0a843d4b15b66fd8dd17eb02fa5400a55fa4e6ea7aeacc4754fe4777902eb0f41b42743bf929e1b97eaf1d4ecb63b6ca11d1f10220fec34925fa2f7d1e4eeb1c700129a200294f54c757a4cf575c810a049fe947ffceaf38c95d84571774b79aa75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7321564b6c3fd4e0925895352312680a00c3d4758967b98f569ce4dcaa3ded4e49f1f5f3f9c975d9f2216c5f12b1ee1bb83ef3a87ee9279fd833a49c8c4db066c4604d7c08c1b96f3a1ef90f7e7998b461abcf42b958f30aa6b7526bdb23f9124f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h798831e1ff79aeed6577be1e6f227939e5b16e32a6a45f1bde4ca07021b99a4f8908ae3858ba46932501239636c3fe62404bff26136f7160ccb528278cefad6afe6ee0caa46cb85e97a8ad72c42e82b14f5e1382de7352335112835e6fbede5c87c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h509985b2b9ce18dfc082e4430b331db44b7dd7548677f6611799b2408ca458840176e17ab5fa1a3d6bf579d65d526e93018e6c4aebcfdba20e7d23c0ae1875c80bc9e760df3309b8d44d5780275cf53d4ffa6b277153f0f1cc71811616afe4af0a1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a341c499853139fe195c33e4468a76b50d1e7079c7340bbc3ac1fc0f2eb6d446e17c2097e0c1b934bdc32be4e0d4978f7134443e1049a82769263f1cfa64c6b191b914a789bd7d1402ec298070fdb9128ad31233faf47fd693ce12e826843cf70d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66040d317d0aca6923935b938fd34e92fbc42d7af4840b3df8ff1f34c8bba661bc4a3b7e0d2b411e8242a0b99e4b331ec6c06bb1941f9a002dddd08a2fa632f9e1a742420896af387552e4c2bbbbf17935c0985c87834a0df0d8920fbdbd81e19511;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb97664a712817ad97b4fe2ff1aeade783fda38618fd1c2b2b7a3b909a762a040edbc328930aff23f7da43d07531d4a6a55513fc86beba43be53f67ead8400111218391d1449ed1595ba285d1f4a40a9f77d58588edf1b0c04b3a365fb8a15aa0a3b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a7fea555d27aa23c75c9674f9116bc8ad4e9e4986da086958310509c98b09ee2d6fa8ec1a367514376ca6814758d5ec04253878d9e7bc6d635415a927528c13f93a4f376e89a071b3bce0de838737c485e0337836c87cb02b4ad348395100ea1da3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2cdc05d2249bde4019f9177904f21cb9a48a5b5100fe7858709fafbd53d8a5fa05359c40f618ddd39d3039ee3958800b004f2ccfd85aa220a5d54a60b7d4b7f9bd4b2054df94c1592e803734f5d581a3d82a186617fe0dba853ad29f99c24e1c305;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c8dabba6d611f69c4b59185d48d706d4a64d30fa7eff039e41adacdca5e84c80e1497e91ba1325610ebe5a3c9aedb9fbbc75d3b13cb41fd6357352f4251c770514cdd8205895702ce540741b11c70ab859189c00036b358cb49b91cd9085fef4121;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha344185d551d270259e2fcfe0e5ad8a2f7f5852d85537d621549304cb48100a883b053ed579f8be44f99196e6a330c3943093d4c95171cdbf45b7d7cc87b670e959337e18d142f84306c9cf98747dbbc33afa1eeba777055887aa773ce9da242470d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a4ebff70dcc0d10e9b11fb276529885b58d62fc1804ba02f705f1da2fa2fb95fc55244d4b97a411ac2f7e3b7b31c6e18731b8d234ebaf7f2c25e2b501f6dc95d0c204e84c9bcbd6122838cdf700c502ddc30eca2466735a388ac1ec9610b0e1438e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ecfd119aacaf42b8317a16f1558eb6bc917d2a6ce820898f0d2c303af72edad919c23b71a8d4111770ee8dbd780d127b8c1c8b558ff3198d750ff0af0de824997991b770df99efa68075f7d57653f557f85b99c4c875e5df1c2ae3a7bce9a0410c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a854fca2885cc4bd4aa4b7818ef2182ee6c111ce6b4e440077fb1dfed279151f0ac1220761293cc10f7382e0f2de74c7e73d1221d2e13a21e87dfb916c919773a5f4ed2b51b0059282ae11ccd9eadfb98f28ba62eccbbc9101cd5c0e6485d4ac5dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had8d1c9075cb12c04bddb9f3c5ca6f682fa7edfe79106ece492b1fdabd135ebda810019846543a77a3bfc1fed920ff93877e16e527d25d068980a7020a47829397131a2dadfeb6c2bde212878b195f7a86307ac0ee555194d88a1043e485f41c5c9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b636eb73325e4c766c9bd12adce230353cba69eb71d0b91dd17311c90f9eec049a953765f67d7b4971cd740fcba772356ce131b3b1103c384446d9c1d87dc5ba6570458b1203f0ab12f0bfa8a06b1751dc6404ee90f2ae6606b45d62720622bcbca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4293eaff5546e85b8f8decb559e4c2297b82b87d57c5af313a20647876b1dbb258fb4c937c13da202d0053cce628a97f4efb2d1a972a6004419e29720a271482e4cd42ccf2825ffa856bd229b7682b5f0fbab79aec92d83b52fb1ddacfb2d6ce6d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e501e987a4cd2724818b185de47b339fa61ffa3c6933e68e905a5d7fcfd77f79b30ae65b7ece167f43f607664652a74a52b42cd0416d0a8b611c8d2f0f634ed4067941b20a0a956a8136a084986beefdb636e9abee6b4dd774cd0897b8858ec24e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb96f961d4703200e8e72cc012eb4e41da087158a8a60ea6f6b5fa421da7c03a9896a6eb4089daa48baffbd931aa0d55d161b8544e05ac81f8f742edc75cfbc1bf54bf6f0468a354af2ae3281ad6d6782e7502a28177548d08e8e046016aacf34bd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4876be63e29d4bba64db08a4e6940babadf8921410b35dbab976d1260a463282a100229481f35b83cb7e4025cb068ab1838e4f49630c801e10f1939b026a21bba379be65de14b0ffc4139693031d35d12c5a53bf8862521b770e31b17c0268fa23a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f1b7112944594581f74eb17ced6f1aa4da01f7aa8f36b2861df27b62947a9bed496f5c4ea569c4fd27fb474940d0003bb618fb4f9959fc6b556945bbd6360978251ede1d9e4fa457f031059c32e746ab9a55bb2732d41f97c5a9283162cb0b10f12;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0d76f4f85a9ce6901a72ab35b6eb2403768170affa492dc53bfc205b58e0bc79b2270fe0e2121747ced220f324675b59439e90afd909972642f28f6a871718864a5e4f19ddbe6f7ebaafab0e10009eeae22ae3f70dbd4e9225dbb0330b37f03aac2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb88d61be4ffe7f2a92391ba36eec426314a6b2db81f3792673f141b4920b22d22e77a636a571c95b2121653ed72685374eb17eecaacdd7fe74ede387eec047dae922a11ca8c541496adc71b76e00fda543b7a9388f5eb218cf8279792ccb076b590d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bc9fbceb7035939b1ba483d8d64ec5421a2b9dfef272c1b4bd1178a2876aa58916b745230f7de1d2651f378e16c347354215c143063104338a5c7d73aa681bd4d3112c6841785dce2a50248011d6abe9e7aac127474a7a51eb5cdf14133ffe33c9f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1987f20343bb5f066e0767c919362c6d8def24e115cd814a346db652628a81437d74b33dc28f36ef897b3ebeb32fd798652bf5f9ae055764bfa1cb932a32ce1dd000b8fa071c28d4efb544e6afc5e63ef75993bb40f31a2f5e0192179cccab40dfb7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3eaf7e0bff4dcf21f0e41b0674b0d5f84cadf59d5fffa8e1768086e96905a8ce8181f4a8d3ecdc19999fe8c88ff01340e5e86abe1fbae167bc8eddcd637bcd295e442ae34cebc73ca78edbf77c15b34678c0790b5d389630b263bf9730a6147b0e93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4744df1c27021acc816a67930d1510b9471ccc7483d8496325b7e3bf59bd91b1511e354458afbc8db3172f59383ca5d448492af812d4a236cd1af6fd8a54f8412214b4f5f090fdfa03802c96e88dda6728e154c0ad70bb170f99c37e0a518d6a003f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7245eb50d6d82e48fd6c2f951fc5667e94d954ffbb387574f961404f57d81baae369b458b48a6fb38f4af1596ab44caab27c1dc3eb2e4c818da3c2c515bff5db1a334b153aae31b21b7015079287692a66b142d982181b2acaa9b8fc04c09b1968ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a178a33af77996ce7b832eeed5c75efd613882b428c4cf98fbd4a64278dfbde226d3f1696451cfd1954ca8c3a5cf3929e403850d161e6aaac398be40baa0f4a4a69e9206bc4553a0780c333c7461ebfb9137124c5da3f8f3df38fa06408fcb8c241;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d760bbf091eb2eb2484dd897b126c3ca9b6567453985c7fa3040a8f9ee10f2a0d022d6cf3500237742caa78069357dd2c89534a4470ccecdac1efc0daf68345f1a35a76af13ec80fa181ddb62cb47304093f391329148a3c747ea81d5d087642627;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc6eccabb32c0d883e10a2952c24fa310fd69271f142b6fa9589f3dd0ad42c8cf167228058955fb06b9c8832a67218e8ae95372786178c940e6b3408cfcdb88efd873df702ec4cfab5a6301e34954c8ea100728a8b1907232be9e3f954f3ffdd121e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77821a87d34939bec8c9299641e4c44b1572b187a07b99ad7db3e439e941f2b0976a8bf8a0f123f30e95cd533ddf2b3bd31663640ef75ff8a2223994e37128754f87cc97b428354dbe8f9b9f6f0f92407c55fa57efe9566005f7b8e30b1b3b620c33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96ec3236ad4b6a3558ec554f9b0c7ea6c10e99d8219fac43e787a1b411adfd7cdde04976b588aa76738731f8d6e12d5c40163a816c061ddb3ab6c572cf847240dadb6469362e8ddec14bdb54a08868db02f85ac14701526ff024e397b384a388ae75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e373e7e487b4776d934e03b5863224dd8b07b9d5609466e8322a723c5ebe6cd536b3d5366a90ba2c332a9f60e9ce1149d134bf2786b37d4590eaba870eb817ebc69d267921002b994e9d7fc4206e3e63a57daf0ab700911477af6d6513895f0fb35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb85e5549a90322dc0d313b8f2a2648520371d5bad3c7f61091fad52cae700bad10138d8016ff34a6df5af316f888b52558587688fc809d1971d5cec54c664ea0cdfa4255df6a1af0d219807b3d2c947b9d1eb0be302e2ecc1980a99f40063799420b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e8230f82f0fb22405b3cb030dbfb61e487b69c045c6525cbfe106ba192466c4d55b1b70a3920a822f01c14e03e66fe3aee21ce40ec2888c68cf4e90d7457b0578de72e7b5ff243de66c840f89dba925437b3be1923c69a55024920395bdc864554;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a4b78677c837693f622a47c8626a387e1a8f87b6bd8e84bdc00d5c39e6edeba2fa06dfa5a86bce0c820b828ff00d119389419be2bc73ad7be7cc3594cdad87d6db42c26c7ed0c8cd76b011cc500bf0d16dc6c8c8f67c59eead93c772234f9ac9485;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcabd974c7bd193d3183b1e1803ad44cfe47f38d0f1377759c12853c30a5579761936a51a416b633e5cd3f03c179d3cf061f75d9b9fda156a179e0d3eb61431e6880e3b5e4f1fd2eff2d0f7adace509ff78338d82d266e985d42b635431c26728f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha14eb876bbf1c5ba8bfa72f96a55bd0e037a3f9c1e5d423c1fb9cac99ae4e97f70d8d6db3e7f8d6c4d3b9d9c61bd1fed2ef16cef9bba45db5ff514b4087b7666d2ed8b8346937c19670350f419e53bd75f552a01fc6e540ba850bc98d60fecdefce8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9cd636bfe774671f073078e5fa7aca01e0be7c0a3c21710fc4761fde42e5d923dc49901414dbe768077f7b6e6b7ef86bcbbf166b59275d5f643d060da83b7641f9bd7777b98ce25b25601a59abd41fbbbd0882da496b6c694aff6d0842dd2f9aaf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha769ce1704f26574c1ff0d325280dd9b673a4e46698a98c5a1f022fffd293065dabdadfdebb71b9845892b3d3727d32276601b7cbdabc51605a41d51b568787fbd53345d2c92ccc5be9db191163e4d84a0e9b0828c30674554a436345ebf8d304724;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbec568d5645c1632c162b0ee00be411403060086d620b8e40d310e5891f5f9173efcc90caa605f45ce4924a6a46908fd6a72403a875e806596fdc735821d1988ad6a4ffe64862ad3abe38ab44b7f0cbf45abfbc89d68d4f3d859a74459dad4a6672;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa607a8430cac5a9c8049038c47bf8e3123a9615ff1ca64e779a258248951d6005b199e2344c355319f691d53506b22f822e9098f916069e5db144293397e6f1e8b0b1bd6b0a21ba75f85cd0364f16aad19a92ecec2aca548c31e2939291c8a27382;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf7f78f50bfd6e763db0f075d3ce74cad9b42a137304fb05801bfa42a37acb0aba1bc5cee40c1f3212c6762adc0b517d7711225a736510853082b30abf7bdded749ebf4f63e72e684c8516e8d623bce24d942ed54825672901dfdea5126a78be993;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he33594286a00236c3af9d74aa4d3f0bdd5f691112fba103e8cb3d405e73a0fb9a4af69b78b8fcffa771af224ea0eb1af941f978c5aa70ec70d77e547912b175b5834aa0eb920a63983ca7b90ad7b683ea888c3cc66856d3b9ca1d5a5c958e16e01e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedb3b21b8183d5ab0f076efaa026c1d020c562956f33a83930871d8058c76785fe1c4d8b9d5befc0c033a2ae43cc4347d341d4add8a8b840d0cbd011a5ee15531a9620c442ccccdd5524c8d750ad0cac3912b0cd47c8da18f676f06790eb2f605025;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa5f940486e828dca693b9fc5a60a5183949c77f41356a22780fe39a27c174c582a15f775fa05d85de64978e922f2733662a0c1905df861a5a8f0a5b9a96ef05631078e0a15f959a4d21625a5e180b1c029417860495c57cf471192a89264c356b56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4571986415dfbde0acf981e42868bac54917349f7eed69be992cc845f53d3eae3ab10f24c042460b39e89339fa7c2165db6a3027c4711483844fc2b14700a1d870b2a8f7ca41104f5d0fac6ad55b174b6f167f6de2862a20bc981f7ac20b81ee7cd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd841ba7e2c915a204758bdaad8341ca7652028c488760db38bb238db2f2718f6aa037511a12cc61be634f638d05ae40d6ac5fc2a58c8a3a960c06ad8570c9c419c9f59f3d1c152ceb266bb78145cdab1ed6ce5f4653bb75476f08c9e4fdc9c347613;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bc40cdcf38d634469479d18dfe160f5fb4ff635c642879994e6d7eda71957cebe037860005e8faba3fc23e5e0a72e2d8b233a0c9c51bbdeaa1795ffc687ecb39e8d5d190fef3359845a22b37ce0a1c1eab2af04b8ee525e9d418aba552e3b1e58ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ecd9425d64c685ec57a5daa71ecf786fc050dac5f016abe29ba95ad3e33ca5adcc961a881c6b576206051f47fc20e4b2cb6695025b900390f37ef3128d6f404ed648361f43c8f2f177796bd102c6ac381c123e82d9d4e17312fbac5d6dddb4c3a6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87de936ee1b85d90d47bc0f58e8fe3b9cc20bb639ca67d53bda750d833bbd0853896cc7f11ca41690bb8f5e97a058f0417196d7a0ef33b360c0e02af86d4d3878bae59582f357b8066aa84b9bce57f472e7bc2beab73274d7758fd17fa3dd8858b43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d2f8a2838cfb6d81522b4acf835e3bbea7ce48b7a58c6781fb1d424c23362b6adcb53c1c2fc9a4ec676d74c17b48c1d86deba91f3b76969b0d19533fa1eb0e39fdf6ff4e43a1f00ecba0d5fb752509534d826635c16e1322012803612539e6e81af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10d47149e8b9f30939a55624f6eb5e2d21e6b6a9cfadb5f956758d4babef387c28f9d5c9795478b79f8ea91724ca0ff1bbc983507321a3304eb3b8908cacc2599a95f2134c38e30128c52dcc82443b1b2c8ac881343692acef2bf394ceedab99c637;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h629913d9d9a327f8298522f69827922d56740c3875822270ab4d9781c232ed460e212457dc9f9998742e3994f4dceb41c650e9955bbe538cf89326fac01c772c2a13bf1929f5ee60f9a39c82d513cb2faf64e33fc573fbfbb2679fe0123639001738;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5ee2ef6e5d692ab34bd7f1af46e06f096df76d9ea6b56092a8c071893684fdf468780d8f8d3d994b7ff4d2bc7fb808b023a4aad4dc2a6237c25bdfa98d203515fc53d725fe3f50f8c1aeab527f4a53d9c2c000a6d22900419e0dd7eeaab75bd4934;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b148aaa344b15cd60c2ffd14d2e686d926b74652453f3764ef98d9388793a3b95ddbaf5b4073b5388863f2245f7a723942c3d46415f009acfaaf740fa33bb701a657a290462de762464c30dfcb2de2b1a471d67cdc3f7988550a120b51768751706;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7bdce6ca82a3e880847dd8c523790a69c113a2efeee178475a6b1212a20f65ead18e2f75edd269275506422961c6c1ae947c72945403b31f5849b8ec3d7715008392a6468a86b06d10278f592abb45845f058ba878b8cc4ccd994ca3e69ca52199d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77c0d1fc0f4dc45666d20bc029e90217fa6338570c2ec4b55e1817f1cfdcfffe3b322fc056483d8ef4b71d53fb42f031cf7b9de13bf3c33d067110ced681802fa74f7bb1ad7623c5e027cc3a5ef7ca82c370293ea238f8f7c92221e1181ace52a9ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h185fe86bb47733a8ce5b36593cf153d9e013da05d9a8e0fa40e5f8cff7be98bcd1e869426c51c6914006ce85e11bbc180aa4ebb51a70384903fa867fb0ebff3a85741cbd1883e21c740f198594f423696fc2e41962a06fcf3ed8a185ae14a33c71dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0ed0ba709e95989fee67d51bc161ddb2d067aa9d757c102413da9448f38c59692c2dd6539287ad5b9aae9a048ce6ad2a4d4bce9e57216d43f471d739747d1798fb9611f75606b4c1b7b84c4a75a6d86049bb5b1f02abf5aab4e34cb0f5ab077496d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0629d686db409d979877669829bcb517e094036a1ac745accde2004d9909ed3e7f1437c2fd7e715ee268f6b1f2a33cd5915d1f37ae01d3cf745bf18b6ab4901d250642c8add50a93c5cdacef1ef8df439f4c52f8d2770f67467cfa040a6ee1f794c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2a13799962e802487a58ef87bc93749c09e2162831c4f322a35cd53d88423f44a34dae67642a76a323842db9c3cbed9b7d709b8cc7dd54b15998bed14190d80b70cad704510fb4e319fbb99f14cb9476852c8cbafdf1d858e99ce965f4b29b42a8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bd5e814894cb754bdb9e50f1d2ca84cb8a450858686fe009963f6ff8a8a40c86a82928406fe6ec6f9b3408a1417541410710a54e80e14e4d68c778c7752763c66701fa0a83a18a6b9680dff844e5efca255a5008ce7d492abb403287a068f0aa4d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83a0d3d89caa1cdff22accdd19b682c53e1a0dd13491cb3c4338730cbe4685aa4a663d6a0a0ddd907fb08ed0d88f7a13e3f4e8777e2902e0b29dcdfb7b36ffbe95dfbf92710a19cf7227a4f5b13ce3a722ac28e62beeab177d79fe1dde55cfb8f4ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h638f06d5bb1848f0b976c78129338b10077d2c939145be88033675222fc63cf3c790b24fe4908ba4333e235328709368e010c100d0ca715b03ede74291680979e72be45f0d3cb36374013b27adc1b75f9b624fe0a746d5d1d0aeb9d3997dccc354ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97cd40d6dc4c6e6ee94bb4e60206fdb5784a9060630e99d58250df82838886dec8aff173cc57a691304f2735397501718433c3effc2dc4b89016df59b9bab06e6815ec732cdd4345e2d1458b071113297f3688af38b8f0afbce812df87d0a15ef410;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha94d0f4a10dc2b9a654f588ab8e710c44ed19ad4be8fc94e50631b1dd9a52b3e0353d4e4061140a6166e5a1ac35276c5727f4973501e803edd5c3786287a26586352c007d9509cd3c7a424a982ae91fb469adc3eb681376507f23d887d15f1506b7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb782a673e05c10d89c108b61b97fb759b79808b9f335837602d3346178991484830dc7174fe3e5d274398ca7fe8eaef7d2c703b318badcbd965d3fb252fc40bfe0360e8333f1b6fbd2515d093ab210ebc69e8cb4a86d2f07f4744bef1d1c0748b75b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0e0d2d05591b71efa2b69f5ff827532d9be9a638ed5e6a9bb343b4d8878c63e2d21d229306038f61084ee0fbff0b782627e01adaa422042fbe27bef00cab97c0164c973c903accb3a3ce8e13b35fa1164670ece5e8aa1ba8f07fc246cb251a1408c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h602ffa72114b739f979742951078cf9767f3262526d343fbeb23c4a982cef67c27068919b77ca38ccfd85e7f8227d55adbe9814b6ef2c0b04055be0bcc5d81cb9b3dca43a34e6966b26dbc336b64f37da0a0a197658087b23148c2d896dd956f1efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8320f913f75cb46cef531350425a7eb8e139c451e2d6ffb453a0855a4566408dd562b4ad86a7400008a1cb9b804994568757b47074b3ac54f3323818564b56789f7377f134157298542c509113ef176165739265917cd08e30deaf69ed32b944eb91;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3554851b242c50787cf1aa0dc8c1cb6483b1d1c93b555e6a52e9137c5bf47517434875b59f7c3f0e3a539920d72a9028e2a6023558c18545914257cac00bc72fb4e5d047a4277a0ae91b5d940e01923ffb9d220f765857fb513c5c11c4b8475c846;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h164ba7709fa3d420dec4dfba46b401f6a659eb41b4af729436553fca2f97af67053de895de26553c8660ab615fac2427cf041f58d89ac26e95ff28e1a2183811bb17f7a9ebbdc28cd0ecc699e96b4f28667546c5ae39702fc49088c08b949c96adf5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae6f3fa1f38fe74c4ff50e6de57f362117ed7038d5634debbacd548a90882429f6d56f69a2ea12923b7999ff375b9e6ae4d2c69fa549634470ed8a82e4793f80df51898453ff85c95905d6439157963e69d97d955ae9d0b7028c2bdb2b276d7d5ad7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bdbfcbc57e150e6f71868fc355046a8f998cd9329ea6f794f4d4da678762d405840cd593723178b63b145f0b9756c5867f92457ab4b1177d10aed8d63073168b5031bfeed65f797e838aeebbd36fe671484de225eb8f46adaaf99222b263953b575;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59293d231b50f0103a788b8626aa1996b2e8eeabbfd2f4c2bf60840eaf38bc7d2667e146a6bfdfdaddfb10200b89f8aa0c38f13034512e408f0cd7586a9c0f4a42bfca8d871e89fb3aa1890ff97362f287e682870cb8565d948186e7be26f4906829;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb3f78eea7400502fc4d3250b853ebdd31c592291f896b7eb8cfc19d95b3952f3dfd944605aa42edf01724a9847e416f5dcac71d1b86751ceb109cb60d73130bf8d1d918beb4b3cbc592ea5f85647710c5d257e0183e95d2b490bcdd3a2be0398407;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3437ab441b097b73175fa76a6f826950fe8b49b938d2d325d40cbf9325960549c5dd379e5ef7b4bbdeea35ce415872f975fefdbb98a2204923544e2364b4c8b956c565cc6382f64787099b936d81c0b22ac4bb5d6db600c68147cfb9d0e5f395b81e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f7ee0d1020080ca80318c362f7c544c9ad11818ed0c96a07f5a8541b102330f4bd752ddc6ceb68b55767d3b2747a9c48f9790a88851ec6cb6c73c4368f3b4735fd77315e7c6732c7bfdb6c053d8a42d8c8ee31ce93775fbb75f5753b75ba991e7d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bf4d8cf971121de19b8c168b79a6899e4684cffeb4b8597ba4c535d503f062f8f89889be857cc782e3f88b204af426a2267509a86e101feaa0809008d32c566eeed0fc4c37044ffeb094c8ffafb608f2bde7c6db6b7210f3b100dcad7de5b7831b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a38c8ad633f62f265ba2b897f20545a9d1a0cb67ca35b94bfc0894fe6fdce37010369afe989563b336d7d340f1af142749e14a2e2b02ada215110794667db74cb6ff210c26f083dc260502ea0c0682a9ccaa9db2e4da45afecbd90a5bca3b3701d0;
        #1
        $finish();
    end
endmodule
