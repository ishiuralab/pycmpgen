module testbench();
    reg [22:0] src0;
    reg [22:0] src1;
    reg [22:0] src2;
    reg [22:0] src3;
    reg [22:0] src4;
    reg [22:0] src5;
    reg [22:0] src6;
    reg [22:0] src7;
    reg [22:0] src8;
    reg [22:0] src9;
    reg [22:0] src10;
    reg [22:0] src11;
    reg [22:0] src12;
    reg [22:0] src13;
    reg [22:0] src14;
    reg [22:0] src15;
    reg [22:0] src16;
    reg [22:0] src17;
    reg [22:0] src18;
    reg [22:0] src19;
    reg [22:0] src20;
    reg [22:0] src21;
    reg [22:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea8d41fcc71af2cc081c37ce94f8331e3dec31115ff5c313f778db1bfff2f9cf7ccf87520299cfa733820d0979d6ff928b27b9f38e93c687f73637d7caa8219260d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he07cee7c41b7135cf495e00d14a826a958233b75647894af57789df891dcb7f28a37a2f2fe30aabc1dd55909296d49e5e71e351d28e5f209b2f43fdea443af070466;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c66bce0ec89568a94a7016080191440e324bd266a34d4ebee1e50746182da70136f806cc39f5e61c5fdb10cb97a9041eeb405801080dd8590892b6fe9e0b0da9bca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e8dc868e9a218bb57b610f7628c7eba37b8291e81017c8625a87766025dde24479bd521c67373d2ed13b2c8439f1c42a7e099d29f51a38ec468fa1cb914dafa4c04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6783aa2a403df4841b0cbc0f4b4aeb92441d56c6105e4bee47403610c761d55dca31657c0dfedbb0cd1e301306e5609f4194dc431221f5e71097a20e7407084ec5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf91197c445c2d1fffa9abd6449c0a69eee19a871b9330e2d904a19cd1c63c61f33a253ebbfd5843d420d3ca597b0ad008c551a32c307f0f8edd001bb2f3af4df5a7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1abb80b4f0acc7e5b073a0ad34b3a436d61320d492280d335b7f2376295c83b4cc46b0e6a5b48aa85d1a1fd828f4c22a544c74a5a297270254ca5018a74f577ddd74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7735e42d0512eb0303b0c3ee974dd1b596f9fe774f8a32f5eba90a3efb940fb4197c9619353ab63ab59ecf9c825cb378976df505f11689687ef66516694d2657166;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19528000bb638b4368938b5e7875d8c26a90b88e3647bf7d53ac78fa5060accca0181c4e2264c658d147bc861dcdc721ba8b1f0c1302ba4aaeaaaf8c7c9fcd8bb2d64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1f9916e60cbd14bee8501df0df88e49ba55cb98d7de296c688a02c8112a28089943b87928a1e3785c591ea7c347119b7c5bd99bb426bcf0d36b1aafb8aafce3469c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebe0e0c9c09672b9017d43c4b0ed581bb8ab221b72d9affe9be43c22af81cdcbd564559f2d2d0cfff8dfd26170a33c83960bdcafad127c7cfe223047b71c52143b04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca55691820c4fbbbcfae5ca4e2ac96973c93cc17c9001b731a8925f0f22b58667ea99ef93fd2fef3e9c6042fe48da0c6bd23604cfa8f0dab1d54356c210b4324814e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f058f28463fd939c46ee41191a746081e57f3d4203c509549650093569bda658a9b0626e9387e97dc366f210ca5413f0e016a1a2fbfe2b654ba64efb37851635cdcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144845ca8cb10e75ecf81ebd741a64d1049b7ccd39354514e0778fb71e73a0da83aa8ce91c2dd860eb1acb0f7a68052d471ff25b877a290362eb0cd2fab64bf420611;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ef605302de2e70ef9e29ff70be7249db154b9971123e22625c7ab0e9134d3ad4e000df4fca82a57d6fd1fc4eeb9fa7eab631f6b2550f99670886343e614277ef448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a6167a04ecafc5a198d2e2ec06e16f2ed3b763e4b499e588a11fc28ee6f4cfb9bbd81781298fc7f0241c8229ec4654da3669b00bd7093e9f6efe61cbdbe2ace4510;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe74989e74f5798b777f8d519acec65f63f3754453120fdd08acdf2a04d3b9c9e82f06ef01cc5dce8cab7172513c1cee34a8070c12704eadbb34e0ce2fd96f943d89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h465f2a62fd9a1f2815bfa67e4031fd6a876931ec21cd33af925c31c3cbda2b2bb92d46a5480f95e4a9a0b717c45a8d14c3126d8e8ca1765034ab9ae4dda4de650311;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c55216b1360a533d51f3422a78306aac1de308d4891a5594d31e5d138d003a78c0994f72e6ca5a7ea7ef472cecb8b107587e37394eed12100066c9aee62550af5e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18763bf730646bef02024dc8b7a5cf8f9de165e9e7a21c09a8ac9a783a2f98214921b4574cebb3f799afccfdb623c5bf616befb97461d85fa3a0917f0d9cbb15950e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56aca7ae50c11a5362553fe19ad41c771a4a5ae866c6e8ce26ec76f63ddb76f81dfb14dddae114e75670627fe93be2d10a234dc7670f2537fd4e9f491f23346f849b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fead7aa30b78b3c0b2f323ddb73949584ca1f191f622cad01956aabbcd2e402bd209109e7e849441f05917dcb0768b29c6cace8061efa975c9b4fbba0dc11e3ef3d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he788ad2129425d7427570d0284f00baea3d6f53d18e90743305baa75ebf962fd9f1e9a79fba99bfd4ba1f3030bae91ed43ca63fc5bf3813fe3a54fbe81ffb27207cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebdf54750e3b3be36e6fd723d800531ae093f078981dbacc9f1e8d5163cf12e4e36a7eee5503c6074d10d92677e3236b275cbef08d9b2541a53b91a4be8ae8e19d50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155a7752a085ba365e0c4782ffad4f87b4cfeca65bce09769fdc4d9947dbde27f8fca9adcf544492ed30ea97fd7cee4a3b8cc6b49a1ebf178f5bfaac4a185bd89c473;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc0255e76e55ad48dde0c59c215a01269de689f1529b42398e4ed3ffdf9d7dc64365fc46589b971ea8f85211f7926a66e929528a987f99ed76eeedcdc336112782fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d54621a160f22ad59a2e8641ef0124b48becd374a6728549fdf34293e0805699f82944b66a71e0f94ff48969994d6cda1a61986fa0d63a58e12f1be6a1e1fbbdac42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79b63e6a02b3dbcb503e528e76c4a4447996803575d8391d13de0adaa753519f5acf9a47fd7c8075941953d8a2b4442756e8a690c3664e8f99b01098ea943e3f9000;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5a2023e6286424d80c470ac821af2623fe6a726600f7b55fc94d69831626d22e66120043bbbc737951d0ac566767916dad4c93dd4f0258190d96eb9457146f0bd20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb193c9dee8f1001a66733f54428488cb1c371432f8060bd6bbd466a0750c9c4144e2aa947d83c1e74ba0364651e8a04429670b59a87087350cd531797bf8dd2f848d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78e91e51d38cdfec1a901462428188c5d9993ba2f56d129c92369c2e7896d980c77efbdd43ba17a4f8534f99c5d48e37c6fd453db59ebe8427d719bd2f59df375f7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb934294c4564d22f89c3685d60434e19f736b9ae4fb4acfa0908042360073f2adafa6b23894e78bb2a5495cd0b6375241d776a8463312ce476fba4895cc4809db5da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82e54f7411e94700275b63f628f4543be3c976681a3509877c48c4eb988ccad5878d5423d9e776aac94eff90791bcb0d57e5e99540d6c88997858a022853f0614471;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da336b89866fb635c9125d3a940b23ce4f13aea5655bfcdeaf1abf98463dc584f921c09fec95802f69614a59986f76fd7f7e30e6010d97039b11bcdbd92d1eaa4b23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b491c23bdd9d81a028b3949a8715c50de03a09eb2d89d5b27b3b513bc1abd930af246eca9303a2c0d940af0d17ac51a5242824eda62909428ec6804dd598f6e01f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcec26b436d81969e22532cbe6aad734bdf1d8a139475892c7be79ed20ec3a9d3de1c0e35d66b63ff0f17ec5f9fb772321f544e694af93b935cafe424bb46707bcb24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88b03e6782ba782053c29ff963ca6a29e442146ae127cee97f019b20af2bdd9900abdac360e75df008e1e8197b87d97158fe992e38728034f7d97ec4988184091419;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73f73daceb8f2aa32c436e1248649f702f70838d76acd6a59d0648d1db830e63ec44706282450b85c4a4bd09426ea6595c9c3cef5bd795137ff472a737342ede895e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cdd55d8d3e279e3dacc31d94250ff099b8a4a5ec552e33aac1a38096273bec6f609c9dc7645c9163f8d241b1d0ecdf9cddcbe8ce1532a95919a146986e46bdc0b58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177788e578622c95a116438b9b3795ec5ae616859a9cfc6d7dfe12b8f421d2c0dd9cf44f75d60da4fb35da25b96999ec37f55f906085c8f09d9a5092823a97c522ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e2af0c0a567f4b8086a91964db804a2435e448411cd0db392f20de6b8d78bfe4db1f64eb78c29890f31c1aa0bf51becfafab5bb28f5df968b5009bb134ea8524af6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd980380a2e1b9f259d7f377bdee44eaddaf94c6be86a38adf4c5bb3606fd54da1d6292defcda9179458a251d3350c36da31176778acac436a882b05d19eae12368bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f463da9c692881c7dc4c717dd84a47d15cd69e1cbf6cf14f716c1545f78688dfe84d8221a5253208fedf690b969e67df9f03b0b77921287318f1ac2fafb842ca4684;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e94d813542bf221e70b406502e035a4f4dc04f342213c7d728c8b9e4141fe07df4f90c2570e02413caf532ebbfd101aa1bee27a6823390665cf39db37c85ebfd47ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha61ac641b0e0f139b979e865525b5565f6f84f516393d25408a8b2b94bc55bf0b58c3219c46ca4e475a392b9dee073e2e82e2fb1358176997b0af5f8f77f1951d74c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f9720fe53cbe7e1a1172087760cb2ed7754cdc6fe12ca0d4f6d600c898bff33357588604da5e54396a1008b59533c33c2b19ce711f080298091c18b397e1583fff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h239f4756df10f3df54d6957c94dc2041cf86ae7dd0163d3bfb979d7bb0512aa802db87830ad661c516e38f7b82ebfbccc41893a9cf93bdbf08f794deb421ee77f65e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b7ea4219d973d443d6c7145ab872db64f34f6e30b7c0091b6eeabd03e3ce64c1a942b82f92378626819bdf256f7f04129ad40717da9be1fef017a08bde6a709f940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183a46a6686e19bdbe1562a14597c409c885d1014af76a3bf98b717c629ac9811d38552b1bbc6ca06ec50011aa59ae8390ce6c76eccae851b6f8d31cb70594d4cf734;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121c17d2e22209d1cef51bee7c58b59fa127c3b31c53bcc55e9c8d23d14faf67c1414ee3d3e7f2a5f78df1d0af1f95ed98f5fff5bbf3cf267f612efa71c8e4b86474b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1182bc56fd6d67f11768da87cc244aff312c2101d9de5848bcf315b92a4310610e263fe8edfae7c0d7fb6b60c80b7f2d3a4303db68a6c0d36fecee7c6d2df26990154;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4abd0f393039d66a62a5cfd8d66ea859ed867b85828b2b750aa6c48c3251fba177b292d0e0bb240331bbff05696bbcdac4dc0b3c5228bd7b1748a7db98c6da951e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef74dc82a42f66cd8d58b0478946b2ea53b609cf5ae4af100187245f0c4757c55e456b1f313d1f338d8674f3fb2f24c2c9458f3e14ceb0e90db974b9229ad3c2c6f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1967bcdf65101b1cd197f0a49c7d1867126a6142f121c3c40b426bba6ca76723555d0e89d38c198683cf00dffc1124572095dfc334ffc65aa9cdee8db67ad607c0bcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b5ae277882ac59373b56f92097529bde015b93e5763dd17a194baccb4d1bfcf734dd4bb0be64e1fe439a664cd18c8c81c133fffb6811246fd120c9f0d18e73d8e50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c48e8859d75f3280f46d96a1f632c531555c7d39cd93ef2c97f531fa3e0e1edfee00ae0d5f878af87edaf60d028c1fd66caa36c831911d5be8c3ed50dcbf51db8e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc33a18081158342836e598347296c908cdbf33288606b76479db3d840a6613e964cfdad34b0cda96fc622605e73ce3fddc810a6c2425083837d014db28ca561b9dd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37e61855ad71616b14a3adefde58af0ab822955308add61b2519d45554faa7a213b82b715def2a313a464401b65a5bcc5b75bc85b5410ff41e4d338e7dee9fe1a0c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cfd4f37d882de607bbfaff615a1fa43978602e75361fcc2a89c23a24c0c79bb42416f7088db7452d016a6a8134ab953f6552c0e77297bb90000c0f373aa99962093;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138bfae8bb458c6f53f0ac35f3dd18653005006719cc4d1487cf508ceecd1911f7042840211e11110eef3973c13d270b186fb8e4881fa562e230494bdbff565d8b499;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd7a185ec591eb26d1885208470e9e178e33c9774801ac24a8351e6cf714b238af1f3cffa5a10c00d846047759c6c15cb43c274622e1290217f2133fdf006da4d3fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he39c53638af5a5a3ebbf25a5e09173786d919a4838e2c49edb5e31545cc983ca5c358db2c3d8747e1307a936aad7b18c651b0c649ad24328018b78c20d238bd0f959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff7dc07f9549d3255c1dc47d5e93772529a7a6883305bc33f6cdac2e4a082c6f57c689b97134915f6419fb28761a5eabe985d910acd1e9888af083c7927b5fda0519;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b1f4cdac5f2f512c7eeb82ede0ac59483edc1cf9a685922a009becdeeb5e7561c34a4014ddef27e29552e97755f855a9473458083f7bb4e51af58633428c577e874;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edb046f6bbdbfe4aa8b6fff40377142f5c6c3d11e2b6ec429f9382044f365a36d8cee9e11f8db399b39148dcafd57b5a6e2e624aff63c9f298dfae2e2a51119ae279;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f66c7b7d5b72436e3e661fac756e507216c0d2323ed88fcf9ea94a26080c9d66a3425d62c2a648681b24a198eae656b7f431744a59ac61fd4e89b84f110aae854faf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11118d3e1c665ed11a5077ad1316811fbce5791c31a95f750187ecdd34a78906fb279ac098571fa1373e3f784964081e94722071d18cb467fe6e6ae84fb3ec9fe27b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hecd26eefa7f81c62c0d8554ea92e79a96c72e70ec897184f15b62addf4b3c8a2e78dd305b27622e6020bf5a6f201a60028dbe75b3a9bb34df125a0c3edbbd1b2c4a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98fbdca5af6b5c190d6652f0034fe94c47b7cae008b1cff618c676b87f53c8d37f7a30e0fc935f0ba659dfcd9a9254fb14d0a8777c58bcd5cbc7aceec854a10a7937;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f184f4ff3ec7bbac73d401fab73ed016ba8f53028c91b9715755f68368f455415a858c35a3b870079e06dc7c00e52a5941e46197ab3652f6b543554d0465b6c0c90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2e2b4b260e9fed091174312b14119e1beddeaf1d957222478ac4121b027a4e0553bd817cb118578e7fe863eadd2e711a6b444fedf95ec39d9aee2201678d8313198;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fde80dcff3ef337e09fb6a93f35bcdf8909f6c43479f94c4e031acb396e5bb8d76da970b88ba226676c36c391f75e7b98393e944dafabde9c21e0387343c85c82c3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h791ba89ce8ddc6a4c62303fa79ff7249a2d877c7eaf74f898c1f468bcfb464f1ad6e1862ccef1b3291e9947f0cf3af82581c73ad47a628bdf9ce4c435904fe1f6d95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h629baae178173ce289d42fb4617638a7906502c1c456767c12bc05f91a847e0efeb300435401f350523343c9509a35940030681d324e7d28adcc38a3c3948ec4bcbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74922b28df0c1900eee5d7d2b44354f6723469645626455a9e2f1e3e2ed012b27c3b49b44b154214b76596f14eb2d76abc0b1a03e15babc3e00077e27ab69303aa66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18776a259cb259b4d01c61dbe766113b728b95e5ba5073725fab943c16dab854e410f7f885340a2f49accfb50000b5c1e6355d3c0050067128299ef8c51e5fdd6e5c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31674233679414dbcdbc01d3f175052782fb4fca9244578e28489c69d84877c3b5753728daf7d9aabd2ab571feb86d1205eb99101a2bef2cea0e97fdbf283835cc91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c4f78e6a3a5ea02f2a204ef112459053e9bc381fb6adecf5a94477129cd0d9fc8566eafb918be91aa988b86af7902e1968edfb767fbc1f6690e379b7521638790c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he90de24bd228a884fd125bcb8e1600c4afa48f310e93078055fcaf6d560c4f2c7bf0b544c4a27fa9f99ca885236a1cae0a4a7266a5216d3b331fe53485dd5ac54b3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c255465d22590a8258bf074f33c7cbd081be62a88314559de47b9351315186321602c06c5608f8126569aefbad3fd6f0f0a4a3b89dc58b67abd017616ef02e1b34a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14dfe40a501582e23786d7f094fc01febd0550ddab02088945c84bf8454aeaa0a0b71dc27073ed0bbc4375e56a5a8fff8c3fcde8e9e49c38bdc9564cf9f542fa7be0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc59b62cac5659f1bba9f119d2165f9b5c0c8fc6e0c35e6bf23c6f329c688fc2757873e60b75b6d03c85754c35de2a298c22bb3246adc2af89648dd7ba2dc95f603e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3818935101e9535639ef123ecebb6673f307ce48549b63f599f6b8326a4f98dbfa86a7683b90cc774f41dabf353f02628cca8907c41d51148cd903cc08121aa73fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a0609435e7b461c7e7fa9e6871bb1d7e6fda9d62e79b254dcbdfc855cb30caf191c0c066a88420d4987a79461b7243cb5200e406e3d1e5a3d0f6f7681f9d1851cf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hacb7b468d6340eed51cf9c1badaa08de2853dac666d33532200323f46ef0596f924ba8dd3de9be70410dc13c1fd63b5af10a1faca1f032384e380f4741ed9d19728c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dd7f3e5cc97d19d82a0b71760c56cf036543abebb4221983505c6316aa4b0c8c8f6d667f5966e4b048f79f43a0c645c14143397716b42a8beaef65a298bf791c13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he838e242372dc4790ea9ef9d727adc9e5f1e6c2f088e03aa66c773d3c091ca210a77db5f4bdbe6fb9dbbf15c1f6afbee683c5db9f6899f2131d71f295818b862eec9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27062948973231b17d413508d254d3e13471f6aaa136bb024ada235f96d1258b9eae5e948c4b5294d868238d026ba6e526c64b5628fd2d81ab766375e23d233def8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142fc08a3b4f0c5b2fbccaf94d328fb40f70f37716a81ba906410107cae80ae2e99afc42691b321114b6d1115552262427e075b396b374e53e1d14b301d087b54416;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h473ec49a9f2f10acc6c6dacb16bd025e8693a9ef8a85f976503f7d3c85d7d90735bb1d3fb2e25f15965702193dd0056205ef9622046bd8b24a1b780499f8dd626780;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166672746a4a78c01f6cbcd9132177bc2c240c316968fa6ab55b33f26c0c56182e20d2d12c5f4b92aafe44dc6cfb7e4736d9de786251453e5ea237f478d686b153cd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1971b2f88ea2e9f61144816a9ce1873823a3fcb301bacafe72d5aea2beec4aad14a24449a6b1dd22461793d46eecabf7538f12b0ace27880c2216d49bbf9a0346bb84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1169b40c0db552f814529c401d6125515c67b639d3178917b052a4fe52f7eeea03abffbe5177dd22891d4a565cc056afbae71a75db556c7b9c5624573587f974ef520;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14070c91f7355ecd1a47dbea63912e024097f483490ef102a3fadfd4e0533d5e6d907445d8c79a0715ccd578bd26bf6e0ab6ba7329ba012adf4ea192be055e001ac06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b351a84b60eaa57d9a1c5aa926a819e0d60cfb858ff9f6d04600814f607508d1c6e12ce260121cebcf60892d5576f578ef3b471af4b395da3c320a7f31ff6960b6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81f6d458262b6b1c40b79e5c892286d4c3d35811921975b3c0275987c6e0855824ad7ca6ba1c663d290cd2f7a21141ee2aa38e884dab8dad0c1aed4f350b70ece5df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he258a7602303303f045f285ddd486f811bdb0270846b094273ece3c09e57c1deb1545bf54b2feb616a4b27d7862ab7fd2c9bf00d537f2204bf55c821f66f83c53beb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f1f65c9503491d4007843b89ce15eac4e92269925f7e0a45c500072890c5397e0f349398ad025d32028888788620cd073e22a2f7b0ef7f57adbb0b4aac642e0f378;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf2c168c0abf7821ff791b606e956f5db244b705941c5f60d8479b46e23735f833a7b8e0e96971abf39bbc5e0100b593af1c2dc03590714105fe553ee1c62abf425e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4eb430868e45abd3a5f226f60e8d1634671da6a727878f4362d8d4f88a691bcefae746c6dc9773d10dcca5884967bc08f0029e6a3f5e70fe6e1181037f84349472a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h939579635c5eb035016f89c7c00e3dbe50c2833746231dd3916457cdf2a5ffc583ed61f48bc7c81d246e2f17ffba5295a3e8dc621b6d958bf4257b236767821a33f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h869d5a9664d4de7228b4f3e4c16f2dec82810e08b5352e55c4287b4cd0dc6c02b1f3a2bb1deb1d944d1a324263f6c4cea7f896fbf978490b345569d9bdef388cb100;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c65ee12da471de811f776485f06b4ff1b1d09897f1e1357f6e88b053374fae5b052e40ec3ce51ea38b3e6cc890b193eef5c0e97500cde15dfb02d701340f9eedd41e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102514e729ee77b0926125245df11649e0933494bdbf2a75bc846d0751bde11ad752bac37dbd1eb06138b0d4cf20b57b45aa505fbd95cd17fa2a41b1f37880f304fdb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4587331e3531e5e95d467db0a091bb14ca2954f59097017f1bca0da15ebb985db2694ceeaafe80eb4c1f81eb3b129f8b09c348272442c434ae4320b7af7b669706fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8427ccf9167ddf15984afc4d962439f3aa2028d5393fdfc21ad5d9b270f7251b486b0d96b6149ae45eae2f24d24cb79e8e412fa2135e6ca2ac4c2972d8a9e45f8e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b599178631f326b3b9c80fbd9e6a48086001a3186024b6161ed13c0dc5ec2e300c7eff577acb4ecb7036224df8339991ac9e707294b0a06d6da3210a56dbc46ad05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b7302de72be5d8e272e1a24502ae5405d3b9870110c799441d129198e3647656a34660c248ecc23f799fa4c15376f10b7a0841e3f903da51ce336c86eb3e6a0da9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e0c9d9ac567e8229bb820640b364c90820c5549af43d1615eb42f17bcad7e5ba0872b5aa8a10d761b5fa5ff01c283a137dfabbee1f03227837f739947aada90031a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e7f588d5c2f8541ce1c7362551ef839ba758a68c4516b7574f2345a26185b87b6298f881e27fc39bf357b6276034287eb6dcbfada14ae0d0ddcc5b4a5395011c507;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5552fc63bd7443236befb58a7165fcf39c2fa96b265e461b6c52726e5f907af70f01ee3ad9e06b27ac23abe1150bd1ac716410ded7f94d870e2d6a4454a7c802dbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1e9815bfbf484e31509d4a33cc8391c2cb0ba6ae029ee426721fe37d39a516cbd16e1d684d40e14804d59f4692350a9f2e3eb2915284a0cf2d2fa462fcd63743256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0acd339475b3d2a602a778f7c9b723bf95ee9217919c14f049d47e9d44697470da85796171afc03488841dd453ef94dbd6eb750f96e1b6aae126d19d0021ece3f21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64966f8ce5c9c740d9b7eba47707669ee337788fede82392f6028e35a3b1e226cb63f38090edfeda5c2d727327ad30bbe5438b51e7b2dd4362f8042066978d9294e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb15e6f2dfb2cadcda7f62ffa49c4298141d82037a33ff5afe267c7f2b90a941f6bab96aa99b63b7b8f9f38e16c7f6f7230897cd4a7d723bb056143a1c70f21bf6569;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125a8441835807e3063b5c93e0bfbb9892ac2b887bdda14b425f8b5bddfc5f9b53a64c76df64eed5f4ef17e0eea841a93aec4b6398e4392b37c505b134f0a3d4587f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e2d66a5e2935e6879cffbaa1c6d2ae77e1773515a624a3060edfc37fc63d9d2ca5ed4be8f07dc8002ed35270fae1086eee19a8b3eb7b7af4a1ea682fdf1a6ec04c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27429656869931ff1e46adfdd25f4adc07c95315a7d02a60b418b57ba9dbc97008d9d86674908bb73daba4ac30a28b58f81984a211082b8539c27b78fb863d68e40c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa643ad8bc148d488dc84757e9c93c0595abde7d08f87e9cda9334b4061d44adb017bf6c96d321f71909bda6e604cd851ddbfa275aed9065bf4937b2221ba702186f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca5503188fbab2c757f769844333751ccbdd2b40a176ee4c05922ea689e7e7202ee23b66d135939c7408e09a343ce638b9ba63e67f5bbe05d94b2b0f27f0a0f3a48b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa0c6618d11b01ca861a7f06fd0ba009305af6923b1d7f37de2eea4b5aabde56c60a01640d28ae280dfc4f438046462a3e2f745c712086a4f431dd93f92d9251fdd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d49b3926c1d023e8129b3c61d7d8d15cf75823eb32be25d79703377a71f57b6e73e6d8c6bb93b878dc0c03a36e1bbd5d3121e8a4ca382643f422c96a9230fecdd4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d25acc1b2817ecd0de6e14ed455463e73ab43b6862e0b4f881c9cb68d84519a16a177c7fc8436e70d7a077b150488b3c3faeb57f6d4bf7c324990c14e88779048f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f316da6234be49d9854daa835d99ebf1f34950c4e38f4256aaec8fede9e6cb2b725cf19a244b88666c17d84c71a302a92c3326b30eab2d062d007e897c500e67335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c18e1f0230ef400661fc4f2793cf39be7e31b930cbd0eb0b2d032e3f31a753f432bee4b3aa56dc23bb2b3a2c59e337053a3918bb9a380c5104d793c1303a9aa7275e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h967620a1ba42f4acc82ec7e92fd2888f6749fffea65aea8f77227069e0d50b2aea3a7179419a4a0852df974c163f5b2f0b198775f5caea006ad6e18e326a2255124d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf3a6b12f43c305fbd4cb4de44c8f0ecdb4627b227fa3e1094efcc61b699ad4d562a0740f9d6ba74bd22692558247c29434df1a8dd02ccacda124d8629d693dc5d9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf65bf0337ad2e6d130c0f2acf48204cebcfc6a3b267d681be672f007e74e52a1f45408e192978e78553c88bb4469f72b21bc6940dc4b41c869463c6a41933ce8ed62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a95be5900b8386b04450614717e5563d82c9779e1ab265934bb35f5a1d6f4548d067a2aeb0b7e97eb23c21218fd2dbeee6b93c3ef3d0f5530197ff6c9a4c86313ba5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30c02f6bbfed19ba79db7a70ac49a77e0a645ed35d58e88faf4724eff719808f967c6170c0498e3e30e2638a89e3707f3738f7cdd4f1a31d0b7b8851bf7286df4a98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd19167e602c9e6961b4b62a229ef4d273454d79583680e571b3f49f580e093f3c89e22cd2410b78f1bb6eb8113fd7d6e66e4b037a35a4a21cb907cd17803a8dd58e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hccea548e9aa89753b22f791a9f7211a23a786ab76f8f957a5fa4f91b01b8acca022678073f4b8deb711004693f3702e2ed8da5f2bb205c6149138a5cabcb835c60b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h603bd5b18f6cc2edd86a95410e379916f2d1dcba04d9ffeeaf08f1b201c8faeda9ef4f30e11112b3d7a87609e8a52af1465c54b7c862c08b3e7286d3dfad9e3d72f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa88a0f66fa6abc25a6e93a3e994d208bb9ea88729ff1a272089abaa0a7b60de735f604227430e839ee1d5412ce6f66dd649de568252f68323529cd8b388eafcc7fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126f47b1b9dccf1bddfcfefccf1db007e1e495a5dda441a76933ebad8027b2b7e8c3fb09505d3e56bd003907ebd18452d89a5a4135ab38adc310110216703a21924b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a2b70028ab27d51a6ea74d6adaab3729314a692bacab00eed7798373f29d0c7a724edd9d40b71dd228f9fc052ba5f88aa4b4e29dbc3e4e4d09e6ee4309c8e11636e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145fa4c3cf015de66f1034c9051329b73a2f322d0af47b96d5c78ebf1247bbeeb9a6cce3b05966ebfcb7dd0714325978beb052662472268242ede2d05e8f0168e73a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dd7b3e6de87793fdf0c6275538137eb38a067464572cc784013777e5c6b1d0c16964fc8b7501db6bf347f5ce7684d1ef585fde9ef7b4478ce5ac66e020e3dd4d8f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf32eb3aad0d0f50c669d1e0ecc896f2761114891a628e420692287e2c04ffb3ef9a4f880e1263c115f56323a9fc8d71820605d58480074ba69a38489eaa8508194c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73e96824b057d6e14f0d187f6002ff70fd3550cb3017d42eb33c0171a5bdcdf185e326832e48b38cfd3dfad655cf84d19d53c30368acb33b4f3e5233e95515b66a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6d2bd26fddbd2478f1ffd9c775be02d43b980e63612661bdd17a0911ef5e7e8b8d64918df7d63ed154f63a7810069b5401a791339a02aa2f74774aabac395b59959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169aead9bc3fdabff7edf2666872af8df67653c99651733e72515a8c5c6a5e7e917307b5100f6db5c9aaaf70482cf7e01fb21edf667ff0a200d832511ae830b352d16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154ea8e706bdf72befe939f8ba86cda86199c7bed72cf8d133018715b6676c55c6ed24d5f58def2f7416575a0f959b41f8cb748b84bf4432ad04da9546d2649d51ee4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed227e0984bb84bf1ee574535e8e4b81dd16e4ad059631d6374eb57f2661319dc467b0641c1200525bd66cef9d08ca97881b279a67f76dfdf3c7b15be863971e5a7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e21fff343ec60cf4018096498a62564a4e58118999d2e022c570096533f52cce1c9bb227429a9d6e0847f75c98dde2a874fdfa6e1d7ef6d309cf9a6f44160f927d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f33282d5105ae74158f9ce30d0059e3ce3f64b57bcccb79f00b0ff1ed20032f302c1b767eef10b1bcab88d63404df2108f6d653be4cc61735ce915cb04b22a65196;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafd6dd92c3d74817dbe3abebe3c345c2c6005b1031261859128d9f4c812cd4131a7aa2af96697026ba0ef4cddfe5f1c301d710b53786e8bcb3ec14e4308007aa1070;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0d4d88d7a1068047e8b449713c7c512f8084f1ea3c12a22a0a00ba0d3068f4d7b241c929703224b31cdc4f1e6958254ac87e98e574dae125c4d5c0b48803a427985;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1053c535abe45fedc2b4b16f6625946274371cbe158d84ab3568567595dc8db119d3c5a35fa02fedd7ba4fd1167ca09de73521f910c96f08ddcf43584d4a6f771c88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44c08752c0512ad9ad36bf9d55beb8d92ff8f1ad01a58c68270590a8cfb48b2eff8362a5312d7e61c4ce36605e162028fbe3410693f25786143fd426a1286a07a530;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171c958aaf030f53b8b90c01f1ba786f9318956229ba9fd58706202430c8db26f3de6cb27df77707caa86402e6c4f8639de14ee281d8c0cb5180ec11335717dab9aa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebff631af8325353865732e3c314b78d87dd2acf298b77b005df421929ceec7f5b425d6d0b816712ba56e5286d59dc4976b8b2c8644210b23219cb30c0c78657ee7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h531ec42187e08fa37d28c615169b7dcf4ebe9527a739106520768ae970f0fd24a46471852362172a7eeb75e414ed99f3ed0720ef5b7ce5bbce379fe09c4c75729fd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2e20a0be7ea1a9f49d009af493dd9c3a54053d50dc068489f9e4d47ba2c504aebe8192dd6e599a74a02e539cdfabaa543d0e2d73f056229b42cbfdc46f96c49d6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd24b771900ca07c39b96debacdfa3fb11f7ae1361eb924c36e026dd3516f8162d7a0dfc156687a7c71bb2efaf16583002fedd3353c79b68404c57f5514c5762d60a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1970c68b47e81b80523e4d17ddbb79407df69ca7eb5ff14e94de2548d9d0ff848637cb53c93ed32c04805ee1cc793468ccc6f8f7f345bcf4967d46d65678517723d10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c43f0bf8fc2c4e0f14710958f17dca5f2fb650a7feb6dc1afc1e11ce7041ed92066c38232320e73388b202aca19e6c6cde9822a053b6db3efc49328fcf4b5d647282;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1771b7301df9876f1a6697c27649641db31c769435827ae07d94f188ae7ce81e1658549644386ab7679fbee81df23c4ed742b66982d79ee7944aec520f6e866cd9801;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafde49560538b96ca2d23e25f613eae2d54bf53ec3a2572fc3e00a0c208138d3397fd07bce0def977536f285645e5b455cf6b566da9726b3ffb97abed420202ccb96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3f80a22afcb8f5a250ab3db3d723d981e2f31f366a9cf835fec6d2189a97097d02125683fb8f1e6cda8b7527412534abeb21b4a475c7b06b81f561c90c1e81281b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h203a95e51ea2b716ee8592c17a30aacc0eebd720be5437fb57d1b50ed63019d3a37938031b01c4d853b249785904f7874e0d14ca7032a1d3826ca8cc4a333fb0b7f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c1d5e40a5d84b4f9e6452fde4a0839a8d7acc3af718990b8a6a3ec0be63f5c8cfa6b6eb7d6dd210f685e3261ce3ab2d408d7894f5f5d4887cbeecda8f7fe365a50c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84a2dd3aac25e599ebacdf6298291d202ab76e562a1162bf1235eadb680980fdcefe2eb5381d6ee50302d365f9bd7d0a0d00ccd127dcf0f9f9c2dbfe03090469d8a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c69e75a7025f7c225479a58175a6abf2eb696f7164ab234aa178cc9f96f748cd309d81fd2790fa090fda406546d08ccefc82656f098edf264551c93a1ff6392bec1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1357a0f2f2498a8a369162e5c5ce9e3077d43da61e7ddd53c9346aabce8098444b434e3acb004a3c03cc908e947ab19eeb12a775ea8c146b741703c5cead09d515963;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194b586c674505906a335964f9cc84aa592384206d31c353811eca1ce8ae917391b6892696fc4c64cf2ebe0867106deda4b9ecde61f443df840793cc3d09b6277b571;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e88c202ea47cc949b3153aaa1cd51e4c1e4786a13915f9c5cadd9cd532e624c29ecbba4f6561448fc5a20ff369d8a37b2f80aff7eb2cd1def8945aa1f1a525c1513;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13597fb8b3d9308303257489b4d9c5343d8747f2d0aa86048f20c3d330057abfcd0a364122421107068ae41a35071c68c2db7570dc6ccd47b8073a7adf871856f12ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2b3c389f91039a8f22808b5d4cc146e27336dffb133bc508d3b9b97617cada93f68bd809bee1056b8ca6ad4874c99b30e3a7bcd14eda8cea80e0d854720789534d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0ee28ace87a10753223594b29b37155e904d6a4ecde3db423b93b24cf6299c6338481600f89d1a6a4a28d8bcf788089d1d34cb0b7e17ec845bd157cb3ff26fbb27f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he232a5ece9e09492ead2d9432243f644c0f73963c82d5b6b5a522a74d8d5ef8ace0120042d27a794482af35d822ec76b26d9996d7061bc5bec82e90926ec85e4de37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d71e9f000ab6be3a3a09c1e9a3fba23131234a8cfb4a52f567228f082da4ad87ce61c577132d315db465a99f233d600663d2d2b4b0a1bddc91d5878528357f21596;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fe80b61abe4c0961d789b1727300fbe7e3cd0f3a578486539a817f5d6e6898de30087bf5754c82190af8f6c6984787e78071af16e79d3e4262c9277d2363a37dc34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1257eceda48494ff005962a8c23bbfe7b5b242c6531f7fde36c3f319d28b0b51bb14148d4e99d6dac7554f29a39183888b2ae1287e0b50eb30d5014418006b915644;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17731634447cd34a858d3759f929c15fccfe357b289b7161bba1c346a552ee50bc68c9d192c0a2e78c8e0f4c6dcf34031033d3e106ceba549c5c2c0e881fc223cca9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168fc7e5e141c1fe19fdd3c724f58ddec0fbb1a651ae44d574712796ebe3ee917eb27e6545e797ace1c4de3840aa78b9333993a68ef5307ba73877cc9ce8dae6d32eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df99b37e3c22cdf223e239784db1c97a00cb323eb4b94dd6cde43215c5450e716242a1d0448d745556204013f95f4620e11fc62ccd1b209fbafc81202119e94f494a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a291e06688c83631a4c852dce4fadb06c6a3488d3cbe512167ceff29fbcb307084da2ea615551db31de36b6d31b05346528519c22e741ee42f3497879e9408e7ed09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112ff37bbc600cbac19988de7f9fbd97620660c3b8f6d23078fc5e09d024a5ca467167ab0b9590fd98baeb1bff958a7ad14dc860c3e11ee6966b6dc6a1eeff98b1111;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1430748eb9370958f743a5b047e66b7451d45631d865c924e63d0af9fde0b45a25628b50b449927240072919a8d8ce4de0dda798a94f606735b2fba61813e211c2ff4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h646f4625103d4ecec823ddc2fa66cb553117bd4cfe53d4bceb013b4bbfa19a506110356d47f9abe1d314b9203eabc0e94b975d82c35646c699ba391dd3a728dd978e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12441310b95495a4378914db93b65b800ae2f4f67879928d8d09e1b71c4f08f92db94c64449307b9c0c0f76a478eea2c0586d782ad40ef603a7f6205af6699a4d699a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e6bd6642c6cdb210e94e710563455fae7fa4310d4d0a065f30e20da7716fb1cd33442e16846d38ee24c6bc838fb6c338d9c8938eb4842273c80f942f2597d01257b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1300dd4d2123bdd96fe1f181a228943ae0bdd1975d3b76689d89d14c8e18dd78ddc962baba677dd88c89f206c903bbaac6564984b72df5dff508a7ac1e79d665aee65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c29a4b7a839e2c3b06851ea892ef38253994b7375cecd7c4375e7ae73cb87b618ebe003bed9ee68b7d1fdd22e0d795987d952b1571deee4df19e02b29ca7d33e9ca4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h432c9a575691b1f8119d37460e58ababdebcf3a9ae8436af9742e425855fd4c2e6038e4f3aae8f8ef378b0c6e83f4776289fe524937f48fc0c0c9d742dd60f4809a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41c0cc1c1a6afdefb5dface4d752196bb36513254fa9e5e41555c3c76ad45aebcf1a6b55231a43cbd113bf03beb7f736975fdef21c58fbdb7800949ead31b9589a3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb279c5eae78f6ec73c3fab6596610145a0e3716f65812536ff424058d57b2499cba5a4b78ab83034184bd90484af708bd6247bdedc9b9ca42d13c74beaee78dceb50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f06cef0085771940158cda11f4141821eee56ed6ae4758f98e8b2f0fac1407aadd6dc37e5b37ba117cf7cda66a6d7920b5be5e19a40e16ccda2cc610a6b6d78a4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a6e7ed485b91756dc8e0dfe4d63a71edb831e4e97b508bf6fcd18fa02a26024fb10b02951c5b55aa41ad7423439ed1b05c67f26db13e4589c4ce68e9fc132ef4e5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3fbe716f89ec38e1fbf78a0ec4b3fa31d34168e13d3293cbdc037dac3d094197b22979afd91c2f4782fd9d5531285d44eee1f8fcaa56d21c380c529f8d834abbab9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faea928af08ada2a43726e38f3e07f7e0e78d9e752ced4d81c5d1ee85ec138e5964bc37063a30301044d5c14cd84e2183225013d64b693db0182fd26422200ad4df5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h842b1bac49e6a1ba90141f68f971c614a8a4efd51482f6030c9caa0c19d488506cccf4337ee17733770d2790bcaeb5688bb079abaee78ed5834836d7893c3cec6e79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8052352e63bcaf9c913b9fc5fb044e2d6eb0b372d843348eea8c53d1aecd6188d1eb209e07b09720c87bc4a28dd6169c77ece49f37ffc58a573227d5c9d7b82e5c8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h213d82bdd0a59810a2867827d24a03de1f4b22228bfd57f33403fc31251d1959dfe435e114d3d7677bb51b5182655afe4d6f3b3a8275c2e0c0386bc051648fd43b75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f034106148d3b5df967ea638f8c087685ce40bfe07f187393923b73fd81a865725dc483ff896f87178eee392413afd6e16893e0f72a1f0f730e31355ae098122e0d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60fc8c40d9add838e421be235d5ac8f1db1601e3bb779b7fc91e66f62eed73d736b40faa813639a3c868e76a70585c81ec16399f539767eea5d6df4b72948cb33618;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1618786cccc2fd5b21da47bc28ca7ff344141bafd6b2cc8b01b41dedf4753167c6357333154f41e033f913c3e9ef66a7b5eab2a3c4228c0d86d29c46e14acc086b0ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73dc721615d3c5208fda58b2e385f5a7c4a5174e0144b620bd905b63a33926a0df681a2b3bf77784a1c91a2a2253e353f840bd9ff17b0be42a981ed363479cc78d92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a354b73d37a508dee01868c18ec4e480023dffc4573beb1ac4b407b0c9c3aac6b5c93050bd005a1f0c8792b78b5c156e17549e4de879fa2f3f500b94cf72c4cb7cd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a4984ef78d7e48329bd4669a1adf14c7b3ac8f3e7e343cf1f693b636476e18c08bb01c1c9ce0a06a7f74ae76789c53a6f7c88fe604e95489eec52b686a80b50d3ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181d0990dd371ae19061d1c9c9def5204ed0c1e704e3ce0eedb2547171b486a3f751922c317ca99de2e8518e6b0635d990d9e1ffa3b41aa78ad73e92a88af00af12e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e104af945360af3eeab8451164dfeb55eb96c7664b8eb3d499e8f2e6276e29930e9355be2cc3e15152db2e8acf877602e74014d2c9f936ae7a2080defd8a44f0c6be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab204bb56239e453d80d66c736a34508e561e5ddb2529ded9ef8f96043371076de3bbee06c5e9531733669a7d502b4214f1adcb704136fd66823d6e2dfbeadae755b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7d0c4b3e11e744ea6d171dc6a46fbc1f45284ae9dbd1cef267a335af62a104a2aa98909c634e1608a85d8df1cd591844d1ba06479f8e5266e0ea88609b89f650987;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ca1eb2756407c878ba12251f37524f4d7458a666d28fadc5b13613037bb75938ec970f8a83d00f9d2cf61f0485d657e7c62502bdb10d6f36ac5127e4c6b7193511f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc87c36e743f4f24a30d7e4971a653a98bb135cae1b3bd85c3c8d471a7259f416ba49e24b6e7e7d0f4084be9257d573d79613d682674aa8fd190a3f9e26f181d03ee0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1319386ff381c6a2f4839395b1b8c09d4274a6a7ef0a64c1d7fb7a4b7275a499264fe91d6947e8d6e9a43e01eb01da07e39b3ef777a7aeb5990332dcac117f4aa8854;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9df57eeefa752db3733d2e9026840ae28ef6e082af3a9a3844fba802d79b14a715237f8539bc3c5474f1cc596f57ac3068e7fa9d40a9e5e1fa14236e1e4981702003;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149048ffbd6eae6fd9d32c48fd10dffbd7e582507285e5d5ab299857975f5bb5c18e1560bc2e183751012285b582339524a7b10f467952d6c806b14864a65cab0fbbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h239e074410f686920f99463c2d080d571399a52d896ac7a78454f9037b4c7431242f7a211969fb73a342c0abb7210f82beac8f3ce444024dd6c7261150ca9b821ea3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdaee746e06ee1378867e40e52daa8413e5c6a179bbf930272393736187016be4a3d744adfa4965111eaced3ff8cf4c3a1d7f29305e858508797d35c67f96cba8c2e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25b586b63fb7f02d4e06be9033e36f27c0d2ed69a0a8cc8a910e2b6162b5115004118dd79b7c3c667a83bbc8206f5236c8fc51a01578af0ee50a3e65969b18b1bd25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86a6e47ae68163120e03c9062f884db398fafdbdcf5c99c3da5bf91aa304cc8c981258847f1c3604d37e7de8828fae4f115b45d6f5bb5119e8c01ff9885ac089c4bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd9cae54c4abc5d229ec193308e08157ea11c5ddb00fdb8ce45e888d2932d6fcbf52206c53d9f100ffe885f18d4021f3ada466d09aea52cbcfc4756b54c03447c1d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94f2cabbf8f89fc3e609c295a9428c3634c18eaf112c17094227b08cfe2691265f8865a8ea22b95c33492412db0ba185f9a9935640dd4dd115dfd6e11523fe6423f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14630b4698fd694f18d7f94c35b359eca22a2650074c4cb6bd5409222be5bde4afe3222120123a62c84be826e5b0cae5a7c6f64d6cc6ce7228a72ad990c5a29061abb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69afb8f125b731e9b1f5a2f2cdda364fd8a8b085a7c17ec1b31a59f4ede0f73c329e1d00d44f924c2de9c014f52871953856dce651161f317fdbb378eb65ca0fcd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f84334231577f7226fe8431fd0f324c35101c0281a7e51e9c1885b2affdda519dfbc5fe8684043c55c0292e0ff9ef4ce265ad749ec5163f0b4438bc762dd53c85c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e434c9c40538b16aa76ba9bf7f51d18a47e1c8038edf9e7c0299322118f8736fdff22373c73ccc117388e5494ca6d4637e9f49973210b09483292f56b06b1dfe27f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178614bb64825b31bdbcaaa91de3ce564a00a120c314a1285a962f34b6b26c34ddb3c469b181dc0574f6efe599e363a9b5d34e32fa40cccd24c61bdaa892847d5d1fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f5da4781e751b58faeb70d19eced62d27ac431726b71db6ab08fceb720c6e02babd139dc6762c6265f765dad772fdcd5def395a4b3751f1f558686b4271e4c71b4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1398f38d87e3d266ce4d61c6185a267e9298302ec485b943befb493d8db6253ff13f1c9f179ca7e59a842091a325cef70879da060f4d6fba50fc68bbe0af1127eec7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e3ae8b26222f7211c5df8ed768cd1e511e482a9af636ca0c717438914d1b3cc856591dc8d160ae9c26bac17e1107a6875e1eb7eebd61ca9a8131e7f981aead711d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc35d9240374aae55e1bb62cb27deed7dfb00c6c57b4672b9f210747f0ab831ff6b0724238bbeddfdb6bcd0c414d4986504de74404a59208411acc33d9a72a2afe69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c8cec30750fd34d309a4cbbd2c4b4bb55fb63498f836d60d3636f7006f3f2b70c251b0d030881ecb8bb2a3d547ca1cce50d2ca1b80f3920fb4f53ce1c8c654764ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfa2b1335d90832f65b3df099d429200de059d77f2e99c4961f47f4a849a9f0793bd30da25dbe5e4b92e2db55882dceec6f1ddf33bced752737bf06a272bd8b24201;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8db91685214b1aab7738156e31bddefac6e63f95b76ab0fa1290fa927d81a2fddf1298198c1ecd5a02f405e5ba29e200a8702d3ca16a39d03c858abd1dc77524497;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eae6bc6aab15ddea11b82a6960c2f04588f73385a8a23bc195bba6c2642a75f53e9478ca78b269b25102e48550a3ceb5f07516950d2d9b1a3dcaffc887d61fe3b778;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d362eb45b386713d89df178dfe0bbdafb4ece655b495e32b8f749f46c4618c800bb75828c3426c5f66b9781ce5157ac56100e4fb0d58856e96b42f0dda773c44a864;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dc8960f1914c8f133be59ba4d82fd38f803ad8347f3dd389b7a3e9c404f1cda31b10dea0349ee307047ea2045fd23b03e4d4515ae8ffa5c98b97b92a33f66aeeaf2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1defc181dbdc4042df0e59b979315f528b08eecc592617c44a1c5c958cf4790225be2dcf0ffde02a2c7ded8f4e73a36986ff34766825c1e42092026f6d78e42a3ca39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he942faf51184a3fa2fadeb1c7e46182924b086461953cb84e7b1033bc9069045f1e453c2fd83abf38d0afd76681a81eb0a67f71dd8462ac6976d2278f86386566a59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91106ab0b0e7c4d8c241a7afa7277a376f9ce5bce01715586e94c07ed581b2f17fd9a9b4381942099314988d1042ddcae52ae3929109ae09d9fbf5bdc8399aa21abc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6445193ef411bfe0059dfad188a20c4f7a4bf30392ab5e4b992b8896ccbfbba322c78d8874952c226a391dc1fe6da21401df21a93bf92fd654372f0a2653d72ae43b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f9f9f683290160cbb348c46604bb2351f25e95766d1a2cff453beaa8a72272f76fd5874c51b2669972bba256dae0144df2cf1876a0187bf071bbddf8115b6ebf750;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h460eb30377930ee52bed0f6d030274d925e91d1178851911cec204e6ee796b775807ff3db8437167eab51dcb47c4917c6722bee39a97a966f7d622f1c3275ae3f86b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f42c1dba38577e740f175b186359ada1b16283c6bcaff2e2abc18123f3c3a9f745d9f1eab3068603905e3d28e923ddd56fe2f5b06e8bab3a18bae57bcf27dc9e3f28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87679e55e60641065df30ecb90251b464196ecae416ca8279b79428a9e98feea6af03e4283c6409aa93af2b6c406f11009ea08009e62270577eaf65ea52578ec5d10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c428cab84d4b22a83088f2d2f7f195ea3038ee33fb7d5da3b2b4390b35880b5b4f9c750f1b0441bf2fccb524d34187448d7ffc2a48e32518b5f7a02c928fcb79b25f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172e1c205e149038edffc2ab37c7cb7cec9a41efc903d15616294284e9b28851c214b40db78a2a7f67fadf14bb498605848fd95fa6abab06d2e3b4851ed66a932c451;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78a6acbdbf923213f27054968bf02adcf743cf173245b88d54431610e7194ed4b063864f75fe83da4e954776d1ee79626209a2f2f915bbe9c64cb315132b3f34213b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151a99822db18584275a7a11971b7ff297caca4a09a97bc3da44e7136d10cf6b6a12412e95abbe4c569ab0c4e8b39598f109590fd3df1fc12a312c96bfa94692b2bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7061b9e2ee80bf2a46d41e0a77280cc908af7774fc4a333b2db9d3d8e6131c5a7621a671354d6885301d253209397cd0cdc160ec91dcabe6f6c12849b9d6e3149bbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfef6f78981953fa2de367b2b5bedc3e564012a3df92698f70dd10da0f218a728896f4632d58ee654e2d81d6723af988c73fec3b3e509c04d2287f058fd9d9ba5e727;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he509909dcb030b1faeef6e3a3fa0606bebd419e222390b7794aaeb52a17750bbd861c354e55b9b9119acb98c1d8a1610bb294cc9c25aecf2cadd22ff94d6e23748b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed468347b30d98550e07e9a3f4102d4e819187fd0674eed9caf5c3d5b5e494143a8efd64932b6408b2358c3c9945dcf5d22b65af3cedbff42386ed2463bd43bca5f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119551d82c51f0cc25002c602d414a8e89ba38ee1f2239929cb2400fea1fac78a08b1b35ac1def6b1c88083587b2fe33191c365bfcbbfe4f52debcec6656b52c8a7a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd2f2ecd4977f87599f46ae3c944ff08fff03258fbff439912e565bf0f683b16d494b20d8fe4a0ed617add409eb517510797a9545a01cd6fe8cfc0e47b8dedc5fe7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5004fe89458fe5f08e45eb4ac93783023c02be687466b99b70f251d26498181471073c278a20a36c37c4fae7e77962a2327ef69a5d4682cd4a33c90c8da8bd90340;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15daa5076af68329a76b2f38c2b70897a86dafceb4b9d7a489eddea00dd0279e751ee2028797d87a1aba462d2d4b04ee0df1dcb44a5dd5b9c0c3c02a1039203f0e6e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1231ad3623ad8574545cee522e33830cc27b73bb34c49387ab3a69a11667eb3329f5624448717215fb034b7673390b23fea60c91ceffc65d3fb627d063334435e821e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb55e5ba60242a750d441f919d3e948b74c63ec02b0e6b5c6c302eaea03a5254c26b4dde4b38dc553e6d772d83dab5b1ae03f34db120fe8f78a86ad311b959817ce2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b814458f37636f8027e1dea4ca695c42158e20bc4d118d46d0072f1ad7bb1584543189c42580b269a4d5f10eaf00b3da1218d0557877db2ab04dde506400027e380;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce6483a65319e309ece5d4a27e7dad104bb8f101b2756c46f5a2270a18a045fa58042ef06c26d06c31306fd4a78e1bb74710ec236f44ff34cb638ed41ecd646a2d6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fe8639a772fa091f108aea12c2a015d2052092cf5389419a474af0b65a70ee1984933a44eb6bffb404a52650ee4862b63ebdc9627f675e333ab0b284889c3d47f3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79dfd033361680f586f09cce7b46eb44f4d51ab1bd7adcd6554eb4077fc620a54c631fce4ded9c3930ea06f548fae3cdfbaa70da01de06da6794126c6a010b7674d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9a6410c90703ebf193a3bba9b263a2bf613228610a03fe6e2f1fb9abd12591c0279c7b10683f95fbf6a66d9298a237f6669cd3c9d934f5e829616d14eee328b503a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9faf409f0b7ee8f5309c2989c94cc32bd40c4233f8f1ee9c1c368fec267d79d7e044c6d259cf2445b8fbad40ea846733bc091b45bfc8d4aa51e9e45f1013fa58dcde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32e3051605df2105d13d7559e4a0924a9bd17c52fb502f9e430b3536309c67b952db7991a7ee836afc7761658d77678389279e8fc506b295915c9e0d440006a1ffa3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0865bd97a0af9f31808d59e86e660e6fcd77ff4e45790f879cbed5d991f8fba1b9d85b8d3b164f8e8f34f2322e6ff5ce6cd9d54c113c19faa353a9cdaee38d804c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174ef4039d8d53c74c66b5d6e93a4cdbef2d4e04fc26ac02191e98c0527c3bf3aa4cb502179b9835bc2020a6dc52bd275ba59867a858e723d279f150c7db0045af891;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e63d67c18f669e5ed81b8d5c8616ddaf9de9df12a1504e692baf5a77cfd1b0fc4a7ac168003e93d8ccd1033d1e5854e466150b3bb36ed3ef79b477c53dbfa3a0880;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108cabb2e75f2a26c96caaa270e51582580dc86fddf84791ebdead5afe7a9e610561ade8b0531bba444c6f13ac4bd6a24b9c383a8b6440ff4cf2738d9e6eec87f2671;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5a8b4be3a20cc7e034dbeb76299df77d9fda2fdd0525e27dd53746247b0d3f33e27ec6cc1275e32bdd59bb9c235961aa97d77d3624032a66f133896fbdfe129e455;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9c4b82967e4b08baced2aa06e23b4f88a76ffad9d571b353b74bea922bde6f3adb7438adf15623750d48399c8b3696c566ae0c36fcd9c25084940728aeaa8f3e93f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab197af72217a073b4d2d36fdde9f9d37c2ab8b84a43fc5c86374673063193b8ffd507fcbaa5be9278749fc71033c259427049392fbc24fe823dc5326d71b9a6cce5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h863e34fe9de91e51e36cb460da02296579a8ebe191ed695b6e04e1b42ea9d12dcaefd90595901b04a4c1d94f2072be78a68f6ede4d21090aa004a18dbea53e9d158c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178527c073054c843f09906af1df50dec19c8393571162486425ef9a45ee6b4e8907ff2184035c8a6da2356db2b56309c787713925725357f9434ff3c79f85d96b782;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ec07ab7d5860cfd3e70e38deb1c3d3e9352f634f1bf3e0554f808c87749ab3eb1f2cd61adf4b26ee548fb2741925370f1e7c078431b955e949c42ffa80f6ef021bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1183d1d160b08731a1819861902b8021bfba346c2e8494182321f8a94706cb3bf4c1d8f25b2c4de43bb9ef0b246ce7f118bcd5fb250074d2f7bd8d0f7dde740446ac7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153c60563955799b390d22f51922ff636bfdf9b4ca57c45228a279f23a9eb5041ce445197fdcf47e6c77a6789f31f83944b7518281d42202d3004757e1d1d044838a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17eb72cb69039ec0050b43f57260eca91a40b196916f6d9c199df918098644192b2377992389d2696dc685da87d6801b5e301c048c087b26bfb79ecec2465921b737c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165111377311081964467305da5cf848f7526fd64f7c035bfe47af49a84a70b12dcfbf249888ed4e805fab986047188bceb8d61764d1cabc42c85510cae7571cb9fb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff08eeabb9f344c65ee0c867416fdd9d0a40a8447b2b1f4d2ba710fad34b776517f6d463ce23d3efaa30812c4ca6ae8b2733b5afe320beae15d28bd49627bcf2b5c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fb236f5630cb7e4b359d5b8e373bf35caa91d8fd038605b27460ff0b9cd7bdf817f759cfc974df1c19323b516048c05d6a858f39e460db8e4fc3e94c39dcf6d4b58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1369bdd034f12e253527de55ddd76673d5e5602b4f67293d82cc376b7fa79e47bf4434c8ddf2882e88303ae9314cc5487c1fd1403f5e80eae9bf356a4c91e7027d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96064dbe3e60fb94ae93dc5b16eb447db15d840dbe3d034037fea3d8d5c45e218c975f6b3caed13409cdc4d944384be14e6672dbe1b784e4f94de1f4adaa850d1740;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bd80e518c927c5b72dcf3bc52e1f11bffe063e0b4fba058d7c523df918a972f78b965cdc7f6156b67e791e3a1e4920bdd9482e2717b2705ee2a47a3242d0443aa11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18537765897241f7cfc80bf02014b080786b26af50b0c5690be6d28edb46ae62a68881dd3ebbbbbd534c7e07e9241416d9cc2c4338b1ab23ee73b839f3f3cdddda80f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3c4eb6a103ce6f1f89e5fd95d16bcc51c06e8ecbf802221f582bd44180256825a1aa7b4b8ca72253c1166057d69f9ed142d2009f74eedb848b33202bca2c7e4d9f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4349d7bff7637e0ac15e1e52b4991c89f6134ae204edf90d2e0284516e8ff90f30403dbf2ee2331aa42ca566692a1db1e848706d8548eaac04371bf45bcea7a2479d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea0885cbab6b214a0ed5566155052d4b8700bf0e71e4adb9497c5bb9ef1c15c889ec7e64968ef63da56237763e94ead75510bcc80073fcd76d9999e3a08d8c5b8c9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9398cf5a546d1cbba808dac9f409fb820fd72e06d11f5d61420b41d00348fd2ad49497fca3a8af3967df3d81e60041ccbb11552c7ceab7c66d5d73dd70cd87b5a5da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18426fff7777b1b5e48788f645b6dfb055ede1b254f61ecc200f6ec22a811e4d05edee7b7aff65970d620505855cf615d88a3f7a36555d55d3cdc211d7aa5ac119113;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10942fc18003f45de89da8326d2e46ba1d9c3b5c2c1aea8ee607445877b24c2a79b19b8bd2ac0f98d66c397d284492b120005a5a3c84ded45697fb30ec708aa3f5a0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10997cfd477730945fd4eec796188ae50079b4eedfe602581ee1f7ccd81aea099dafca6bd04610ca654cccb877f599fd116dceee57b8cc45772ec82ff09555f783c09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2056c5c8052a5dd8329e2140ecdb3aef5e98357fed00367a5cd30e14e63b9afa05645ee241583caa376bb054610976f514abdcd744adbdce024550be911e9fff55e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d51fa951d1d1902d24a0e74753c4ad807f68ae0c38cb31bcf0bfd74019f8792937dd4e70cc1dd95aada60a0cc17b57e9d0dab799d8843ef51de81b58b8be46a0335f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121231fed910f69ead1a55fc3a095ecdf9cb971702129dcb11d99ab3ca9129510a6c5efde7e7b69a74b9d3d4ea0fb57b565666486699503187852defabb9e21d5572e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65a5759494398c3c3b813577fee0176a9bac5b2081ef0c08ed176b90e661b1434939b2453dc7d47cc112bd0682a5b83bb4fdcea9dcf18f826a46d26422784dd4a4ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120a8c07b9df57e6b7131d4b5e6fc9b6a2e8cf67a674b8707842f2799e8a316d64d9847013d65173d09b25eb6f5310b3f6e6f457daeb47adb022a891eef1c7227864;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d69ad18b134508031224a336286785f648ca9f5de164bcea491e5298b9f0f00223cae52e9f43396d1b4249eeab4c3bcd37257d150de956b9b94bccb08680696373ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h455583a075a0028ed026e8435b3fd8a73bad9d005b5f442fe08770cfb0a830ba6244281340b03726df01b1f6b83c24ed4bcf39e96c12374658873c53a3cc5f597a73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h292147c645a0b3da201ae2b6725148ea0cb9453c1f7eaedcb550571017132f6adb85d5500a6f082da0fd65ec88757d9d185914ba073808a5f793b04181d95f3402d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d9c2fae391b284160ee76a42caaa4a91ebba393359500331afc3328464513c1794c5ca4e4b5b7849d7462b211400751756d37750df1e91b990516836403b117766b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125215d90e4b4de5263d72d63dc6ada4de9e838afd994583d72931acfeac3e228c71a616b25a46926274140d62fb5ae4ad0caf568145c1fddbe7c9c36c62cb25f112c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7084aca46b3b47da46c60b763ff6f9c4683b52a3fb044acdbbc131b542845379d76edacccad4f04eafe3b4a906af326d8e7cd352b77ad9fe5513a370d3a46f4ce1d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11cc6c379a1435c499d40fc5600eb007d9f672ccfa6190109e111a0f76dd0238b2cea098e4f221366fe468ec53282abb186534d010714fa9906ee022195832c7a87d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c66960a4ce0708ea1483040f79d55ec01ced4ebd7f7b44bc92f07e90804b8e67a342747d7eed5b297fb5874103a2eaa2d31f8dd941af6957046db4153d5c1d25aa70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c331f1aaa94b41d12f9db99cdaf9ad3518a958d83eba4164d4aa5c60dc15e93248395fb1185455d2630368ac1b423aaa839cdfc8474f34615d60d5bfd383d6f0ae92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1441a4aa0bb34e1235fcf6633825b82f896184caadbf533a5ad0de53eb39e6e25c55c2463c486f8e6ef0c8a2da3b8543da25ffb9c8bf328e4a7f15a1c0ed267de10c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17add0e66696ba12ac0e5f5d58790767b352d7223989bf28d5fd84d05ed7b7132f875ea9495e375684cf80e1d7f1fbc1954ca700a39a407d55750aa2505dff73f96c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d41c4ee000b7ecd7e3298ab6627ebc8ee36839407dbb99ffe87e7d053f11e77a45ed47ac542bcf62c77592ce06dc087619dc799e54c07350cc50fbe704123bcd2dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17dbf33845a4233efbfe309248565fbdb85c477845dfd6c6add2b205391f05ae53b4c3b268adc2bac3056e72f52b2327c06e5367844ba701a256fe9e643b36907115c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea5dc48e14ca7dfcbcf05818dc6eb80463c5d936f44a7558963627c80df5fee6d5086ff46b71e6dff4945f8ce37b97fd0152113e7d4cfa098e0f6e7728413bd96f4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b8477173942b1764fec18c4020542cb5235e27baacb2c0442cc649c6d5d7bb98b616f8de5f5ece47c753a5aaf4af73a2a6da70d4a7607d9ff13378e8d8343bc308f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h367ee03e0480910618d5a37c26803569280ad63322cab35b8f80251dc59c08850c5d037afafceb566e415094abd479ab87da090845319bd7269bb96fac36989a9f69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7ff377adaa1525f39860f73946cd6983ba6aeab4818b4ffd92319069da7dbe54274a0bc2b42b661b4b087868f3be6709e4d0830e0207c541e863ddb81edda73f57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha637c4803fdd6872003fafd0eb093ce0c9e95323439e44cc95f1e39b0afcff7c06a3ac4c93a1956b22df105ad2ab24cf1b6496041a0e9562419a3f54a1c61aa6a4e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9d379f93145b3ea9b5f61afdbe44bd9d376d415bf39f15ef576b021be6a53995f6bfa9cb7974aef68ab7a161961637cc623fdbd445f7c0210c6160400e94822d7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10125cd42fcfdbdc82abe54cb713dcfcde9d495a8b6adb0bf79100beb7958ebdb633c2a7aa6a1c4745a664ee46398fc96c25916235de3bb1041f0affcc4aa12b53fa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25613b4bc4cab47ec3257f752c451ef54c3a6b9c54fc80dc1ba9e0b167e9c2be14d263f4a4d77ad349d6a030bc98e8917e4c8979ef7465f61ff6fd0b0336ace2818b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b0a27e4768c0da7caf842e5aef828bb910e5b6be1a5b31a669659eda9c1c3487c53e773d3815dec040c5350c90baf89a8ac95cd9cfa6033aa2acb424adfccfc4b6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31a02ececdfb4a66fc4e906a4392daa0310eec4bdb5c4545cfd41d55e95ab82bd6bec4499ed395952e25b07b883da9c089f2edc9920c9e62071f3066be2ad1329e63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2c7c3169f4bfba96cc92f9085ee8eef8f3ea753e7fb379e91e6a53b328131e6c8e2b96f057f1f29c26e5057d301323e29b267d52bc906940fc2ce79fa442de7b5ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189d6b35b96e4789eb3a84d176a509685babf4982b8ac2fb61e9e51b206a01c32312f508220f93e4abb42034a45a94970107ee50588b893c46800cf57f6feaedd4ef0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70f4ce6cae05e7bc2f3fb9c9c281e2a7542cd075609eade283bad5a84ebdeb8e370b9eb9be547021ed4a738c5d35759ce54845ce7a5e3a35d03c69726fbca7b6826;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35b5e3721a35c240663eec05e39b9c5f3b352417196192686f89f68ea513460ac3064027ef585a1fce7b82df0a21b3b02f221d214ab8037791ff76dad09044b5e388;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8c684c33a5d40009f962a04f54912d5e8a8da2c9eb760bdcd038a9fcc2ba0458ea8349000cc593430674d121c4d5f53c9a84905da420fc0ef6df116e889a09f8838;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5eb9cbfacac925e7738281eca41019edee6450c28b918d873cf730dc1677ff0409bc744ba265cad69150744d8d9ce41d3fe22fc0e293dafbba24a285b9673dcd5d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd850f8c23f4859fc000c61cc0981e4300839580ae38798dfc4f9813a45225fc17ad144fa7f5743843a7a5901de9b4d58ab7bd23a1046af21ab1ff5eb98f2098f9f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17955fef4c7adf408c578503962912efb7887278160135b454b801240879488401f9d14983cae96f1f28dfa5803dee64f1baed9e7713607bb2b8414338bf3f39a318e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac1332b462b31ccc359c7be835ee1361b2dfced7cf6e0ade50051f46cebdbb62b2f6138f2636d4591d5109a66a9c2fc448b8134d8e54ee25408011fab63726766ddd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9be6f68623c9b75f6eace8ec021a0f4ee7cca862abd4a4ad2bcb8ff8b3ea004ba624a468ba4d38d091fd11ba39101674f0db79c141a1a74289e0bb1fe151c6643007;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f23b525fd5c48c41c7c10fc80e1c371f28b02a3f11f9637c362dfa7a24939a7da9e9cdcb5163d15c1c9be176b6e495454ce1de24a6a25a841e9a4095e5ce56a80a69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1352e2a55e11fd255290a67b0c06a1bfa11fc61af90b2b2de6f2793bc7d6d977a2522c3b65b3a59f959a882001537eb655cd9970188cb7956df9c362a075d14d2bd97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79ec231667be0fdd8fb788bd5f83759b176ee6763d8a6db70bb1a438464e3f33745c68d861a25b9903319063b9a3397cffca099b43efa9d23d9c855c2ffccaac8d74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h386e27f6f1d03fe11ae96ec8fdad179e58792bcc1ed1fd0b273318271b3df0ff32f7d82dbe6b6b1e2e5ecd1d1b1421b098829506f572db02f4ce735dbff2c2ad02cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5489a9bc5699c72475c2bf3348a88eb8dcff0c6b91c0c7d3a826608c649bc9edcf6e240aa637daadb4fc8d24963c6dfb6b5623b642f81c5c8cf22b7a3253b968f10d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143b5e7ceeab3c0a18d97beed35c1311e953ace8ba858f08473540c163e9518b65ab53fab6c980a8bfba530466493285681bfafb91d7a59f97c1fc379104322ba596b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde27607dfc534aeef9bea8e7d2be04aadec44a7870fbb5c1584d690882fd2b267a2b72684af0e2cbdf0248d4ab7114c7675241be1991b796c6934ef238e7b38e59fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11546ed82acad47d3a2ea8d6bb658ed8a3b129037d2b20c971b8336a56cedc0a5a233f2e6e287a4e0ee44c55a26bc7d887c57b87013de2d25d1dc2cbc97126a56b766;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d605e33889ed2447cc96ad6442265f251ac3c67a2a2d42f257364a4a9ef3b61fc50e7abe4fadb8964408e5fcfc35ca1c9cc269fd7bff8d1ea0cfe56fbaa80826730b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he79f48e530aec4e852dd902d19265305460e3b9f543686066e86d67e4cbaed46bf4faadb64ba3a866d53b8d0dd29a73129d656e4a5063fee9c2ca2ecc0d0dd67269a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7653ec810df6706c01e2c4bc1b50bec474bcc18c00e31be76e73cae80734d91037e165bf1366e27a5fcf39493f7b3a2135e34f1a372c6ba5311ec784b4c1c1659c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5d664e333467bfc09a2ca0ac0017e50ff28902b5e5f61937bea90fff2a517f33688713c77c5832d7e2eea8e1570f460c6d4153e63f589ec3162b5e760473d67d027;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cef8e1cf29614f70f1e49504630dc668840407b7ec8a8c1659f1a7db425c4b03bb6e197a313785baf83e4d0aee36448a88379dff16580fc0a401bd478b48af5ddea5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h405196d024daccb5497e31f4a52be517748569d35fe51ef5d8b2cee8dffc1af214ce9e114e2848d9c26e9ad4d26370647dc066924c4cebfcd8d9cac0772249e40ef1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41572ec260ec73804380fd98d19d611b39c0b08d8e0f3da92758f99780c6355dbf7420ebebcb542cc1db431d0713e40159b55f242da4d6c9acf27af39ffa0315fce9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106c5df17eadf049741584b66941bc8a1faa2aa8ab6b5897dc7a50c74de5da09cae888f4077ebd7a37f52edf03a4ac48a2d78080a3daccef825990f5c34ca48c18208;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a4adde5273d1d1200232c8dd18ca6c256943ae2e0f6d31e50769eb93e261df33100c60e0cff76dfb9694d78a91956b18dc0804546c4a360e25c9bf45a49bd6b5e3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3d6699c32a6e2ab783726c39a78e3c3326694e4214dbabcf0a3d50fbe7b5e10a3c9ce5fa87ba0fab73577189fd1d8ae352bf4cc5d2725d79d9bf958b3b2fc9f41a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cef2a7a7bacc847d9a3e3c94503136f38e5f2d3f6e9f4a0ec6d48635b90fc2a986bec8b1bfa8bd786facb5a2a121c66205760f0466ddd774de7cb6fe43e7c7f3564;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60537fdd46acf0e637f270c8623e2c8f42330923f271e75e0dae1d68a39dbc87e145211ca460722d943a487964c2cf39409a8840638c481cd372e3ad41303a72e230;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc5300741de840b30a59707d72d0ebeca4a0404c066bf02d6abb28313d3085176ec6c03666ca4ae5f0032bd4819e5b5b43480f776e1b0ad357043152c30388b0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e94e9b192be650202fe9abb4a32a7f54031cd1e23fd7e0e6f3050a1509a86539d308d42f86f01523e802c466f82847bac543a9709e41ca3b911c9e2a66cabe9a04b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdb8925e96df24b1170b4981b692c45f0d04349a2f285cb2637d0b987a71564479101bf05a7e2cbbc37e3b4c7e7ac064036e318b59c4afe8c4f00e7f73ff012cfa35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31024dd8808f2d88f403558559d2446a3bdb5a20d6ec824eb2122659c817c157e1129fc0c85ccb211472ed4fca3b7939984a3a33120f5e220e9b3b3bd07f17bf22a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c880e3c64872089938f84b2e6c1a986b5cbf0346554796fe050a8475ec2d73cf5c86021f8c30a11c2f1d8c67fc10ecb406b5c12d660a0b786c9ca83daf6d3ab8a26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1858b8b3bb716fd964a811bdc27572b09ce4a9d8d380c00821426a9db47a7d3a383b0a47e0b158e94686765d5b4df3104144cbc7dd465e56e84734007a2c814a94a09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e19b1e92c63e3fdbc1d8c739815beb33af7b813d99b10434f7412754d5c80bbe9d2362910be44360dd0b7fb4c8e981bd747ccf0449ad4f420bac845792cb563274da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2de94e2531d547b64175f5e8e6c3db23d8e5fa6333b73b6b601e2039f1a32cf549e81943e5de40429cfdd1fd112bcb7506a64d8e0af4848e11ac953d5685d79fe47c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1503eabf2628c9e7f8fa7ca6b204420119a9ace55bdf2d3c60b72ce20d921a33211f380b67ac8e134ca0bbe18fd6be104934bcb2ce0a395ca7df1632e5e290ef27e1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1361c6b00d8c88e5856293640705311030562652f537d45765ab24dc693b784b520a7d4f357ff2fba8ff92d75972038354a2a73dc7740ff61a6d38891ee19d1c16bcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ef1763451f6781df2de85869d921cf2bc4fc50997b10d484fa177c0c581d039d83d46afeb6e3c081c6040288b66912677d7cecfaff7a71d50d12c5771c4164b8eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heef29f7793a36947679dd29c7b6131b0acb1d4912ab136232fd1a795712085a5702747f94fa422730967441e01f09b415c9ce9ef6733e33e73af7c2352f2c5908a47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d2ce23d799793182f19a31c5067093395c395cca33825642690e55562df7c92dd90362aacf9137173e15f7ee013375990da31aeecc6858460c257e48e8ed6a6e4fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b64462aeed7c7e90713bbfeae64b43772b42b3f18888954943cbe431a621bf3ef557cfd62285d1ee10f1005cb5d810f5520a63c2ecefc25d51ad8962f371f8bf34aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11de462f3da4c3b9067f787b0b94f0adfa15a113d6e7f3c9ea1a7703a1cd9d09dacfd87ae60075ff6f9290d564aec5a3ed76faa43eca2586b1bd89016d24686c175af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5de2fcb347e7d92cbba07aea435081a0b53a1d71a1ff4466d5ca26c3b8a58f24d025a75eb6bbc6674c139e5cba1a42ea0520ed15711b2a62a4d8e274e81ce0cfb07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17215d850999ddc3d5ecf366cc56ed7a97726c492001ea8041e3d3b0576ce11a22f3842125f59cdba72e4d2cd17a167ab01381a54f9f5893da5435feab5da570e8b05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf553dfda78d47e4b684f25de4967d209ce5ba4aea4039a6b79608c3220c4551974cb5ec8a919654c740c14fff32f3346a8cdf6a9aca02db47e593b758ad44af636da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176308e902a5cb08bc5826e464136ce824c853c7e47da9f92f15c180e9c839a28a52cbaae2ee7617e74281b354b8a9dfa6b0b6658528936473ac555ef12844a18d16d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4caf61c89e876a8092a62458e780a443e0eb93bb4a6881b93b52a91f6bc814c27233cf1a07ed5e01dc4dd0d0a2fb08fe600f72b2ae72cb329c1d9887ed2007ca44e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196c6d46886404ae35fae1851d5879dfd78cfbe4292dadd0f12c08d12944989ae471d4c8abce9b0f165e95e1694f63c4c9d11df25dcefe8f35e81694dc55d85162381;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65bb811918da751fa0bd957ce42c26f40e20172b77c5b6579b44a2b0270e0c7f8dfd1dd927d8bca1e4f86170854db77a2be2cf06a570de4a6f81caccdf6115fa625b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8fe96dbdd18512302251f5f04ec177c4db2c689c5d83f371856ac8a6c7b5db4a61382951aef4e48b7aedd8e51da4f6826c0241b562e4d3497c69ee015c1c77e0fa2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7ad7c5bbe4d6863f5bfa4a8fc5e12b0f94fd944608e76d1167059ca1622d238a9d96b1a248974f3c4e80bd8b954ac348cadbab8c28943035a7f349e828d1fd1d936;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188a31b44bcc2b01557ed9a09b8912a7c45e52cb485b8e8a6f82adc7976b2ae46bd923d0ec2d32bf95c733811c1160c10017f91d02f7ce63bec85bcea94d393563971;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d2b8504c3a57a903d02d929d30ef9fd21003e66f30c4c5b51368c39f6645f86dffd461563991461192e782e9d7b57f27cc99f5d8009b7a601b56dc017b3af29c01f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113c20394a77d094af45dc5d78f09b31ea81400c158776a597b9cbc498ab5d8fb29afc1f2367a239b1c942d4ffb5f9c734d82eeb7cdfc71e991d74629ad46ba1f2444;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf98cbef43e4d2319f1f2522ca2c724905cdd170d2abd5cb7d6ca4d3f296db7e5a7d354d41731c242b54ff4f33074e63fe7c61ab28c2b5e09bf8d9504c07ee3dd9036;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6732124fc0cb91452386ad5370e56438c57e13b469f646e1e55ae11391b47aa90fcc026fc4766c0a0c394cc8d5960e9f84b0e7b2e576b89a812ec9df4d010e0e644;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1048e01188af3e2de3d5549b5029121194dd21e6154faf966a39de1445540cfafb967a16dc1ffd917d85d96b988b168b627398a3ce2f3804ac99629403a829c81c6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bca90bf585e8a612e9ce598200ab08a068ac198be2c15740fd8ed24aebd1d572ada81dac3cb222ed2ffe8a0dc5e835532d77b44790eed170bd6893d80c3d885637e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1041c17c5577ddb4fa866e13ca788bf3fd3c499a3305aa8d1ea9b1e088aa107c5e91858ccf7b8b1903ab7551553322e4c60d94ddfeeabc92eb7dca3f083b80577db9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151b7282e66b6603a75033ed1a748bc72877b1d897e3cdf2a6463954713a7fcde24dc4434343183b0c5c5cba0e6a06ef240e41bebacb8f7cfe43b69909dad3c37334;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ba3abf1c3f252ee77ec0c5eb72701151a276e4ebac25caf4de3321915789bace94f3bcfe37918835eaa5d45b5366585de8206064b714b38fd31fa5f2069666992f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d9527b653014fc0a2fa27af13e6bf73d6d8eec0856abb8b6702779fe490698557d7e9767fde2937b42a108c93d03aee406e6497cd9e15295e2342bd9b0769638313;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7f7fa695930bc62905c3b13b79beb2f91d7b959b7dee59a1193758e8b13d8eb35a85a4dcc7ee1c45c6aee658ac26223efd14972a09abda8faecf5bee48a853376b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h695c438a97ad5b3bdbcfa00f3586ae2c7c6f43538fa2883de5fd829c8913a8259c8da022f824bb08f734e2af0b1b55f28577a0db75bb4c4a9138bd89e20122217927;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1640061e55b69ea39476188fdd857cb152f609d4958107c6c8586c7e0a3357b21a0b88a14788014f2e39e7edc21a5fdb761d00925f23d40c597b07c9b1f3bff7b9c3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8b866da279c0e491a438075dbdfe0422d5c1f86dc4739d56d8adc1692f1b644153d0382550fe502e364981b34a415327ac69674d4abb371e9ded6a64a6cf955af6a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h665321a25276e259d678e08cc61cf2dd19b28952d39596a2d097803d58fda04619e0bedb04eeb646e6631a3b40ff6e95deaab7463ea54c20c13232e4607eee9f18f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41b081e95b8f130fd4a73642113a97fdbf001acbaab4b867bd4f58e995826ea6c0db0e01934a75a62ed0b4f9d40771dea9602c56f649eb91ff49d8fd423895f5aabc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab69cd89a501f26174a4c258caa37f2129db1199b4ab9755b62e113299b0915a8140aa31e2660bf6860d9ddb7da3f1ee151bbe793752a8263e9b6e83a55f7a98fa8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7dfab5b207ce1b961cbc89f19b5d2a2fec4e6336e8167abdc9a686a3370376427605dbdfd8a857a6b16504642d8239d47f6b4d6ccdae2cf129a16f5e941d98d14483;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h959086d7d4ebf101e75fbfd5ce70332914e1d805245d2236469a0b8034761888c82f6f153e689803c0754f4676372aa3cbe0edae6f0eea665a1e2265dfea71b93aa5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e75f6f20410f38295eeb60dac957a321e5ec7cc135f512e95e7a1c51c947cab80f9e70c103c42e6cff5ccf90a614be814fb61fa5a45ff7e593b7f805111f278bf358;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bccff08d596f07990a0fe7d063c78542f41ac2d8eeb9e796a74694c66541985015df24e293f65b74a4cc4926da49f351999adbe7b0d8bc3ab20685ffead688791a0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de7b98901d4dd7426d9d9796bcb5fe20089425e973b2bb78f593dd7510de1846edbb3bf66476f598a08c0eae4d891bece5249a9a996dc0d5ab2d57a00f82215655ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cee4a854003e03c1b48282c62d3a807eab385ec2182ebc2690648b6ac2be6d75d825daab230b3ebdc955479f7d3ec3e215569570019edfb83e7109a023cb8a460cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9136a35c79286c5a665ac6a26cb663fea9b7f8ce6fdc20bb5765ccd55f69d10f6cdd91aa92000332781a41c52e43a4a1ff2373f6cbc775da1e08948287e3f6b1bce0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb47603fd4fc99363b612528c81c9c57c47c89bcc73317cf254fc5d586b5d5fa567c6a4199c8d78172d8eccda4d8f6b014027a2944eeaf70010288f58d5e4865e6b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143333b8aeca3cbdf1e14fc60a6156c4580f78647074eeaa12eb73bca444388b3356bcad327d7a84fb05858ab31b768b94f9a75d2d1bb5865869476fc21d577fbc659;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15016b1b64886f2284c39e1a86bf0e6a301ebefb3c44b560276fad91daf59c41b597a049a0b196080a2b1285922b8e88f3924ac4f21cd730e22069da9c11532e80683;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0f9e75744f37a2e9dc2fffc8b7e1f437ac1580d5b921e482ffa102f9edab4a7dcfbbd1a4457bff89e995d74104334bd7b7f009f72e39e256e9b9b93a420f8b60fef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166f9f1bfeaac06098a3354f02cba54457b0f6c1808dc79bff5ba2d03ca594061a623edec940ede033ca3f1bf8888076de6c1e429367f1f1f7bde881de12d9f474bd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7b69f7b2c569943c0248522e44b7b0e14085517c01edcae5161fc475287ef71a4ab132eed9525e5d99601750fd65b400e42df6d2d46ddb870bdeda79acdb1273dcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb87f9dca67bf62641eac8cdc4cca2671be4096bdc9927f5940b2a746240784d00252d9384e3d798b922879a5487ac6232bd5a53b09d9351255fc5f95b44f58ce960;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d0a62b5858850f517f4c126bc677f88491f94b8837c5e0555752e3424681b4e391d470750c13a06882d13773c8a1a1ee3752f0cdf05cad7ff30bc922afaeab925ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eea11041627033805cb222bcd969f4e053aa08d56ac323f96cda81cdb2163d18db51c71596f295f58af2586a0fe7f5a91d3d8faf8ff1b57825a247ae4ba11f35ed22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d431560d0f6698b1a31ffeace45bb91838336abab1b3bbe14c65d8cfd07e130f7bbbced3ad83451d792ee91554085edda28bdbfcee49937ba4cc7798716b5b16959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h836312e98ece9dc36b942820b4a1714fd52c7bbd3f330944222428972950faf1bc8a572afe22cd78d54089c85fd8eec71f2e402e5346af7fba073df9ebc867dc9828;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8c5fca3fef23ccbc3b499e9afee9ee582c9e107325fffd27ef925023be45b4253a50b40a063c9c9bc55097919d354be3684e8973af97b6adad1c9dc58c091d8cfe8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127a3ff89bae4b6ead3b4b913c65372896a8240b14f94ce73702b0888f022b5960a381a31940a660705f944dfc929fd573995321c86228f532531ea478202e0a5f18d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfae7f36d94e66b67683d87316d5bb04bc5209bc17dfd9147d249c91f8c48051bac4151c1d23a0f2d295ec1a27757d71de5e289f758be7e086eac4ba70627759b7d4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118044e304226f01f69932a214c7ed032718b240c3265d6eedb41d0155ec705af3541a78f967249cbb9d15362366e61ecfd94a5f3007891350cf3d3d10a69fdb2347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdf3eaf0eaa97a6f05cb36fd141bd34e86365b87de6b831245a3d1c6b2894329ebbd90b1e34ec96085aebf04c6575d391350481216d323c657964aa41ddf63d17407;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b8e02f163bf3e0801f992510a2fccf05c4f89f0bc34ad018b3020c2d6c1726d69bd148a8ef62fcd68c4e317ae84ebeef64794998a2235513ac49a03364c8e6df9d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0305ec231308a107155409eddc879d0c37ff8e84eacfd472f7e95eda104828a748c5a836d8963ac0250c3e9393adb49991d0ac554ab2bca1328f4e9662d8c4b7d91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d12498914c7650627626f66b12a00ef5aafcbe064b110c482761a931171c6a7155b6cc9ffe84c848b6ef11d2e62de64b64c3da484f0814c4e37f0a09762a8b74d6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eef89bb7b45e71786f6fad8c7689bd7b4918656e76e515d80e21614bd188ddcebbb6ba8ff0a516609730081b2ff8311f0534f6fa1d9c98409a626f079a6ca214a7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1771eef1813d622694c9bf6b63c41a82579fd509735412b8b50e4c94912feb20e9cb1c4b1e5fa037c5b029d752ee2481cbb6aca3e4f12c60f8ca4f5f9bf3604bd5eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112fc23f9a462a329f26a4165ca5c671135e44d8cf04f2d0b33ee09a957592987e990e14619b4d910df99b45d74feae3b4b8671afc0afbdb0c2044ed1d8d3c24d7bb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb0e7f2292567d5675163f1e5766ef68c29af0784c653033f23bb50f655261192a84f3de07dbc85e044cc1e0bd19b9fffcc4213453b1d72e56766dfa003da8835981;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe9af4005aa6d515bfa189cb06e0c3b299e060cbc20cf8e26d1532ae8e2a40242420bc35b09c5938d304f9ce5e1d513c92d443cb44b333a9ed79aa15b02b7d9123ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d84e9804bb9cd1c1b4a1759bb420402471c92230fe138636137a6235ed7cbb8505001b5c7071a9bc3b23fd298300663f763f130589a137eeffb8f9d7c07682ae89d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1494704b8e7159b818834ce82d2c553d2a75a7e5e545cbcc6f36e51bdb566c2facdc97880ca7ed4f3643e3c4ca62eddd75842520e16999351534f2ffb3545e0758726;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1343c8549a95b6e16b1b9e0a56a2567e709199d25d90d88c03089d8ffb4b0bb072e75aa168d9752d3acabcfbcf4ef710e39431b553ef4193ecb8e0610af76bbd45c42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18eeaddf6fd74432becfa21f9739aea0f1fab0a856b4886f255e469be6a8192667fbf50d9c60e30e5427ab4202adedb739960e9367078d88332c5a9d13a8067e48a06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3286c08a00c1a14b7d38e1d8580148902f8e85efddb9e8e5f465d2dc1b50036738815fdc69bd1feeab351e8ca0fc6fa8408eba9e24464854cf0e34c8db20f4ab5f44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef805750f96bfc7671a5281eef89c63cb75220b545e4101a72b79acad559f2e1f3f4d02e53cc4b2adfd9839ebf2aca57a5b73054942ba47dc8f1f30d76e68c6cc327;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121c09915ddd9d25e0a0fd54146041857ffee7fbc1cb96ae6344b855485965ed05379db95d27c55d6fe51b47ce2e901c81aed0951b30e553ab96b46002c7f4393a9a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90eae55e200ac1a03f6cfdaead90eb4233c2a95c883634d59ffa180567be1487a43680451d017e4bf2b993ffc4b977a07ccb7dcfc0896075a2dfba369df9a19ab61d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61c0b7874502b11e28995f2e2f6bd2bf7d429ee0769c846d7c1f12b2f7c2a4550e67182a9961fd8246652475f7be85dd8a44a7653ddcadf8f36de5cbef8429b24eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc286b11114f715bf3069d9c2e16b08c4dc8677b6a9723368adbf07ec59987225cc274c5358e1072581d5cc0515082c762d67e89a84fd2bd190827440db6f5d977a3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2207aca1f589b423a924f21c4d563b9c20c94984281c43d9e7db376c27e3f23de1b568954ca12218f2ac1459d37a1c50e4d1a689b3938968e0799f08b59097c1c38c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed65537fcd14cdfa692ac85880b4d78410e2a09bd6663a814d00e76385347cabbe35fd18e2fb85f59fdc7f662c23bccbe3ae4f1f82a55f5294f05dc95384ba9c8738;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16164c70ac9de529389f4c6d5a72e6e627201727870a53ce1b174c0e8aeab3455963315d03b648baf11fc9da6c770024a78a615b5f2d8abcc4ac9c9252f556f35313e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2b6c0e127990dd1c1bdbf911d4a5d1526e594365ac25029abe5aab776b00d5b292ad8550641d9276ce5f56a945bd821bc008afef32c9633a3657e250072c587cdd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe475cfaf0ce64e07bd5d47b23ce8e9780189e44f5411ecf9e72e89b193369d5dc401f81f41c28001a34c3639af302acbca9149ad2f2349458b042e76362462fe0a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf32db0bf0b6a9ddb912bacf9a8e2f02e7f338cf219426c4211399cfd5e2686859c4b392da004d2eeb687079c03c7e50e94d95695ef84fddab2c209ffafbd805415e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde23fc8b933d499cb599a911d1e405bce647438e690ea921eeba0bb1499cd83acfd0de463e5eae6853d6ee7bcb33e7b5cd661a4840acb532dc0d3f1ee19a4b157a01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b078bc90967a2b04ead68383e9f769cd2e8477bd4c681c8d27b0a3a21b0872b1cfcf3891cf1e05e02ef05a31d5b78043eb886168ce49eb2208453cc7f58bf9e2862d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2b29635acbb4f3a2390c424b9bf378c653ee9daed50876ab9a536705f35caa17e1923435c77af5dae9e6e86bc9903946cf04192bc44bda62baf93323af845967f19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9aff1b992bd0b7a82411be7bd2cfb7ba0f33ec512c6e188dfbbc656332f4894edfcf6f2851a2d9dccda3084b99d458a1f6479b0dc17bc9731382b3a4a4607bdbe20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15dccf5a6d9a97b3aca6ba7435fbc9ff3037e614d035fec122d0b4ff78f55bef09004d736345f8c2f4c00f76f0a084d266e067f578793ebaac3ab99a3859d2c4bfba4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa53c7e6c31327cc79f92ea415809eb48a2fa49c88ecea94efd38ee3376a850725e80150b310842fdc09f2facd135e8943a20415439188ec4bb2e185be74e71d6a2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff6da016bb1499813f370dfc0b7ede9c6ea94657562e35bece1f36199387644fe050a17506a4e2a9a03d0be2ea4b2a81bda11eb328925ea0a1c6629d04f24cce26a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a3fb85674e956f0cf95a09f581f8890a5665c4dc28e5ac41327e9ae753f68360c1358977038e4330e166ed6814c457976ae76b442524b22123023786ea4c1ca4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ed0f3b5fd88a802bb7c1696cfd360ca37e14ab9b2078d5f7429349a7ff7ab74d22e173752a391b83730264ca1f9baa3eb01a87c403e132d50e5532d7585f321d912;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac46ef733f3bc1f7921fbf1f7a54d4c6c59c91d5ae8bdaf6c505870fd0843a57beb90528260bd39bea18775dbe76919006ddb1e5ee0a13142957608980a535b049c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haeb268fd53cf0e2cd667f62ed32d408d8f46055c52eca7e5479fbe128a5cf61c06d7f528a41e475d2eb82150175fd42e015e96a740c806c9ba02b315618dd81776a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d6cac027fe287d99fb0508525f044105aeb46180c6d86ffe2a7cf1df10d797d273e99936b179f8fee79dc06b9dfad785046823f5ee29011249e5d3050341f696252;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dbf3c97ca67871abfab6301072c4e3dfc18a71158674e4900c468ca8c0f33aa829fe9dfa4285d750934c2d9cc235b100b58bcb584635caa43fda7095e02beebe2491;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1838a166e098fea2a838bba4b6f70c3011c02a4e27d91976370c9493a575bc94f3c122f0f9dd0373ac5ae25f22782335c1f6521202810051670fc7b5165431d0abe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62ea1a1a733eb444319cea122d2ddf81cf818fce6045030f872cc8e851736698386df45171b3c27934a7271b9ca5ca7eb6f439beb37e7a9e3d9a9e6e765557d201bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3a392226c708a296264c4b230bb1319d98f8a1ee7d85c20c3a11b1e61c180198898efd1e64b5ddf559b46899a186c0c5f9c04af3a324ca19fbe96cb2d1fb93d820a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0fdc7062a4979686cc7201f208d2183586d01243e019cb90f6321f33c1a03834561bbdc0820bd320069e8d4121cb24af16e61bfbb2cffa9959a80cef937c04147a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb6ed5f51fcd3ea81ee885a789eebb13e54c8c7a8cd70c0768ddf64853a66964782abd30ad0f3c373b247f4af8237f5195901683b2fbba448909a295d87c8f359c76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdc46ce94ff821e82f1e98722de9607752b80354a372c04f800681809ca783e59665e6df6cde4c76c23d026be894f47b6df404bfdef5cb430a569b7fd1afd5c2045c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffd7a003363aa90e644eed7984be7e640cc008930698e2be8986e54a1535c61d4d3d214384482c7ba110c1afd4c598aaf1baf18a559807ca5ea48e3b8aa3c2ce5ddf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcaf7cbe562d6722eb0ae2ec1a42349ffcd97f2ed488d8a93b9bf8f8568a717e38a8e51e1ba1b24c6c8281b1f05b24e0a914310703c70cb200b18e624472283a81d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a1ea7e7ec150e612ff0b0eacbbff77da1df035cf9829b18532b89ca6cef5b45825cb60f1d8334a830df0166598e3adda52951ba3a5812363f5ae084b6bc94ca829a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb661de2b518d0806df6f68ffe187c6208f748f5d0b5e2a053dcb3bf62f68e75bdc0dba3e2fb2aef837020e4471cf73cb19da3c2585861a49baf1a8dd90f54ada36a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144d2b562b4945676cf80a6ffb8b18851644302ba10af6cb389e10e86408a9549b69ddfb4917dddbd79fdccec2d5dad918e70820e413b42e32d56971cafd0fed189b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h723dde11588918c638193d0bf065a4dc2d1a4a61a1f8a1486f83d555b6dd6b1b2fef2d3a95e575a4d822525847d9f028b20c4a3ff7901b56d10344dcac65e5ec2456;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h314a188bfeee0655f0f3395871b1a6ad1755955c3331d2013cf1464821d0d83a7fec4abfa734eb2583f2be503c64af44ca65b1f8516e668040d59c94857c3146dfa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ecb87ffca5627a149cff529acd993420c854f220443e4cc1488a357362abd3c11390fade159bf783cb2c6ec981159cdb022b4473886490d41103a81c47df39c2459;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83904d76f7d02cde5d734464669d312064a480a73c2841023e9d4af1cbdd0cf54a6a98d66716b50cbfb8e4b18c392258f757017526f595275b51b9a590d3a63ebd47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1959ea7f1fc36b5338715d8b5d9195c43980b3cb82f118391f39e3344061ca5cd28150d237f0b37cec2cb6fe8ff569806c428afdec023c5deb6f3d13d4737279c8e03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152359382420021cabd7c7a21f898154f1782e35f10166804cdd15754400ac7c4dc9faf957af1c2bd5d93955030220fe8b450e10d514d763e883375fce7d91bc63fa9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14250a9f7d0793987bd3e88d1cd1be628837d62cc9938225e12343e5bc7a00a2f2739874944d8c9ab70c39f15c0cb03780b8c3136077823e1381acd689627750232fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196602987fe5255908c60669691b6ebe59e4c6e382b780f8a36c1c2372e4e214f420147b6bcd45b9191aabace64a2e61218b5401594b0d865f04b97b9b82eeffb7dc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28a89f2657384df95ee55fa2c0835126d2d409122408935e7f0b119c8975d1adceca53a4c768d503c3f15f8188aa2d02056cf474609f90bc790e78a182adf7a6d26c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd0d58ce1eb729d81d6fc1b0bb0cf2f3c2b7c6fb5112d90d95804620840b99c854e37503427e476aad24320a457a60f9d9e7a8f504108a63cc12e4f49eb2e20268f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4b6818854c0480e7c5722e0dad76627cd956950fd7dccca6b0940ca2ee663c52a57ad11d0f593982eca1bb34e41be26d56319bf3f8ef533f80ed3131765b8a06790;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24b92d81802e07d04cd2f76b44951fcc345e072fec08498b75c9df061304edc582135f35b7760750f70845d8819f865534b105009103ad43c99db03407bed4a4720b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17167bd2b5ef3ae11deacebc4bc34323f0cfba3c4284de6532080d553c8ff532aeb61ec58faedce0738cefe8f9649687be1549b26c884cb0c03c0fa55d98623549ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139f00d95470ca25feb66f2b51d297d7a1682cd1910ad99596bac454094556e36868dad52bdfdcbea610f640bbd2a2ebdadb5aa8407c9d3ee3b99d81759a5599ae519;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16bf05d537578642729a2cf028de59ec22a0ba160daa24f7a6f82452317a615187065544f3cd02e804a1d5ed8fb9bdc40bcee67f4f8d895d0d2c55faa1b64a67ca8c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47accf4721b2d58157a54217aa91a927106127f37e2df7123619858794badf51576afc877f658d96bd169334e5b375930e2399ab49ff0e96ca8143a94e7798fe9680;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f372e98d0dc455264cec52bb304553c18a28a71f8c115a09c67aa60c3f4610654f0e718e24e776732e5187cb1957740a1fc444989b07f9a19adc2ffd8b5986d369d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37b85ae6a1b64aa8e9ce6b5ba406d358c823baa20cde3726e784f80e983675ee16ea30428d97400b7a1dba00aac896b8eaa12671aa0013431852bcb205383f9d2bfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4af573d553346bc075290ef2b681a600475e8a8c2ebf9323e028e77e112c5feb448641923eb070e13a6762a91f597f8e364c0962eeba93e97a28a10489307f02352f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadc523f22afc02d8e9c4168adc476a09ee13f7481fb9de9b5cbfc9273d2dc32a5716f9b4c9290f003994019ffe156f8956a62f09e6cb98467ae34b3caec3439f18ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff06bcf1ceba54417a71b51a0ca5c740550a3261c16a517ec00c85078d800e110888e2f3b93ff5d400cf608c7b7bc3517e4c65238bb2d201966259fa2afd514b5d42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98e37c16eb21ef6f0b634069be675a46f8c37d0eabfec00f958d04f466dc9ad67169265452923c49bb578e8d4f28c45309253a6bac8e6f4c7204acc72e1a3b4279d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f81e5b1a31751d3cf9e55153b444e1a7e28a22446da9a32704eccef2d513e9bcebae4aba9f8196e0e7272a02738ae59969135b4c37eaef9ff33180a94a76d2c9e45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15957117d06018697ce9b45497d4993bff89a898855477d8161d0132a142a154822a67198f609a3c697ec605ff2970923b0d6967a37612b2f9f0b0533daf51bc78d93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7962825acfcf22d944da065fdbd3dce8bc7f5ee4c55984662ebfc1241ff15fb5db83a65b7a343457acfdb9419d89beb800181591c06161034e983f358a97ac0f14f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6710c8df096639edee6b4d9c5c244a7f5954076abadf5a7360bcc6aafc807c37e3dbed0d258026b8dfabf28fbc787478980607b6a277cefb5bf2e46cf75677e9adb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9a12f18cd1e76b65952ee4302dadebce311ca82d4d153c1d52cf306a529dea45c97b534f59fb30511e1346a50b9b8b509a9360fd468da57997978e18e87eded9074;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13464e6193d8cea1530a1b93cd4585dd54e53ec288454df25c01bda453c4f6bc2494b45678d1136ed3f360f2205ede7b56f42d037960a43bcbe3590bb0ebbe1c76d4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc3f70e659d87e58333a60ae52cbe787c5e38a354eacb777da829c19e9c36408e1dbca5e8a889866dc487e19e5634d079e9ab1daeb0eee3e6933b10b6cd7879b3d56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74b73dabde707aa1398a8bd0cd59ab602ab6955450ecad918359d334655198c505665e1f4d71243a1d3309af6bce7f90a03e69557bea198285a5b2f4680440989af2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1251a59098681b797cae8a46c6bcb67203d18a01a09ff4eb207b0c329b74d27dafb5510ecd0d47ad3e380fab8cbf2ea8cdafad0703963a0e0a1076a7c684dd2469c93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1accaaaa09ff3e2928955e649f9723ad3b5214073f64f31b4740f204cf360ff051ea3e2c6cbb642110f6856ef337544f5539d6c446413ada6df2d9001faab7d60752f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h487d0804c7187ba01277cf74d0d04c411e15e0d1880d381c5545fa757741c55050c1fd45b73a76e817fe220d688c30df573e5c7cae8864eb007a96849862a90158cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35b034c4b1cdf4a8b432501ae78c6b54424ddbf9ffcd179312e3cb1671a98c4cca903dd8ebebc6a74e6129b6c52bfaae2bd7aec48530c3663391e5388139f0b70cce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187cd59d4a3573fb6328bb47873b15b89c5cef46b163d481794b03cbd559d12273044b75f55c7b2af862831db3008f187824224715d2c57e955dd86df8252e99bcd98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc62fec0d1336066cc4e4a93571b520c7b0f36177aa1c678dde9195e770de4462dc6eec77265674a04afbe02b8589435ca516d933a8158d9c8ff9bdb57f1b470599d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2b9fc4004d21c03b6eece086d93ad24e106cf1408cd09c06ebc6807e7030125c688fa9a6a72fc6a1948e7ed0725b1daf9b09a9a2779439b7956163e760b10386633;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193f8494bd99eaa99021a91f45d90bd582d14ab50050dcab1c68686539084caa28c9a8e84b9e4ccbbdabbe28c669a23e68453694fe5ec58d87691ca1d18035598c218;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107529b318d185f07ee5b898ffb57fcdd2f334931b26bb258eea453e342c3998b6e671b660e7df35f268a1b7f870aa7a1e4cca5b67b10e99a7042d14d2cc2dfd48ab3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7ffc7fc0a695471758226e56d003ab65a8259507cf6d7e69f52cae7201426813e393e607416ab4dc3aec90d94cc10a727c631859e345560015628796f16c428b649;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h905f3c19f296ec4dc7afd5f7d929ec147126efe33596f773aa10086633e3a0b85463c0ccc2bd620b62fcdfdfc41341205bf9eea9e1e5d9f888e1de6011592c8a2d01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118d30d1c15e9982ffd17da2a0b474a38349a5293738ab76eaf0315697e0aaf18d6adad6257d85c0c81de792707d871bd4aa1f5d45f4b8c2c4a6ee9fbfec2bd81690c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c96f01b3cb8b3955b8e2ff7e800142f590d6a9fbd32f7d0130f05733ed7bdff86d88a7662ae9f65e07577187cd79185f3e5c78d60e28bdd50d08ea03196bc147d267;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70969b6e55ef2e60fea3a1c73fc8a837f45b42dab1f99abb242896a99a5dd6d834f45c642c8ecfeabeb4ca1d0fa61c5481e089f4d77d0b28936626cf977c4747f7cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b12e598038a7c2bd166a5b74e72f7be8bb8733a72e5814064b4b9b85e90468d69666330dfc958d422e37db3253b0b8c218f8c404028a40b4037fc693197b0b8a002c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ded0863206e58098d87fbb0ce6d2cd31a085b34fbab42c0c1832575099faf48d1a8da1f8577c8ebe5a76691372a2f9ac2c61a82d66daf7ffd25fbe3da07b1dac761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1540cf2bbd21453c8eaa807cb131705ece31eaf16b6c071e98701dc9a7a757f2a2f7c89b2262aa65de7f3bf73a50b3f8df52ce0d0981238988cf19aaa6e250c031512;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b2550548abf3442791f2449421acb626e0113d660aaaea287a77a1fe3daffa5669d3abcad7f591ae0cc8f5e4847bf74e5ab2c34b0cca14d67cf4780be874a5ae8e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18973edb0c15f122e237470e6a85e45f321fbc56cdcb6fb65dfca886fc7507d5c60b201a29dbfe158b79d375b2be722d6a81d79351be3d1f178eb7baf171001adbefb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ba2bb39845cd9b1aeae01b431af920c7c6dd4fa862765586cc66e4613fd328a9dd7b4f9dca96ae9028c7192cea85fcd6bf54f80fc23dd0ba0df4ef40c49d75dabc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d79c94028bd60427fa62a1e8a2c51bebbf056c81fd4783658fea86159bb69b84e7f95397d07a5a70df0b12f40a4db374959623dd70fe4f7278548b535bb90063c13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h520a289153a9e6c8e19e51ff1007aed54235cf2049548218fd04e594a2732123dab273cfde5d962fb98471e4d4fb1bfe7ed6419b865f1d1076de5d29cf24170110ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb55658f62a287538bb56b0e215a10a73ae3a7ef109778ae0b595006cbfb775dd48fda189fc2248e0bdc5f40d13e7343f397610ac9ca10d589c1f0489d9f9aa6c225;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4dcffc3c5150ad670feef933740e1190b5779caf7593bbaff9e8bf12115200a33a07382b8cf81a38effe2be56dbbb138ea2eee7847916f415d40c3b2d8ffb6e0d55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h502441a9388ca9909807ecb7ca8c7c6d508db180a75e08007686d5849da9b60057dfb257cb7815ca04261e9c434866b89aab1456c1928c111314dc7b8fbb18c01d49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8de3663ae0beba6bd23da99558f9ab5ef5ff0716e8b078629d66587962842bef0c8f815ed19f9e1d70e4af0908d68d8184c6096370f81a8a6d499e3f9e060d7ab204;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e785fcc0ec70a9b4dc90c422c1a4717733fa10c516106940e6f1d47e8c7d6c710875e7da89b94ed8f2f2a922f140ef6e2887a935dc008b5b23dcd16040bd3cac6bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1070d465750bab6c564410d4ed1c92324d199453ecd2aab062d47666d561d6602e100cfb51bf1fdc78f2696d5b48a08118b8fe92f32353dca70468c3b6abdfa0807d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7c60fb06a08ff718da783b4b2bf2256bad8403d0cbae013a95b29d3665ea08bba6992c50e4971a700198080cdc5857035262b1a0d680ba68684657670bbf6d4470a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e183a1393ee710aab4086793c2913cb28ff13fcb6b14a25a154c42b40e233f9b86d359736be4504d4fa8a70c2d54c6ed1bec6236d398ff886844f44664fa18d00e60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1619bc52e8d770fbbc440b523f520b8f6b30cd748ef839329ce0044366a1845f7f3b7a796731c8af2648f4338669b1bacbffaa338ac58aa0fe230550fe5e3639b8175;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d81819902a8f7624987289d34015c6efb468e0ea185de2b5f81f87f4508d12f8ef4d039d908359a26934d6f104fbe79108e379ebc7bbe7e40a8d9c8190be6a135e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184a8762009f610ffa86aad42a2238d0132441a48103f16b5420ff7b7fe43e9d4718224edd5743445cf91fdc516c2ad8c3d1c38c9a1f058ed9e8467940c24f04a00c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd6f4bcde429f5c5dbfcdc99b957f1eef9d36e8c22734b058565ece8a2d1fe3f035f39b453511d99282ec3e5c8b1b996edbf6d9ae0675cb21c62825d7755adedb3c26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161e3d818c2776fb11402109ebc50ea1fe318edb08b3bb49c70adf9f0c8bbb264c03dcfb8861df36a79cc263b96006fbaa4aaf3d9cc487d9f44cc3bab91ab7e9c93b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16193c873110920ce5089cb6f164329e987c19561057ed7db5039f1337a22db69ff4a2f80def73cff63485086f859bc5af5bdf7d4c20aa3e8aa3681ea508b8c675103;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f22e6e311872a6535de3d7c3b15a340aa2cf875ce4749947e30abd496acdb509b71d9eb8daf724c8489a912552f22624b35479958e729b9d77cce7029ebf407f608;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10dd22717bb61fa51fe82035bdda4d6ba5c12dc294c59722453ee14db3f28ffc086e4a23f4750c1cd1a1d24bc07ae41630f8656326dde48908a163fa96549873770a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f561a51ceddcec91faf52b25cab0a8f80264ac39ab8767b04b6d0a466c6072c1aecfe2422d299b86ba635f8a2dda8f82c48e32d4069c36a7bad90c966f1ab87af25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f80392e7a3f0866dcc4e4a4d2bb7de6809cd879dae5546144b808fcaa46f9b4468cdbcbb8848e79b0c8ebc98d34c0f9f212e5ccd2da1f15868256a6e65fa90ffd22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he89b23fc3270e6bd2b6c69aab4e455f5b70ff35fb5ecc671c8024a8572fc324f5352343189782ecb469a269ce170dd0fead6b5233cdf3ae3af8bfb4251dc52605fd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148c5246bcbe3b494dc6afcf7f24bb315a9f02dd6cf4d7bc5563c76f2e6ce8bc52a57a5e7fad63cf166c0e12979e9680aa31a7426efb6e55c21e66569da443b8ed5bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192da2da51449c55d554d1825691768a17770b8b17c30bf6e0a6b89e3dc2b16e3071149b5dfd1decd370f5c1cdc65f78d8599fe988be705bb09bf29c5e7d9a78d9907;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19eab42065a6f4132d9727c8968332191e614588eb95f4151d318e37235ece064154637a61eedb69889c558ef82749f2124969fe94119c5a155ff9828a95a45645d34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7305cfc87f15ad1336826b5fa7c10c700bd0f3af640c0a8d4bded3a4e1f1d7cad74c3a147805431d1584b705df11f21cd18cd19488658123f9444ae7345bc6c278fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h412a66fb2acf09f958057e6f808f87b0294fea2d8b430c2894c9982094da32cf111559957e13c61be7e09306bc946c33f19b9fada6a8ec552739234f93b86b063df6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1561c814be0d66616250f95d574625c38ebd5e1b456ec4891f86861816c887ddf58d85dddf514abdc063ea15fae53caa43af5ae14eb62ddd1f7950dccdc06049c199a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b2cadd10eaf4d2ef965c2da7218bea891a362566597a5c7220a955ffde826422713ed7890721604693896f4ecec91c74e587880dbb1497edfde53d01a155c209ef3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he44048b5310f74b6fc48cba6f36e9ee2c9e83427bfc7bb4f4030cff1ff60273af2c58db2015c6cb85bfca458eac7187a8dfb69327354d7e25f30c1593f442f4cc43c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc547a8eea9a9db35f9d7c2c1f1d8c5efb3eb0a1941e348685545111dcd77cd3b9436ec084dcf86178bac49b05c06435ab6233c365ee6787cf9e93d4d51c2248d3717;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f54770f21efa0db4b068c370388f0daaac567996ebcf3b32e28d503f7d330626c674f5b9c5d7b462d8b8df7a551de51ddeb546ae4abf9f579e0ede888f580b8bfdbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a50f3b450022b36b1bbb1dbe41b3b77a977dcc35a31430a90240f969aacf8a922802073df8ed97c3035bba529bb37dd503231a01f30b1d563df686469f8d9c594110;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9469ff5dc6402f6a23e40806616c61b9ea2674976bf437998a654e2151c5d572fda149212ca89cb1a220e4a4be1d0c8efde511c82075c0c5e56ecf34366652fed818;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159122c6b031efcefe6174dccb02553be023682c48dbc06424c535fcb9fd10e5469b0de7d1ae1bff96ecacfa54be6fad1f379c8d9add70752b9f13e0a3f6126230d7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h43d9621ccb6c37d3cabf0bf3642cfc3aa8749f1dc6dfc3ca63f8ee18388a3488986f856abbb007a582826adfcb6569052687c675a95afc112d3299753e60b646ec18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b2e2b92a9829b96dfce788860c508d968ef690cc52356b2bda79d7d66950ae53aa7e1b31c2a2b622243f93f3de1762cc01cb572d752de89608760261c805169294f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135c6d5f895d498abca65e9a35d692a8aa14fb563f1abe67d449dfb2592b8842fdac079a51ef0182962c9463b450f99528fb51fc0d532fc6df4c942ba759f7478dd5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123c57b5f19b998c649ebbd578057803b04343295a9dfbd7b664e19b74a6e16285f806d02a66beabeac9e0f99fefc2a807108598464c084157a2170df9558d7fbc44b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e1c7d5c0ac83b5b862fbec87a07b8ee9c22da11f86e0540ed11e3b401d71613c22348ec31e8e82c40e34cfd19dd23c2a3ad93281c0a16e390a8ed31aabd890e92d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4a3c8375575a38db1add70aeb757970cd0a4adffd17130d4583527c02076099f44d7e3b52e8c8b204880d32a995af618a898748d24eb9deeb01850d9f0738cbe518;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3fd354aa143778b1e88d54a39140bf70c79bf6a782ce342386ee1eca9c3f209480beae8b6a98267474cabdcca342dcebe454135bc429a8e080c0e56020242b2fcc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a9a7ff75a1b3e92111ee8f5175bd6a705db5743813aaa7c1e49def682c0dd2dea3863e5bcd1a1a1a4526f83812f705d7a6ad6ade47415d825a0c177d2dd3a66f9c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc86ae273d71b56b073ea48ef6a812dacc40d097d1cc33f152d0f14b8ce0aaa5e4b14bf9b1f8b46e9601fe84222c4cb2ae0ee068c00ff0cae7fecb0b5145d20c8539;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14bee9bf85ea021348d7e1108b350438cb2c1951dbbf95607037c36e62b7fffbb4b79cb9267df1ca582a31412efd10b951b25766babe5d9b3f50ae0636d968306a462;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a14b10da79ebfc07e3dac9c4eaf79cc846b1945de28c5a683cb95fe351ab14a33f73a65ef8f9c0003293c0666b5a6feecfa189ca0f01459d431d6d0d6db14c0667b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1f99350f05f19ef63f0ac771b59e531b0b03e2a6401d469717cc21e4653f744e57047ba80712cdbb6a92bac9c1fbc2df9ca97cbcf53a03b49ba808ebb3c806892b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcefac76b2508d559be0f0270607ac9c224c5e82cd9871113e448a4b5e6998f7e3e2c798222fc80fe4cdd10df5b69ca09d7d0b432d937535ecc1091c2d77f88d1191f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e6e7b3bf58c5392220cea88d4798e34787fddad7e7aea5452fa57482a1ab58c8b4dfb24f56208c91bc58d21bc420d86d9fa1510da175e53b459fe709330d153999c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146cf63a4ac5726196d611998fdb73431a123ccc2c1c4614f00ec40c7a0483c8bac52210fbded21d40f36f74526e7bb9a858c68888599c763426878d8fe14def593d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a07e01b7933b2b6ce2017d4cb3f77b34797cf73505bf8da05d5dd0d05a35164eae6ab1eba12551679f9bc94ee8380e452738e98ac782c69386940ae79c1cedb4a88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0eaccbdcb8034f1e5ac5dd492f392a48083564dc56ab17fb4f6f24c05c45c33f20520a4a6e5c4d13f6a14d142af711b68cf71e555fe9c7c3527b929d7c9418782af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hecf0dc83c345fa7cafbb6c30e8eef85af7ef374ee28a29a601a3c340fa5f3c4e9c40496b0629e5280a48b4d0e847ff85052dee1bf07d3e45c79b984df2736c3411b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h486bab599763495816f484e97a7a90350a8ff4cc90b5236379553d7960302ad6156820697c970bc1e57b646426cd9508b1aa4b06acc135e277092c5ca3a8ecd60f01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a860800d886949f441a05bc82882cfe5bec12692369fa82b2fba937a9d3b4228a6ba21fa615b7a3abebd169bf0496890b93e513c1a610393ca070b9942ad9ac5581;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5eeead4307b49c1b42646dd702c7d7c1e892a609c0101de2b8adc7c22b812f0d842bf3614cff21b6e09731001997a3d1d4082b69f63275de3c7b6d8f7ad213242c40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3609889a792f81b81bd1bf55e36fe016d8df0f3691b0061de6cac4baf5f604223444d5bb23c1de3cc373d6eab3e35b6b8431f0f87562c3f13e06696cb6f218937f7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec2fcde542a87edd338ef89c406fef55c42ab3eeaf41d9ca81ce412f6c0fb385de602b3ac5d1a809e18028caafa8e41ba90b11b28513009da8a7889a395bcbde88ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fdd1aaba744fcaf090f37fa552c6ed33ea864f19de6a7447c60d09645920f54bde2263e005502ad435f6fad164a55d268d45d002b14d8c560116b9899733e17356d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afb2663e061551fa6aadd942076504ee726f6669f761d2a4f8af293610f4daafe08d51c425316986a12786ad1ca4f80ea0a982abe750257d1d807fb53942bfddf8e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28acfadbf214452e9373c8c4b57f35a563d151a8fb4fec052ffb15cebb98de60978ed3f3da7e9d22494ba20952dcd90e3eb1721438e4d072216202c90c21dbffa837;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d484fa2b794b54f7bae11cdd71473bc49739aef36b3871c7156b4ff9c41b4f8c16b0a1d3d39e30792684212b6e667a00d05e6652e7c0de90854a629d6267d3a4206;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d52070b2634629aaf12974f42409188f3fd5bc2ec24b150b9fbc49d0a32265610045d755aa3386d34bcb9eb179be7d9732718f34e34c42176f03a08d929c0166f18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb46c46cfc39069a61c15c4a1bdd2097ccd9af6a31c90c813f45bee6049c4657a711aa305af801ae179812e6aa4461368080ba036e38577f151746899826334a42bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb275253e697f3c8b26a0dc3ecbd22206e716227d33d3c3501ed63736c87d6fff0dcb5d7b46d3246bb6d8e28dee93de50311277fa9f95bab46eeb5e2980b6341e2b8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h768aac7b62b215abd62ce6b9e2cd2af17cb4b11db48e56fd7f09a08cb3768ec0aca59ef6b38bc5c878911c53876579b142626a3f126acca8f76675c0550f3bffbea6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h658d446b800cbe5254c791a9927b50ebd45eddf3093f3bc04b34f47db20ecf619694c6527b9f131e95b48917ba84cfdaa7071ea69b4bc5fdbe9c9c52e8bff92f469d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19292e1872f360b926d25fb617cc5800f92edc0bfb651501e51084602b9a981790c3c1d0ca484b3b5c85b61fbdcbce2d8c917c1814900ee557a2dce3b65bd258d37cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b8bb188690b2d9787704275b5bd2b03cc78c6157f8a5eab58e5f1b2ca8d2c2428546d59c50edcc5bb7f6bd2f0f01e9252de871afde1fa94bffbd3ca5a2070edd78b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f46e2fed8cd0790dfb2520bda554201f59d8c4fb57db8959e461e4a63095d9de31593ca58b6e03d1c107645ae71e9c882fcc982a14f8e9985ec4259075dcb7ed8a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c4223344be4b0557554c7e370160b4be6e99bd6b978b0992aa1f00bc062e2dcce03fbb53c39ec804cf8e6be48106fd2ab841fb692a72ddd6caf080ad84d5699b8fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158d2dd5e1473800fb38119b163cca4b0791c61237b823dc68b4b6198752de5035e5aa573fc884828c43e9f74dc107271c3c6acdfcb40693bec6e3bb15cdd54f7be7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ba0f32be08508e2cce46b867fba255facb4036928ff2c111ed969f8e84ae428a599e06218694bb6af283709cceed44af788624e453abd88c3cd3f3b787666ce2162;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a7caac3a856c5e4fb86c42fee85c587a4a760080f12fb163bcf276fb3aa58fe5bcf0487924cb7fcf5b566b8c56cdd206715c718d3b425d48914d306944e981480cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c693891c4cab79fe68c330526d9b017d0b56b155dc60929d52637dd9c14fcb83b2663b969a83cbd553b57151e4cea3f7a77dedcdb535af91f057d332f35d1332005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb6ab6b3175d846d542082a0020802d482c7cce181f24580bad35424e08fe9730a51947bf848f9c3a5fe655b4af30890092b69b3ad74c03118c9dcb1a88cd3f6a1c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a53dfd6ac40b6d2913459f15e4e493bff01e0ba32d3cd2ec7373208bb97212a2b5316f97ffa2630bbb2fecdfc819564cfec44b698cf5a0df32368521f3d903126b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c14b02fe7ce57f6420d24515f0df98d9e233bce27a6598a6be639d4490255374266c0c7ecf87da73bd7a7a5f8e208af9c18dffae6bfd459c2cea3e435d37614b3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h516d6dce2cb3f037e29c9d9cb082f7634c1fe35bbf5b350b18e7abb06f456ba58e3dad6099e59830c353f876275b8c5fa0d12cf56157cf21a5142a7c79e3859dfc12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119861ee7624d10d2e1af4cefe4177ffc1afe4dcec04a6104891e7e71ce972cd01cdc959f9a5a6bde253c7c9eaad2d198c4fc73a3917d2ccc2b1bee197ac126085d9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e456d4a426c130d1672f7d1fc55788b5c2fcd770eae826991f653dfc40bfb4ec3296e2495975478e615c6e2cf7de60a82d61592833952f88a9eeb92bc8950046286;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1114300b568d651295ea78d08f2e76f86875d655402946006b6a6b1b283ebf215ac6314870ff03709f6b33b6a62b868e28f6c23c70d326e65b27e2dfde6250822d10c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15dc8d8d2763f938567ec6146de80ad6bea00f11f3dee4d5c99fe90142aabc7bdd9af50dd61e566956cc603a7d3f084f6978be393e61094e031097fe3c8b0327160d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10eb028804f22677b37ccc547cef24de8a826b9f9e37e61b0e68c97d886869450b748374d835d0e1be53e4c972e8d355ab092a1231b9831245733b20de0c4ff9e8b43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fdc8e6d3b9fa286d15e5a5385dd643ba611156de4ac9afb14a4dfe88e51887fec866c98ff2afbae984825075eebd6b4a0d6508a4f859f51bcb7c97057a091847824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1aeb72b8001e5a8593c6e92f19cd84d2f4a4781dc0b2998781fc780bb6b9468145e705bcbc8f40c5b8c7e3bca740f863b14a3d3647ef72b3fe6588b87bd88d61d80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h616c51f76c0f44e919de2e084639a6abd4cd9f2d44bcfcc52fc2ba441c3f56e77877baeb672ff1d9401699248bf02b2d8bde26c81284692f1ec5e7e118d0aea3c291;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6e5a5f7c1b05f74d7b2121b95bdf12c234b3d258c9bb3f037f321fc080c0e209accebbe3e2a7bb79a5f39c87dfa8ee74f3f7f4beea70c63240034fd60104fab4c9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180970ec164ee63700a6ebc48cf276850eceeb8b7df9b83fe3cf47aca87eca6d289fab1ed1856826b2d43bb4a96b3a620362da1c49debdf19dee46d00b5cf3b71aedf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff714d94498f2c7fe0073c946613aa8ce4a0b6943434389c8b12d9348400a4677e0734c881bc903c0dbf27236a7d4f3357fea33db940178741ae01737de2beb5d623;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef7b375c67c99958d3ba5a140dd18d0b1a5f344a344538961db29af493763f4200ea3edbeada670cf79ad0173f2eed56082aeb91d3f260f2cb487c350d4775684daa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3627b0ff50eef1b6cc7b929c6466a036e70d1fcbf30f7d12c084c264a25563f012a7d2327cc332ffd89fafdac0c8395d3a4e23f0852807e086f43c4c697060cfa460;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e9a9eda4ce161a0e78d3e9ff959bf5198eb949d5bab437f94fc8055cc22554dc90e8f9d7c84366ee64744a89622d2238fea3fc6601da5df97623c70f34e4c3d7813;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164a58c1b6959e20d2b5139b068b7d252884a9a9d7d44436977e0419291d51b1224913db47b86fd89437291ac4c85b1c32b779aed3c982d017b52dd8de9802b75bb78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d13cca07ccfa8c267b2edd63cff0e2e1439e1d5e6c4ed18bf6e27cdb59a540927ace549db3fd171139abec1c59f4e3def8174fba2ef6481450437f1725fd99db914;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a55fc37628244d84bb47c8c2a565fc54b344755dfeda667c25acc281b7f0b97c2849a56b08e38701afdd7d06e8d48b0af4dedf52baa732cffc5300b39df9c8275978;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83028c579a7a108a27e67f7a870d959a60d6801cf79c4d68001f2ca0be28b17d6e7404ae073ded071c25add4a1c917dd8a0456d23e58158534dfbf439cf26558ce1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f993b0c22e1eb14fd6f830d2ab9d5f888fa51dc2f73ff2a3c669ca33f85d32604ee1df49a29cb0dd76f20b7b4566ca1b7e34cef9b2f7893f204386e041edf692d5f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2531c18f717402b812649789e0992c420a717853d51fb2f1028ad14f12bfa9d81a460e64760c39863c513e76bfff4ecc8d4689742338d912c89f20af25b719f8c19e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96d096985b553bc1068920de8c492f9e94c9c229351a20875bee30e1e653349eb0356919b4b9363b6104a218f11920e04e4c91def48c852af78d631ed29d191c5fa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaf7f3f41fcfa2c6e256e7547b91d7c6f9d6f42608facda15ef5604fcbf643d1a69d3ac274deb4024261400b66bd344218f28d69601feba5d427e1ee0aaad50cbe2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d2779e8c4d684c63b26b48deb00c52d47051f3eeb49109f75808d20cf24ae6d5e6337d4edf95974282303192f9540220b1019a09e949f20f77600c48045e689fe56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137c9190e3fdfbd132fed5a7afdf7e2e4379d0421c33297c6c7f0e5dfeadf5b822ce1d912b5a48770f667cb9b28e473c479e792904926e5339a43453c947131588a83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186d75c73d751f909bfcce0f6c1bb1103a772486f06c8c2e278df5aa087661f0f2ff85c7ffcea4586de20bb30e2a70f597cea5763639840af9f14eb64895df8d1344;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e31353f22b7ae7fcb12242425ebbdea761e92a439041897a99789364c172087f48c830f7df1e7531764c09ecefbe57a7bbc33d129111ea0457d2181ecdb7ea81396;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda9c692a03a192e749c41cd7e8b6a6dce77f0c212dc346332f0b925f98b9cf543455a608eb4874acf84fd09c52ec1831c95bb865f586e87f3c14cc48f2718afa050d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faafbd7eb6228c704304f81661bb75fced38f99cfb29a199ae2bcbeaebfaeae6c4a5f3d95b3f761ecaaaf28af71630550a7201efca40fe1b739a4e2821654a4dd38d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4dfc4981de167a1ab9b1c019a12cea33361aff3ebe12ef9865f244c8ae0998d7757cc3eaf61cac8cb0753f94a1878b04c0f883c660cf6b4060798e7d8e87105a50d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75e6b051178a63ddf0f6236eddff6374483ab892269d57ae6aa1647104a332e78b0c2fe8132e2214555bc9b8a76f48abe12debdb60dda3fef65050264641c0513760;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd54c2c2fa5ed316dfc59b0f6cef494de1157194bfbfb4fbaa5b8f38d04a68ef09b39cf210ce8c63f71085fb6e4d5826900e03eb1aef23b10b997b95c472466446f0d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3a8129a79973a5dbd917487d86fc3b9e143ff8ab8a7478a98498c327de852ff9269913dfc2b9634e4a5559190754a4ce7dc777c7760a13bc37799fa823d5f21cd25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124f679c463737752ce496a9a8345fea4c6f5b8a104592fbd26e3cad638243b8b679d163cf2e59ca1444e5809d0a1d8eaf535a92f97cd160bd5ad4444acbb7201a662;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0b267d222b7cb5dbc53bd05f4012c15fed070a69346c8a9914415d25a6d114fbbb4af350a94ae905ce5aa656c3d60a12ebe41b8166d0821ddcec36f0279f498fef8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127b06f23196b7813c38d9234801a9e492483028696c9bc26c8dccf5472764e4a2378febce1cfc1feb57c97cb28eb77347b1e99e2a73657ebed76792ed6f4e33a1ab0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f145cc4c6e7c004c998a9d003fd360c239ac4442d3a7dda84ea7327e4a604b7e310aab55d90688fd2a5ce1f1e13be3843727221009e8f0150286d5dab660a75fe895;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61a4409879948cfae6a510e068d3bf33bfab0f27d5fa1951eb4b9c95bb68306635d296cb2c293d131d5ffd8b7b1d4b9e5961242f06fe0e47f79578a53c3514a1b791;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a4c7d7918b98e8da91b9a9c90163a079ee79b9da845402fb7c68a5d55441bdf62ac60c858b95fc97b1e21746e3e31de6e345d9503673aacd177be26884a4005a2e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18564630335a8bdfa407b5fa4f057e35c97f72d9071b77b522f652a2e4d139fae6cc67ec27c9afc025b485261a1406c246c7130e68bbabd9b9e1c589bb44f82f2370d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95b7ef3cb95da08ccb0a60f262978dd7c1461eebe446b48e149e72788ced583ed50ea46bb49495904e810cb85ad44895e1959227437ff12e5e203705aa9f79738a8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36666f67e9ea381b83b3afd5fb475afac9ce70e4c115200c84c9ba757dfb03ae12fdbd46e4a43fe23268a390bfbeee77939c946fb8ba91a5abcf8ad79a49c9c4056a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h687bf78fb1f0a41cbc746257b6bbf0a338336682a38b30e3d0a3d08e4765d53bda266ffe4dd371691404a3bc0bd7c8d2b69a0c06c96664c5c951d8a17601b80eeb09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90527a639f3afe66c4881d0c72245117c68d42695571720247a3c8d31d3456e9e6aec15149ca11bbf2da8c26564e3d3e3aeb993283370bb22eadcfb990d508e0a2aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40a5ff0d76f4642bded9350ebe032fd25672e249bbfb22af3780225ebc85df0968f00ed018aaa9efcf1419ffa0836a281efe60000a0479a970109541d630ce3090bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd3bbff53ccecd59a20560e41c9b1aa8ed71978659b845a3ad92105680a164c82fc774ecdc0bc231c25c33c3c85479169d213a24c30682472279b4c48d9116e5d493;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1233b2e6ecc706262d20b63aa8ef6efa1fe7ba3573d355440266ffc562982e86326f9510fdbba8799a417682a48765d25f01a9ff65e0553968e9b11d2390bea97d52d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd04052c4fd1ee6ffdf1cd5a66441bcb0ed9484a622f5441c8feb4b97a88c0de689ea45414d336a9be8efdb7772503a115bab20e1873407750e5880128dd5f3abb61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf673bbf97fabc9433bb6d285803b1ade8df6fa9319ef5cf59e0d811e54585e75f3b9a68d31bd609e01551ac0d0d5d5082d42e30f32268c8c2099496277d4e692dc2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57dd1df84ce3d0dd5163440f6fda1bd0a5b97faa4b235e7e0b66279614b616901aee559edeb53bff01c77f423114160918a544861863c8f7aee667d90ed5d501c944;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d2c1ab89515148e9e7f473102dd2c3852b7aba780aa36eff6307de434a3b482de5dee8047d3a33570e6ed76d8fb9d27f46ea99c8200db58aaf49c0544775f2b2954;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6f2b9aa58c70f288b8ab6bd34b22b4442bcce26a40bb8ed42abd266f66c561ffe33e08ecf9bc20f301ac73bbc80ede870fe3134dfdb406abc1d84b081fafcc212fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5edea3369dbf643cb79d0833f8251bae1c3b79857d2745babd8f6dbba5c89a032b67dd0e6bc451dcdc1793c6004b63d5b0377f75d6c779b1c44ea8260727416f44f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7eac523ccdc86f29c56b591900027dc09bd9e7396216b6f73c58690bd4d2544558f48435b1ee1fba84a70cdb1140bddd32bfde63e19ed84ee8ddf55a92685703288f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he536bcf05dadd252f6e88f7b7916bad091bd958dee28701e02d12d1a19f9c3162f955ad1ca81dc8dd4b77b8bac1f5b924484de072e14649166f78016b15449bd2654;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c322814bb1ce1716fc8ff0799ad47e70686ce4013a17da206d26e69c9cf0ab1774286e69b014d16ddf987dedafab012c365a44e0e473688294395227dcf033a086;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e71725f3f966f51b9f064d7d410198ef2564762fbacb0e3fa6a5d4fc4b8c9afaf9e40502a221e2003e182ebd930e9aeab2265d7df108f94551d0ed78d202faa6048c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c6b8f11b85800c9b6b1c7d74e9cd0a570f1a2149f38455da4e99fe5e4ead95ca970c3781f21ab50dba24c8b7d8aa4a1dad1221f8dd89f394d7411c2ab69c350163f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcde08ba415da82d5a84f2c427e39b03cbfa99485059fb048a7dca818aab48007bab991293889569681e825359bd36996fbe9d04bc6c4c07bb03e22d58ad356aecb87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28ec275c6db44223501235ba09213c1944cd01e571ae64cdeca666f520f3820019d73d561d9342d8c8002e670e3314a78511bec5f2f7fe6d47037054cb5d406e7f7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf45abcadb084b6b6a6daa787db3529b7f63a4f7848297beb0e20afbc81dbc419db35fd0a0395782c1c29056b1d2b98e1afcef25f829c56b2a232472be822509486d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f55ca70778a7a2913f9c7a88ca4f4f9d95054b391e27216204a9993b124c3917e1d32c1ff202a5892c7f2cbdeff556317d6db1ecd6855dde83e711eb2e4de4623425;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1057d83de46f6dc241a1d0e9919b3b77a53167f28f2375b4c36c04430db4ace65002a153d94af83e7f4d1b96d9e530ab4250753707e564207bf81d39eff9ca75a2218;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb376fc8cae101b960c77dfcb9dfbeff97cbe904add7e4e7a23698eb943a8c7e9e729e2c8bd7ad0cde6bca388e0e555f4079a78a5d33385a3a0453f32f5426da4a408;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b8e9dbbf168f16a0687c7736c2db1bb5360d8c7cacb725372e13d35d1c6bf3579a9caba5ea6e3c62e0d1ad02a1d23507dd9007f9fff9b9f77da3af22730e5f08950;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b8c55f4a272a9fd01462043cdcd5d6722eb1c2af437aeacb64006743809c3b7a47f2e515294f23f868207bad9b96b454dcdec6ccc08135635008475892d124d7a85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5585c8628fcd739a502b110eca36ea6f7740e21846dde6953e257174998f84c03c0424042734c67bc9eb3085d0f7ea6bafe03f997ea048f5b68b30fda34d4ba8554;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fcf28d3ece302b077434404702eeeb04398c81285c75b9635f788094bad152b482ec0b6c6e7a52751644fd7a61ed02b4e3d78aad2929feb1b15af8cd1d7e88e9700;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9242c5218d143d2c2e7bae8866c63596abd502d3d0c3bf81e8149f4ed9ec2a969dd28f818886cd7a3dd96b1b3a36ba3e95262138ca320cc4d91ce0bf3dcd271ada7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a800705c3e10e326d900140165c197a06efbce707727d0941f4f8bb34cd42d32b61027f20de20d1e0902632789bf1b6c065415fee25efcaf0b310818ffdb46cf7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171048ca2229716af3dd63f2a7c59aec8a337ae90595773d0e6be701b19d2e41d6dbfc48429cd00d0d5b18612c595a843a2fe9795a3631f7afeadeda89357a200d11a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1037689f0bc15ad0c23fff20fbf08cddff2050cac99b6f402c8f244bf38d47601a87e1da07d6eb5c0ad71d3390872cf5a6f3dabb419df394045599ee08000807a5573;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc47d9a006bbee0fca3097ae4c3f8b9b8a112562979b2f5b0ff82f3ef5783500c8e93b598d21f8cb53340e14659f27144161bf698c1e753beb49cfb12834ef496b879;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce5a59d93b41595a6c5e856e51d3b692e36f566f67822f7b9330e20c58300c30945c703cf3a53627c24a7b907682eb3081606feffbe726528154df74214c19a77d6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d886624675fcd97f174f6fe1777b1b4f40f5e1152a1c13947e9ecae6ef3f3a3e2a4fcde59f7d67365ae3b96586c846a3d3d10fd8cb27f351357eab146b1a5324eecc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1606e4563deb8bbfeefa990b725a970861b05f7a32eab9500b41174de7b4ec6fe244b086112ede737dff3937a4097dcd5c118bb2f3604b8100ac9a14ca617af2901e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164fd4557b13d67782f40417e916e8c1810061e453d7c9ac177abf20793c3e3570086bbdcef2c96a2285ddc5d9bf7eb87fcd6e2eb29c2e79f03aa9f314b7e6365a458;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142c94ee91d1751037b3b12390617f8512ff9bf64a3bea6c7246e74f9d77ae5fc382c445316af4343bbfd2875f5b885105e0355cba45e61927ab3e6b6b337d3c10042;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182e9b071bf22edc811baef60c39e8c8dd089dd44f31faffeaf3e84fbafa8577bc6957eb5455e806a6987e3bd62f0cc94022bcd1414d3703b460ff82f626257d48341;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dad42f9491df71e16e556253e17555b40cb587b7b7eda3c1df15611ab759e412a10cd7cb915b74aa539d95a65b78f397d1a6fc43c49d4c9f7fee867fa7ac68805861;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178c293209a676f9656091206d87a056d3f1822b9b6533055cc091c1fdbec9ab894a886d41e63f5073b86d42fae4acacd99383ebc85e34ecab13a2fe505f06adccfee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f03df949cddbe54015c3da81ec3973772d0ac9d7fe4f1b944ac0e78f747f2097b6a2a1092ddfc4ec4f93450e69ec3006bfd58d1e7b51b2831a94b83081e937a0c9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f332ef370a14bff59e5554a6f7165157bd1fbf3815fb0929881bab84a650c25f71a848a1ebe6c98ee75f72fd446ef9e8e22b3efcabaded8875e0e4328e86c4a811c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc26b563e53dcdb3e6143b575ce9b516d20694b3e04b4eee37105d442f3c8e933de2c050cb2f9305c0a11f967a3975ee7f63e29b5a2a7ff6e4509a208d6a090b544e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdc57f1d0ff1d280971ebde6fb8dc65fe02359199b5a51d33b015730d8d94e2941a52420a7d90d4dbea9d180729788d073aa325c5920d4ba8585fd09cde2843a9b17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10361f0653924761b9a2f0578c27a4f4152ea3c6f7cc561c5183ec51db5e8ca7bcfb4e7158d86592b3f1b621ae4487d0b852b5b46851eed62b93ca11b8a479871325d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdc6a3027c7b7db9aba80bfb6d5de84e402bc155b05ca610854d1bd68327b0cb9de59a6f416c3e57197191d85e2ba31b7c36b55ec98e5df1a5d6a14c58fa34c3e96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5301b5d8a9744aa5fc787698b52abe5ce18f02a90a676630d1da5f4676470aed5d6be56854750734548b44d932b9a8491b61a45cc38ada913f4c2c7f82fd4cf8eaaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f0fda8844032b8f507f1ee8ba4867e513564326601355cedb58b8de2a872011ae91649ec20dccb0719e173493ffaa8557010fe19e5b726cb3568c4d76fb9e3f85df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182f1ae509e58d85f80ded20870ab901544696cb63c129500e82e910b5021bd950987c85d8801d6025505256bcdfe9394016688619928eb44e65d9a1578ea35311cfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196e5f350b9e6706e447f159322e8b6db0fe2a0a62f5b8b4b42b48da538af2939f0271e0e6ccfe92578bd666ea92bb512fd00fbe02913ebc40f2180fe14acaa61a5fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21c2cfc3c7c42166edfc535b84514b42155c3682730fad9a9dd7f2310e7f6b4eb79d95be7ee4022922ad3d76619b66e1b68f4c33fb59cbf9b1eb763e06a564d933f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e175aa674a52261403e1e416437776ac72a6ad94b8d01e2d4016290ba7dd67f9b8b1723f44695da6033f34fa233eee1ad72b15d7a9680ee1119388df89fc5a12ee4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11170f7f6b3f645e7fe8a5487f478c9602514c2d30ec42d387072df0278f52e5f5e20a82ac111861f6a5d7908e321c32126f37b5217b9732afe9ecaca3e25161dc7b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had904018ceca241380979d9a5cbe1418f0df03281241b8439f78bf359e62026733b0aeda73d1a17639c3a86932f5b613f96ecf308bfc8a7dc39fea06a951977baf41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18026687c106249ecbb5487747e13991d5b3fe2f65a02dcaf16d441f289df86f7fc24009f7b86bf35465bfa4c37157e178cfe45c201d3c5d491c9ab59cc285cea4e77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2c76be58f9bd19f7896504f2d5bf1ca39e9026354c8d84ad63b3ef1af7b3d2a5301969d15df4d3cb26c0dd71ca87ee44a681ac4a30783f6adc7d2725daeb5e10342;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f91b6499b12174daa70042f3d87ce1fbab0d0929bf4cd1b5c52ced11ece1507804907131d7de564cba46694d7a90079e114a318b167c8f10b4966dd33b48b8916f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha22e3059b2830956346017c6f8c0e109f0c40291a826da4e24a4f01a4be3b14cf7fbb7e93301b0b8261f2ef749a9b12010d021116e4ced8220b710148f79d9b73354;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0e28996975f18ba2c553005a727db114a1e3fbe5bd248dbc081fdba52dd22905d83df304e37cbe6c17ad42d2b4a1e66bed0c48a992394d5420e6fe30997a2e6c301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb86ccd97964de9cb5a2bd14bf9772439e9ebf65c7d8f65b667d7859a7618e35ba0177dc55f3d11023de2b254678894a750975119c1dffd2fa125cc7f5a4f21f3a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d70d3fe9b8f2e241b312a4ad51f785d78bca8147d605d4801c3786ddbdac0c862b242e395b9cb5474c75d0effa2130c97a7dd32e0bbd9ab9892b1717bcbbea3590d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121775f862b39174d86b9a2c884311f1160061d4f6075b76b1fdf7c6b74e4e9df4844cd3c7a3d203e8dca73c6687a9067ad740ca6505d4ced191c8e367727078ea968;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h503f787e6526fe6d68a41f436fc4d766cfd82e3d8db0ee4f16864bcff1fc2ab543395929f99f906cdfd216aeb705051fa19a76570104505a7f57d0e8bd00fb64bd01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bedcfbc0841ac9f13aba3de65658fa4e2f0bd928ca0f81c38fb73e663d28b6de64690312686f9c11b68414632d30875e0552e358bfb0db88b9bf3faf35d8cb608660;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1695f19b4fa77821588363549e26db6cf204d7fd9cdd5627d182260b8911d47b62f661c8ff37e68288d8a563d4b111e6efeb8fbcc51fc7a84821f5402377f6a1f0b87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca9bd05ccdabf6a9590dc1e1dd3d84d5e767706231ca219ee6442df400880915fa67007913e80643ef0ca5c2743b61b3e9be5ce2fa63d9bd1f9799f768b5663bb026;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19df4f6bebc139ebfe16aef52ca5b8fe2b980e4d5ab14cdb5dd57c6a0d82bfe69d39f6b8406b4991b99048ab90c3f4ea8ae3a6744b038b42ed2761645ef896a475a03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5cb7204261bbf7a0d5b424d6097a6a67651a1d96ac6d762988fcece8feeec479d60ce08727cca66eea68fef19a2ade4cadca1be5108514eaa4dac4c214ef296620a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fdd4acc72038dc0fb365f2ce56f08500563021118be42a1c537bf3c199ce3fca0547173f45a13458de17fcb3bfe19be4a12485638d6023bc4381fa83fd3b155650c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169f9f473f903b1072df81976eac32a0240d2722cf91d4f34e442dcdce611b622509ae937f7c36440112df050bb86c6fe6c58435dc0b11481e87c8da36697a75eab05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c4b66d0f8e360ea4b61f5302862308acec8939edad83611634e1e2125546057b30bf9c13020b0c72a4d6551c013a820d8c9523f8c8023b8d87f34e736d7b8449a6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8631271ce4e6b5e97bc757f193abb43e2ba607a0c8ac121b5b8c3986ae69ccd9a585f2b6bf47a6ba8595c8a4e9f9eeb462f307f27c2197785ddbafee8be117a19a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7eb3a15b1feb532875b03afcbf58d99f08a41ed783628432e851f923199431ff902d4fed34610eb8829311bb40fa98741b7f450a82374b0b21cd42bb372635171f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf804f76f2dd17052701c01b594a2df704519b14d14e2e21860b1fcb529c1933838635065dd31f9d469cb1574b16fa5f25136cd584e9aa7147df024e169faad6e85c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3627b9a12f96a6c313484ca445648ff56f8c9132dddda1657795b6ac75925d752d2c00cb77c34a5ed2b32adfc5b538109b9a854c2ad686ee89b89162ae8fbe1cd3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3439589a0235919d8e7342bca63440c0f95e9a6b4ca9ab6d72dd27da0af223c55d3df28ab82a9166ca9a8318d6397e9f870cecf9850973a47be02265287fe0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a4f78862c4fa01bb523c38ad5ce669d249932b167f908fff296dc7c90a5cbe954c86d533f142e349a15004f950ba11153da28698c06d54af7afe8afbf933e8be767;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171626decb880ffc8f7c5a9d0126d2e4c41931b28f0be3c1756ef544ccb304874a4fdbe4c19976cba80bc90866e6070cf27255d5323e6c5742d33a543497a4fff1f00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86d2e09618017122c3783cb3837072856ad69ca2d9f196eaf8a97aa31198d8102e2a8b5137e70ba359221c464c6d6fda77659fb6c8818377821edf31ee93e8970fb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1fac44359c3c7618484930b98be18584fd7abd48ab9c695d33885f6d9450f80db714ddbe3150b3610977d401e0569e3c0340a1b70ea74bee2733e5bf8ead808e434;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff80f0d54bd6f979e07dc03e6ca9717fafe27ec827afc51df62f9b76377fafc3429f10153377f8d7df1145ecc7aee756d584a058353a0202c52f085fb99e1d5e3e67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139587f9bc22a508f0170690505d8b45080e38ba45e72c5c76f533dede7d7c02e1131c48e0e6ee817f27d0e57601aae5c4cb4bd05cdd0980ccb69dc13d1f4199b8c64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h784fe36bb0263bafd394d4c66e9bc788e5449a235557d0cc0fc45f424aacad9fa18bd2d6a8db194e8ae82b01e1d62a46a59542cd3558180e0ae89d2f2c72b2bfb203;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e05154d3d618ff08fd2c38e73eabc90f6a5926544ab1ec889d41250b4374b5f63f626b698ead4f892e59312431ebf78042bdd5c36fc919717ead638ba458f6d1cf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d683b534ff87f9cc6029cbb6e3fb5257030a5848c8caa7a40dc6bbe4addc46441f4a9dfe82d4ac28aef005e116f5526b8fbe601ee262c023a83c547630906d59d7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf8ec802cf7989d70e69e75554288d79275d87c304fbda2d4e9ccdeee1783805b8659dbb949ead6bbefd11c82b160e0744e3e0c7ebf72152d71a778a954b0c932a1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cc5d18d03917f62d6e8d6fe07603d3ff7ef052cac4771bb7866f34fc316aa10ca8e8b26470373bc5fe779288c0c52049540373e6dcba3a19b36c3810b6be28b9629;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ae002ce2afc39dfa0611036ee84f6624e1c757283a396106b936993bc8375353381a78eb25eb537488c76c27109d82d9cb5872f584c97e248a73a177b2b3097914d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f70512f3d6c1a54700047b6d7c254f047869d014ad19f3b264a88bdbf31e43db5d8e347d534db57401ee30df27c06aa0a8534c273a2ccc96c7cf52d04755c68bbe6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6734050c997e3b3a40ab176d11255e7839c2382fd4d2848ee184bfcc8ab8f44c9c1a14b7a39cb20491ab9335c1a1aeaa2bc1eeef9f5971f945c0d3588e32a572fcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h857f7bb2ce0a4fc174a3f724ae88e6a954f5dc1ef1a662fe7abadcf5421969e41563836980e34bb96cc8e6be77c26d2457261fd97a9f78b69eabd8f4abb234655ebb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ededac7e1218be45543c03fcbcf94719e889a367d8328b18162e7bc1430d19ae54830bfc6371b8b544b6c7a2bff6e1d94dd929566b8167f425965731514b52bfd2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107e27a55009a8202386071d37d3a70975444d53a11887ae8af000e4c51136f727ceda998fc5fa9c899aed8a136fc47da831baf2c2e2f8f804fb6138d41e1aed0a9c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83bca66a4ca8c156e40cf6ba23ed3f679c27bc4375ed000fd0fb07cd0ee85f0753d9c99eab7ebcd946cde298455d38940a1d5b562980208476cad1ce7997a7462b8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15df9f691388d59ab7b752699352cda0badd58816cd298e5f7c13ac9ac3eae722d9c2577865b3e62a449ac8c16e17c2b5e4e753ba4e0afc461bea96776c27be0b7c57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c95d405854906adf36eff9da9b1b6d395c7e6db903d5e6f4ad8cf0597275f945b8ef500b9b87142e66c8d7874fb39dbf4cc068af049b9a3aef190efd8ad7679aabe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efda96c87d5db75ba9e3175ae446cb3e10daf73c8861a86df2f998a115b4cec14d7ef5717f8d4475d2bd8c5366ca40717c38e3af2f00cb8ad11c7b376260737b2b0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133538db5f808ae45cc33579f763a8ca71e28cbfb74896ae0eebe58279bfa804104f9625dd7abaf53ec680d185c45d6456b7d04572c7c3b75e1c38667fcf3b720ac8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cd28467c6bcf818aff1c7e5ee31f3ad682b508d7211888424fb15c5dde1489d70de5c7b98997fe5c2f77f7b83daf5443dc1b0c6e79854de8453c3b9ea04c13e2f52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170f119f1f594fad9b8244afdbcfa5f50fa6c52c2e5f6dabe36f35ff73ac21a4bd94ff6873773b6e8d0417f1010a45cd5283d8b426e22e5834caa2e59124f2a64371d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaef0392472389da36cba4064fd5c3f34b3638a70036cea1bc193acb8fe4a713114b68b0acdcce28601d45cdd278267e294725c4c77a22d655a0f0f81c64d31203a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eaf7ef775cf1a25ba5d1d6813f7ce07451a9a58092a4e6cf2fc1cc7102599f24f386f02de17e4f3dd0eaade8f9317427c06ca8311d683518342368dcbad11e26743;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62424cab30160ec74c7d6f63202f6148d3bedd4370425fa40262b508385510e674c9f9aaa979a39fbdf311f4d615df7714e814aada534b4c31eeb6f0922090b8120d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1541f05e390128a064c4a9d84dd6359c0e0cf2824fdf918e58ad1b7ed65241f087955745929f7ddcdcbd2e8d4401df185d68aba6f040cdb2aa7df94da900f38fada14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1debb5976bac87b4f9f7d54da52135c0bafb9231967bcb87fe5135dc5ba6cc553980d69e94dad5c60581fa1835495b596e3ab807566dce276d75346b58cc10da3f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a91f52436708ac568ff131e57f65e9a7c4d5060587f5e7d07c58683d8b7a1d6f3c8edbc6afa3f88d375903c0e810b52a3471f0a00a6c6e0829b520e8b5006ed17ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf27edc75e11058dea2cdb8627d668d3ff3756e211bb9cef72e5de82cb628973e0912c2258811adfbaf5a7484e7d7a87656b4c18cafeb9a03345513c2a8044b0d1ddd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1701b6990ee60dfb5fb1f9af43b292762dd47ebabaa63d44ec9f619dc811df1cddbc899f5a31bc7ed8f1ab2d08536a123b8f3fab071604f3b7321e754c4befc7b6968;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1defa468c7f9eb240543bd6ab5b2db9d53e9f36f3cd5b76b6a19a18a013224b3850949fec2c07fa0052c119bf6df185b019db5a011c2a41025b324dfdd9e5ef57d306;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf81aa2825ece9842ca8b4fb959892082d23322a4c2efdc1cb78118816915d7594f0d373854ecbaee8a0d9e08e7d88df41bfcac5859f2f1edc6863c4850c0a4a30d67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd4a92ff7662197316d7bfa48fe11a954085db929738300c223f7339c6f5c58928640ebd8c4caac680539105ba93e5580be00badb1e598006f7f241239b0a659ca29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a7a04762e606da82287b4061b49e74bee127dfc17159e65ec433328c38ac4af6a2ae6a578d1f4ed1edcf193c8e38d791b18deba43421bfd561093ddee7427c239ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9f7042e4e888d7ef25e083d0276fa9c898509f75febd2c6ec44342c8841d707be17c5fb630582a4714412c8962d5b5bfd3c9aee445752bd48bbc9ec625705b27314;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1930237653cb90edc89fbd69eb2a2f8e8664bb79bb20375a54ab0875ddaa569c33a62789c3a31ed963b37526d78f7a831034b2752e94b7b26cf68f0e8cd5c78f849d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h907018362138ef8ccf6bf095e2fffce07e4695e99d83de5327f75db424df056cb6240095373c65099562cb888e46659f1fd854b7c7ad71e2f75098f8b87771acd412;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ede29600db519277fde048fa66b2041d39ba0ddbd6c6a83619f114e9e67ee1c86318ea0d12fb6cb5e645d815d04642270740e9cc3cda3d023442313024d83f1007dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a763e79f8d1977a84afa8df0bb751efcbf3ed50927317637ec7ab6482c48f5d3d409d095dbfc513c842a52cc2a9aef2f6b987820d77e6c91440b7b9ba9d0d57e26c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebf69b7da0329ba984c13725d1eeae8d7b9b54247d580e00de9a060e43df72340fd79fa69cc56cd7b56772e84e3f6ac1c75b261983f8c1197d485852b94d7a2487b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h542bd22204001dc20637c63dbad9b0e4ca68890adc3a6d150c9c2b6c1787671a5981e115694838003b6ebd84201564d7d4ecc9db169ad674aee96ebd4a6ca5758e30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d48f90d6fb2b04d4b3abf3ef866e3e39de3865e3c3adfb2a1c0ab57e8c6bb606238e21b39077265d110d772ddc60a301bc290e1d5c26e08511d2d40785de4063a03d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0228fa59060d998dabfd79cea09ff4be865d21c176e57cc0a792b8a5231fb600c20fdb18bb264480d2aff4c2eb7dba4595855cbdf5ca16be791e43bd34ef2facf50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1200b596db9cb84e05a7c2b60898aec3e55a86abdfb566c31347eef9d8ba2cb3e36d37438b6fbcd1df004667935f6dfeffd454eba80a8eb582404a7717b13792899f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149aec6cf2e2d93336c5ab1b678cb254d1bbca08628fafd1df96196618a88e00fe86bc632cf4794e792ad3998a9f51e6129deeefdd4f499ff9d07a1b45e3855fb8657;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fe8cbc42247e7f37f21be1a2a12aa1adfa85c11a9546234b835f1015f6dc9732a4ffef32e7069dae5e9899ab274cbb2863814316673d32d443fa0a3ea957bb944d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4997bc5443c10778a6e07f825c47ce2a8601074eba62fb55d7a139a6826356ffb87cd1b42b935854a65d9bb831e287e307c05b8417211e209257c5bba590897ae5cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24a6cb9a21f01125ba41485cdd9ae969c71d4e545d884500b62f21a30374bafc6831e55942c1adb41edac39c7c258fac93eda000114f2123e1b064732f6f0a9b6626;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6a55b28c6c808534c7c229e2ff13a836a1c26d0135cabec1a53078e5fe4a305ad9cad5001b1e5f7cf38589c2feb1fd318257eb8ff024a5d8bfa812a97b472c42cc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14768294e060f82b0cf7b49618f422972f20b892fa18a55b63033323517277677ae35cb5546e3193acacbceebec84abb420029bedbf2961ed6660bdfa6f5f4aa62d8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86541797437fe2439ad17ab56bd8085be6fe245eb09029dc165b07c7db5fd53ba69337c669c5d08b0cc923e596704462d7e8259911bbbc80212895f5ffbb31fe3a47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2354b40acead4909424e712c3568004583768b64b77cec5923e3624fb0fa21db405b3297c83c04a41765e050455ef11f9fa5c00877cdefb19139062250a4973a627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c11962982757609a844dd338af0e4fdd224ecef4b80e3251e9cdeee4f9d7c9ea85b05a5fc679a71b8a63ea46a80180c6285d4d56ff7ff0e74c45dcff8e2565b942a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4b6717e8c5596fa880f7c5de0d707893f8ab6a74c0be91ef5dca3c5336fdb7a97941b82f1d499e0511f6ccd34f4fe605cf548e31ee002d2308d30445488301bb436;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137800dffe53d3c7dc664ffb1bec39674885fe745ffbe81d64e0338353fb703d159dd9a18ab2f9e195ec6a95944dc571666ecd146fa49a8924ef262f08702bd45992;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd671edf5f4d1caa866be2d9e531a351124bedaf015aa7d35b3a919d916971d15e65eae604fd63eee6a21f591f1a9ab25bca32c6f143dc3d1a7ec2435d3aa44cdb64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190fc01599e9dc1dc8ad23d4892f11ef651e857008843a1d52ad935b40049a0cd721d279424a8fa13cd8d0ec7c9f6aedc3aa6b78c4dcb5a8edfad739c9128d5c26da6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187b675b478b3b0c9bb5522c3662bbde081b6167a093f2b4ee43da792323544c302fbd53f9412398979b5e667368e713b03bb9f8909021667e6451493e3be77252187;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1747d3f164f7605e9900e1f6165df204a8fd37faed9eeb6c2dd14c18d92a9d73b74eb7a3fa690ce07dbfa403699f826a143fb1a8c1bf0861ca9f73558e6ea6308a81d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f4f017805820bdced977482f27ccd4890acc29458faa838d29deff56e40853d46d496360dcf950900e21091461ac6a970d40f0296ee364caa2c9ceb9ed3083b90fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd28a28956c00e497d74200ff463ffa2d09d6fbbb4f3cc03ea21069eac5b1feb9bfedeb053728f140745a94a0ea4d9357f4e7cbd72ed173f0aad4e4c74d0d5bb2434d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c479a505623ce55abb79936c1ac1a37fd8cb3e79f5986359ba5fac8517ee556fb1598c716ef1b83f5a5ada85b38f6e27709207d75acf80a0d3774224fb1682452db4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h913f3e76e22ad16996be8cbc8f4f67cf4a464e16379bb0f0cd622d62b7740e00ea8e790ec8f0740a64a546ebb23247ad9ad2d8e2347e50026fee38d5cfe01d5cc1a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7148845a2e9a46e428601af832482e70b40f5f3aba1349bfce188b7bb73d9a63df5fd044c3727ade4109ae7a9bfaca791356397ebd661c28cbb241734a0fc335139c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf077d915517fee7a4b56505d37235d2824bc23d1e16ad81205f16319bef0fc63d76ef0e80c95f4bdd00ec44ed4fe323f5282c69abff432d95b24c00b8dd225f7a180;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f968acf81468edb950f49fb8816e523fa28c47bfb2eaf5721c31e104da3d0b981ef80e475fc14040dc51c370e8ccf659f0ac72f7859bc01d440337ede8dc768766f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3b906f317575b557f1c45ddddfb2f00716b31c0af7b0459064ec3d4b44b76ebaa431c71c5730fbe287ef9194998f55a199165704e1983cc982c8fe44f0a4abf5c79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c28be36405bc84dd111c36f2da3b2269a5b88d784f954e53856405d0fe987883845de8e019e9568cebaf42a5e35e4b98df80d724da8c74bdb2a2b43c8ff19c8e0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12aa3972a75edb0ebb3ecffe96de2b2a5fa9396b610a62f06092bac16e075c0527332ac68a8b5b9dd84adb0d4cced7865af8aaaeba57b0490995aef13ab939b152c8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1650fcbad3688367301c00b876fb7fa9f859b40500f02e669c08f0cdf53184ad7aed0f3fa6e44f0fa33b5016134f1ba16d467c71dcb60bb9dc37c449b4ad3ef2b048e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h934c1ca3f2190c58ca34c95e313e62426495d705c6bc210c24f4fa330d378a1b6eed32a6a11d6c3e5c3d516754a8b35b7aa7f793dd4005df25d06bae21844ee1a808;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed878848d5d4a280275f2c4da0b23d905dfde52d80a2fa4655910ec6e20c7db132b475b3558c9290cd811eabcbbd7993f4c5fdd68c0f99ac16a5cf268a2f0e2e7669;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb2c2dd8bb5206c621660ffa4cb2690e663a175292e0b313fd9cbe54b745b19f008d75098a83d8ae0850129e9eb6601200f305e29a31cd3adefce9abdc078f3f55e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1848c6eb6ea472d94123b3840c04d1daaad36dca81039ab229962e588016d10962f25ad3f88af5c359ab7dcf7f5b1b5e1d490a4084f3e03d89e96287fde40c4faa32b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a2fddfd380a56e7f88bd4a48609fb273bff23fa2b1397501e32ff1168b68a1caca898f36bd7d55e63ee074984188c5dfa2bc08cfe4e2d32c56cb8cacfeb83013af8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1743e14ac8de5935b622e37a1f02296116af3e967ed1ed9689c068e323ae4fcac9296172ee124c995aa1a566cf5afc7fb04205d28d0e9c6d4c2dcfc1c3224e7dbac07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5219a726ae8c83bf67b736b67da84afbec38f21a101e22666d9ea57ae3ce694d9597ed31b8bba2c4ef347d6a8ed59e683d034b1a4f78576ec08bd119dbcd13c8acea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5f588d16b0026491547d987a3ce68c4f10afcd8462ca0a05911754f1bc5b6e3f8945d95ac838cff0ee19fb724ee4f4774489b7ce1ce03ef8de4461140556d2061dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcba3289cd7bbada698440b75451543d18fdb932500cfbae380020d504b4efb81c4510dd3b25268fc2b04f9846d7264631c384d019ea549e0297e5d23b109fa639f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1318381f1bf5feb61b942c8bf210027bc351054d0d5cba47e1cf37ea9b1b5dad3f94ff471ac0cecf6bfff105ce95e83dbaaa7c12e920351517f90d4597f991017c70e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2936e3109289ac74a6259707a37c7da1cd65db9866956a715cc29efbc54a297c848cff334ed64733cd1d69fdf87e44abe4869a20c8644385b496c1d48f6e796f3ec2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195516201d02df679d1f72ed0368bfdbe055316ca8320eba63c54a2db3f8be220305432cca67c82342dbb2cce51c0cc376b80d497280d7388e7373c2d812cd5129983;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ebe33ebb6cf2bf834c03061fa405b5c57e62de56c801583b889e64f5fd2be908d9816a2c7778c10b7e48aa568fcf7e57caba291634598e3e8e4d5e196612f0b40e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h730d4a5463bf0981dee6caf8583a151a3ef3cce53cbe950ba7e5cb140b034f629c9e5b636d14993d72d3fd16d6ccea3ce8edbfc10fba185b609a9130b37274b280df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18526d5678c49e1ac09febacfd34c435021f998f8462dc18e909b916a732723aeaffc7813ebd4ff55b38a01a92f864579ed16aaeab56b6360c610746b3aab399020fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113532d60fee4704ae11100729d9cd74fa9ae9407c64ef70f2186cfd9e78c76d1b4aebebfd3e74f1f6adfce6d4bb93d1cf31cdc9f5ccef11cb0103d4da99abbd0952f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b910743c3706173cae6b0cebb1b6b90b715361e8644069bc7b6ee3aa625afa0f61b87ab4e921bf1d9f065713d8a44881cb086ab974c0dcd8e5ef552bbfe29def77e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb9ed4bdaabe964794bd0f0b683c2461bfd145b9318970540a6e234078c58e78d7ae42bc66db16da08a0d35e3a4cf615b30f18887303c5ae793474d4b6027823c27e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e5c8f1cf56ec5a6953e98295c3207693b17dce89d42d99b686115b70a94dfd6eb60d242b23e28ec58d38ed4c4b4396d28d4500481d564ec56a94257cd8ab4f95904;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec8074f12e464fda9bfcf93f12f04a08b7ca7c345a0875fe6a8bb2a950db551c4cdac6d5923704189578b33e44943221d72322bb4434e0273d0504cb68e06c895aaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f368469dc8f7ccc41b9a7ddc8c087bc6cc2301ae53622697a5a582a9a480c5f78ec43087a0039f1be2d2212747696e28233bdfc2168bf0ecfffc4e090903fe9a67c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ea2ae53e19153649c921320ca234de478abc4c3cf5aee921b878ea6cf4af4511d67c5cbe68b5c0b9c32dd5e74c76bb7bd8c33a0135d4b3fcad0c532684dbd7ed15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c510a8fe0c21186637363589b12da40f83bae464908051328cb663dc478b91c632766d501ee98e45128cd40540dcf725bce563697a038481ec65d3609dd7974ff273;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef9aec682031d766532e9aa5e3bf0c198a3a8e96749183cf03ccf3c642898b18cc8b5822a7b7c9b2a607f81214d0100b1131ae246ca8dead6bdfd9efba93c0d3907e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e0b500b22884563ab1e18944ae331d9ef64ddda78a8884805933744134bff619ec691550ff4c0804ffb84f4a6bf6838180efeda2d18e4797d5927d3ee94b0ba46ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13efdb614da5ecde41b63129d0c8ba4b70a4556809ff6a5803efa17d5b59bf8b386e8228cc5788994a909e9972d8a7a775eb0c258a8ee7d2cca16aecb085455228277;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1cfbb52b788e74a03d2336aaf29277462ac098501793301159b2fe7a38aea6787e16de5da0e9effb1c6e22054b41538a1e4409d21345d8a4c4220e58f02119baad0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf45fd3ebb721d2331354894a4fe0f5e3bd89b8ddadec6c00380d66ab41831bf987c3adf0c3676a11201bb0ca2ed67206730c4b9bf5ae111a4b5ee1b2eacc3ae1e97d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136f1664c07b7b3552019f23fe83324fa42d792e4d48d9a644052852c8959f8daf0550e8213a3cca89c2eea2174113965e91902ff6408a75e9af7d17cdf1233f092f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h262bcd7d2ff713ff851ee60f74788c8a5d427ec36b60c824e99621d28b0551aba4206e7e67d132bf6abcc7a5d86c8d3f9dead5c06af8e9c5b58acd404709e208daf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f32f8ddf40d017c8a9de4af82c3a386d54d65fabecf2f955da7cbd9dab0056fbcf231cf674c6d6c6e5352de686532f68f1cf24fa6fb4fc3ba33edd64c2055c4e16d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d224912813f1cbc680f7e4d8199f25c734f2b06792a9407f9469471cc23d070f22ebef46668e21bf6676ef2105eb6ca3657c9802cf5cb17368df28a05faca246850f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c753b06639173623036c39ed19ef050398c2a2e835768601f9dbe5d9636644b68c68f853e8be7b844710a6ada4d6101b8fc3ac401ce7de2967dab9a69230e7ca861;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18327818f6d1e98bc810e2cd2d4a129dca6d092a9efab0b10c07e8e9acc702df0ca25c2abf63601d59efa2b6c412647e1667c4d3d6df01374ce1281453b8404fc2364;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1501f34503d1cadcd740b51e92b6039877e401ea2b3e7ba501fac27b06ead77b81be2c3c02177bd0b6ded781b571cb9d1c3240b4470602c9f98e22d0946d46c3d86ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca441dab88d082ab429da98ae58c42568b4eb43ba7b71e4b114dd0560889f27401c467d509f9a1974637cbf85024ef137097e1f6da01ad1a756020f38ee50a703cfe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195686b1ae0bcba31b58c9ff9a027a11726335e8527125cacc5d655f90701302274dd3dd549b2075f3c439308c31433040e29e4ff40454e929385d7fa3f3d4ea5a40b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h475b8665008486057be902a3a90eb5386a8e86d83f744b4d508c122123981f7dc0a6da6c1daa326012b0b037e43e2943386f2bf2f4e79a71a74b6748636b909abc1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1868ad26255485b70db100aacfe76c230a58aeef9c4bc7656f04aea0512b985fb8fffdc29aee1181cda055676046693100ff66138a1d1b041a045a0262ca0a9f184d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f236424086d0bbe5412210f85a4be94184f0b18059e8afbc7bcea271013c59104b07617a7e6d550949f5af8b8820a9ab861dd85cf1d7b958fce0a9465de5ac54cce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h929b1cdcdbf1b77d721fcb759232da2f83392072560dfcb71c60d8412b9829cc8e535601d564d5a0b07935b0d02ef8594f8c62299e1a394dc646b97f7ad9be0b7653;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed369c8bf463e2b78b835fa82ec97b1269f777809ddf98dee3e04cf073453dd3d7a0ffc98621f7b958c3db6fa2f8ea2c47568d488e7a58478cf992098adf7c6c2f55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9aa7086c52c1a954370f430682f61b4f9732cfa6c89cdf91bbbd415cbe00266b6b0f468475992e9f676d8624e5b36f6d39339767981b25b3267c75efd8dd7681e5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e720737b0c9d43d7593ad244a863b71a9a6b00368f5208856f46041dabf92c30da645d84fbd23bf69871c40b96a39ef339e93411a6fafcbdfd92996c5f3630361717;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cf07caaa2c9c5a760bc5e1de199a751bb1d041a1c0b06fa2497dfa961bd732e8c6765204bd4ba76508ba82982c80088359c27b77f24c648131e84d15d8be1457b17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a2b00228bff178608c41ead288516da4dad0588677287515f55334dc0e94adf746a9209342ff6cab9afa8bc94e587226e3317e93240b52415f85c18f085e424f019;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104633ec49d6a3052a634102516132ec77b32253ef2683be9df8ea960b879ac8649c3f0e7800602877ceb7cc94eabd2108acbb2d753a95ea3b7ce913a6bee4b5c7e5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df5443eaa3093289a7a455a3f82c41de3145720d2d692a1318f264e572e3c4353249054333e16d55a8e8fd6f9f07350f50b124718e819eb5b64817e2dc15e391f25f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6022e7b68bc5f8e55ba266d2b75141d6e46bc56d70c240618af1fddf95e5dcc2ed619242ecbbd053dc19de829fa4790fe531e3b33065b1bd17729178f3644f95e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1478d668929a60a3f651a985e1cc1b845a1cc78b3a77888823772d68a254f6ac18e8abd88bb6476805af3746f0b94a2a32bbf5abac7d51ba8423f159c046dd0a08a94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f931fc58d7f51a351f0630bce7f29183aba30690e9f44a7211a4a75ea84e6361fbdc59beaf6e9934d007fc06d2e47d70f38064417ee924b111a388488be9cf12e74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15cd8e2b32b37c22944b00b23fb68d16c0700c7f716f74ba3b6ee38bb4103e91f9f8abb451828f50eed5ae9dacc0d34380b4ce7388db873207c426eee84642423bbc8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176ec244fed3e5075ddf623dce8d14dbee7d032424f6ca9c1fcf692752716043a8b523003b9309b55acb392e76b5c31f5e8613f1ac9a963d3b7f65c084126d73c290e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e9bef24d66cad1f6ec9ba9ba26beaaa40ef93de22a17998a396f2de5b2f5b096d1cdcdfa44e615ed8dce02d7c3eeac2697a2aab11f1e25e54dc2cd7bd466b4d1fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136b752be2426c88fb090db2112553564b258484a0862ba9ae4a3499fb685455a5fa932cc699917f136e512dca77b2adc95ece4ccd176b6bff41a5192d7b9539b5bf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3b2622bf7822f9b2be0a98a3fc642c10db4f4edc8927c320dbbec4f15a62ee8a9128739d9e0e64efdddaa3261c4f92421947d85b9ff598ebc719089d975f317c610;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcfbefc02c1ac47aa3815de4de60f8651870f4a44bf5354ac45b8ad38a9f7603efaabececb36b95e970676779129c217e2b18163c6185af309f9dcfcc56d0af32565;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9e5ae5c9f94ffab752268abf9ade900dcf3463c811601149537a1fd15cd876ca4ded3a300fced701e7b413a264410fb9096caa99ac9009e29373a07604b4bfd5925;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ffddf6934f494108ee206adc7ed91a4009f89448f6ae3373bab7751634390c5cb9d3cb2d191f2274b492cd7951c1ab898aff6c7b89e0be779e1579d47048b74897;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132b1286d282f2e2f9237afdbf6c26b4b45190426c8abf145b1bddf108d51fc7c03eee365077cb1de5fc9e25d51e903468b89947b718ba31b965b3a50c8844b6ef769;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha546cf0783bb66ae3f7bf2744083ef88798aa3cf903afe7298f3ebf7a4196abf85a0236036ba19b024c91a1b519e6047aaee54407fb57f5af7d96ff701bb037fbfa4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a55bf6cf759182feccf917ba6ef8481fa4e4542affc929c4859131ffe648c43c0b0a50079d078acd5a7605c8bff891a1dd380442b9b15331d2a00f963a2e543fd573;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf3d62aadfa29c5c7d42028d0838e87c13f175350dbdae742cc78a83c926f884d6cea83b4f44c45c23c162f3052387fc4bd5bf1d3cba34016bf08728e466a49804e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119a7016ed2af08cda10ab2ebe36e79af55f64a56d25a0241b61042f27f4a23c1a0e56fabf1fa485b116ac0daee2bd9c1eee915237f2832c4f51ca066a1a0ebce2669;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha30bf547bacc46f9028edded41de59767e503ce0931bc018c2b61523837369711dacf5c7efea57faa51e4b956a09ff691b62bb4b16e6995dafa35faebff1b59f55cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db9e99c23f0984b28e38e2007766499acace43dbc1926a1fb8fa7da164730bf8d644cb7ca29a6dc25cc739b6d76ba5a5bb41b414d5926fcff1db551d001c25f9427e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1ce693ebd3e44fd73d6094eebaa7ba1daa30de47bda67ed93cc9071e1a343247ea6db534c0ae7be552665379f024cbed86688aa22c1b35ea203b50dd1254babd9ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1779698fd22265270097e8d921c1c21350a48c8cca2cff5dca13d52174751be8526d9bb49bd31cf53a6ddb396a06270c0094a63eb0a87438f5c9f80cc410a70372f6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8722e97152b033d663c3d13e9a5802b446a5ad5c7efd00296fd873633f09313637ca5c5d35a2d96cf2d4e81d2ec8703ed09b91e429ac055a79f82319fb2243b0599a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bdc7ad9e5d529118f073a8cf9e63405be3f5cc2c48b7fb25cd505f22ed9684058cf00c1f544eefa9d0a794d4fd8f3a18a6791a4a9f164c014a659d109ee661e91f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108230fe15d0cc9e75b58ae42f6aa20d54b4cf29d90e48acb202f892f4fb0998022e63f6deaf0f893de971d7b98965fc879e1bd8f34cdc3513dd3fe17cd929f9b0b40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c5badfd43c5fc09ac03c513648d317251c403a0e5c71d4de87f403ad9179a2ddf262505fa041ed7bc8208489666a257ce98147a1b2b237a61639c35c6c8b8b850bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ee50f2f2b29e5ba4e8c847179f8ab25bee013671ce68b2a4c288ade7a474ee2138c22c3a5e7018ddf7f574ba76af4faf7c428646bdb200ec443a88ba0ff11674c38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba4cb8bf7d475961ace46fd77400100461f2b6850f0c43ab10b61624de34e03e0aee1305547da1a994f211cdb5212c328c0ac7818704c80849f8202322704c18add1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c39aae1d34c214b27edde42d24cca7e28ba80ecede90d89447a21449143453a14c0f205107664686e024ece7bb1202ae81d224da906710e386d45b789346cde8990;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4772b76444789be605aa6af620fb2ad5f86b817e75acd22d82a56141ffcb00cade67671ebab2e28d2636e578b8c60571e4af538b74a34eb259a28aa34ec0d017a1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ac37919afdd455b01f9d7d34fe44c5519c7e9274e6eca6ed957ca2184ac3ef407914320dfcd89e3a2c32c7c36a186f33697ef23d42a9ed8848b56e188b87ffea3f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd605e60de9315fde21997137e3eabc9be1fbec631a47cd0afcff3d95d99b22eb4e8e4937b30234f5bec202c0c84b58947c4306b838f5fcc1bd42b4d757e56e30617;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80624a3f924f31093580a88d41b1e11b5bb1e7be807d6851557a70f3dd248fb822e833758a4822adc1cb3609c0f01b75efa42fb052326b969049af49b15bf9048db9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73aff77ecb869b42cc96b50f0155aa18e3065a72c49724b0b8da0dec181ab5684547c0151723bda3eb5f1a3c3ee0d97d223ff089a7a59abfde7d3dcdfb7e15cbec7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1576b2829c01bc621792ae298675d442a1fd38bb68de6bbc3ce6347d98536851dac44f88645182d2f6b052720040588c60c1d1b2dfb4918fa62fc16b6752fa2e5abd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdeccde6d2c14411fadb07da069d1c718748c2089ee0f70c4ae2fa98e26de167160ed0ac5f777d3424866d26dd0a5bff6587d8f1af187bbade7b9127ccca29947890d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7d26506fd25cdef50eb302c8477ad5b0e74c72bb3b04cdd274f0a7b8c86e66e2ca958a0fc3adda44f22397010a823b66c000e41629ef203d963f25f480b6ae6cbf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1037f6e30c94c30c0b1926181eb50e877a3758189485a2c5eb266b4eb748748d6a2d5ed51f8c05dd2278180655fce882e648407b1147face6b10e50380ba0fac3ba3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a291ed0eefbf52050d32d8d21782d4cfcea9e437703ce7459a37a9d551402ba0f91046d7a47b60d5cdbd5e419307a8c9c7402d00cb7fba55eeeb4077be08bc533078;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16cf4d2c57d6a4fff3c5bceb741167be7815f3786ae293257b4860e9858dc9e0714a22cac39e8c70db7d58f79c84fa85e7a8f654830cf593dae2059393c2110c87381;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99435f2d6efd26e6cd7a02b5f41e4ed59a48d19d2f1200ddb86d90355397b5cdc881b9732f3cd13b019da03d972333e2ea030ad7c13f73aa5c53228b20aea7ae575f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d0c9ff4c3c67572ec55e6b8e365a0467b0cd12337dc55aa964d7ae49d614b76e82c287aa3ee9edd35c93ddc09955bcd1a50527c47b45441d5771527991903a96ef2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0a00ef254bc9e6eb588fb62c2e76caf256c7527e3b33865c2c84500465bd83178fdf974fb12925c9e7f4d0e6427fa70c49097afd1295332892042ed12c6da480f5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97c5487452812468d8b8a1122e604257e2d85e2d4808d01c6b71bbb5cf9e954863a8f6e6c048d7c668bb707a3aadfbbab2e8f7e4ff37b21f2ed704ad15302b594a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c082dd3ff0e667b5a844698ed23a2d907be4fb76c01298bd386da89ca6e6cd937f25b04372915963319b18d834551adaa85f8e39f0b5d05c438a6ca9a4960bbe0282;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3946bfd440f4a4e9cbc3274abf42fa03e5350bbdfaca698b76125e52c0374a9ffe1fd6fa1da14676e736aa5eed921576dd72135ae2059d5a211c5b3b2d6282e4472e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20a66286b6524556956dccecfefb82c584db0801309123e62e1c7b9dbc8e9b412a16ad49520af077f8484acadd59fcec2aea9e6f53119d2138c18b6fad60d23f552;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h157e40bdd6b7b94195eb5e7e63a786f1fe39cb5b0de3c95df80c9de2353010ae0d7ed93ad2ac9bf5566fe0cb9813d81f543b3414286244fe7c3e5f4dd87a37819b614;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17391757e87826020d8e258e3c13801277d827647ab679a68789ed11697b7bbf0eaf3647be880723ddb42e17cebd3edd1540614f6d1fb527e3808db11ed2b2a0bd060;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf19bdf37b279879d3780c5255308da14e0a671e42ed3d7e7c5dd2c20aedb6b715ea11b1148b09548e9a00020613339eea9f8700bfb64050de8c3ad760e2e4d0d86c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h979dfc029e5f38ca3acad66929f880b25405416cf57e3b422d1cb74615c8cb1a276978890e05d3535594ad9feb6ef3171668be9ad20bed788c795ea43dcf08e861d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b30aa1756480b23f1b28d6d4140966a502bcd0f57368a5c149109a02b97658ac9b8765fcf4965bfce1dc70e56a6c7fa20745fb80779074bbb6924ebdeed03f8d319;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12aa5b609f6bde8bc3687bcb55c3917ac8152946e929d279d95b159f162886c77dac929d293f4a0d8be412501b54efd49edb58573d9ed31228bab491f3a67bad2e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112d4e2133c298a9bf4bd23c97efb03739d432588626f57521fc5a13abbf9b8363dd4fdc14eb626d8a38934f69080b8ffa1de1f782c010e1a3dc09228aa15deb288bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16740a989f2a4e3d19d7d7850025542ce5678f6df429fc696b154dad61f888e94b6506c323f40b70751d7d224cdbb5af32c97261f39c96e02eec9436c65927e51720f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7a7824c34ba4e550d1f54cf0a0042f35d42b84233ebe5da27130982347a9c5be916d40d936653437959d9e820d58c8c822d2ae9f34aa5d77ddef969fefc6d5492a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1976aa4b9fd96fd70b1bf222542e768a7d2be255e6f9ff1efa156854121e0e917a179766141beb822e300f88bf20f4a20ace5fc81ec72d959c7f0cc756977f9596ef7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd80ab49a14fe1c036d74d6f53e9c3a2915fa52f01ad4564b70aaa28f3880888248a20d9c8d4396d6b9f919e7c8031c94171d19aa93e6ba77cebe9402e0e71a7a9d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa4727bd393e274350318945d1e7161c1046710ffc006a355852cccef3ec1dcaae348d04b69f2ca193aa397319b278869114e918a3e40af7277c002c2528294cc5d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72f11d8af2f2f3000c76926a1b32ff79dcca2139982f0fddfed221febd9983b7150b6cfc570db2e051d0a82c0da179488478b2ce5e2ec4a6789ccec1851075642d79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128a0b4e1d799053110182d93601311303b7309f98a8a207d260d5e56ea33036de79b3d2142079b356125fc012960ccf0a75edf217665c24efdb599edfe51e1704d41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c88adc5c466fff9ed99ea1a461c2142283f2b498a8112948b4c19232c1d07fb24feab46128ddd547497ca521d6320dd5694112e51eb59d957239c6a8a4f862be5f6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3fa8f2b0679bb09af9699b21145c97049d9cd81f655131401a2d35b1d8f98c60df57cb13bdc01b66de9bafae3b99cf4da5244ee5061425951824ff131c1c8abc71d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3de73c49ed7fc0092c63b6a1f98de4a34bce0f17cd8dd22d9adbf3b4883affb75cf33a1d0e647f9794ae10abfec4a1ef162af552a7d46ad9468d02a3aac3029bdd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1469445ac389b192f15f9231d92d49dc594409d7c1fd22168e5ead31c04f5a9cc5c75ff2c29762b9c7ca0069f0dd1a765a9862c82fb2535b9161422e20f3663eab0a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd117b7fb97ba98b43c540c087338dd7bba19a7f3f78b10a7455df51965ed5f8df137734d3761d0e44de7c30af81adbddb821612b3eca040b6e01de6318a7eb4ad650;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa33abc5fbe2e934af2f835151b357bdb0241d6494138ad73fcfdcb7285d535fc135dc7447dbd1d60da6b80f4a38a93122c624660c43e14f66c3b64533348c85f2b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198f046b666b62363d438234d7b41dfe4d4dfa66f872dc920154741be549355f7f08e05087f3d5229b0489e64e452bbd749a92844aa98a3d48646d221dd3608934174;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34a01eb461c0d4294edad035bb3a0bfddda58d230270d8ed0d163acdf820fa628acde275506a3bfb75f99b4d24ba7afc8061c0569fb50a8d8d6bddcecab718565c4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48b9be568051d1d2c8c825dd6f8de9f7f633ffa821aac467201b26228aa9bd5292e2091373aa5428d10abf0b6bacb8857cf1ec281204ad647df4eebe4bc78ec90cb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1a6fc5608c9968d6c019879465fda86f71259f2e587cb7bddcb1cb2e7e4c3d5938b93009af4a473b0da8543de5b147a7c9be2fcff306b6de8aa8094b64798a87004;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5b7cf04587ae156abcbc5341c8b5949ad338eaefb103b6e2ba7722733777f0a5ad7128eb494c166e74d1919376a5d1abfece30808ce619dcbefd0ee401fb277ff6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175bc7fb9b989d9d6df4655446b10793b1947a7e5370f75c2e7b1d53134b6c9601700185d3fc794ba0e0372b0fe499a767c9d401cabcbad24dc67f0cd2f76de18303a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h893adab241996ee6c3d0931f859c83e9724b7d3d9e0e9651d898870dd4bffc9e47cbc233b8986fc30d7a91dcf971f4626689f063a5aeded9e1604ac01423bcdf5b31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e4b3966352cea8d4219b330e4e2b3f6521814b6f72e10ca607ce17fab615afb0249c7047200f005565651390a3d19ba991b1af079c620dcd44cbe6428930ced6f8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10562ec86d6bc801ea32180b17b8c256eaf7fbef52ba46b4b393f5655ca4b4486f7a5db4e097f7e472a20d9dde57564732349be42f8d7687a8293f865e26570e853c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb207c301d597ff6e3f449ffec7427f406e656b002bf768ac5857ff16349f73a330c90e9845de29c82b47d5fe771881bffd5f360192b1648bb8bbc68b4252128bae6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4b54b9edf52abf7a2c78ac9156f44c8951c20ca078e74c5a6f68f3bf7549a978b657042e38c50bb76c2522969fdcf85eeba934e74378866113417946e382d9ce6ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafc8e5eb854efba54421dd80eb57a63d2062a6a8d1c9bda023e6d881d2223cb3c7da01386a06d6f98f2a7aef6294efbfc4a4d0607b8c4dce0e2fde940b8fd908c87f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a6c4905d3bc6f2f12cb64b6f45970368f51838416e2cf90ddf9bae70aec8b46b9b1d59776a1d3a2a923b9e84a263eed23d89f3be28f179213321a4ab8690dfd22a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1beee5bccaf1397198c982a8accdc9982136416d861faabb37877ddf7724ec459d06ac562d4a08ee782da4308af11c6d37ab1fdb9f5c3c06a2aa8b58e31e97002ebaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14940168322e28ca2faa07d9da7b01526af9df3fba3eaad88569400ce2870892d6ea883f79f32558dcbd19fc1e456a45bd4f8a372e641b84c79d1b5bd2c8dba52727d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6ef00cc0333863b40079e900d5fe139e2c760bec503519b28f85e65c094b16641306981c5d989c47a808e3cfbdd82fef9b0c942df9c055811a6d71a1c46954df3d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac2621e9b3f6eb61c6fb9b1af72609eb46fe7b618c82c5ff7edda17289b68880c4705b2b1eb1b8626412091e4199ae66aec9fa4f5f7ff1039332fa7b05d295631b9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a8ef39ea97d0cc2d74492770bd4da0a0795b8b5b63f94244601bd0c59ba433baaef5b17c20165b30846dcb54076af39ab23c066014dfdca9c8c6c2759bd6f28bac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6603f1023b1a5809da8da71379f00b2dd5cafdbe420e9f2e57eaea294172b86a27c2f953e50453eeb6d3683cedba0dc71a9cd661a323b63564895fe1282a40b06cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bce03014f4a31162ec37579cecc4b13f0fc506f0ae51eb93b8a6a185a5fdc2eb6931e230c78eace2e6eda27763cdcccb2d5f833036215146e97186d11b48d12cba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d6a57f06a2c11167236fcfbd22053c6cd2ac3ab54e4f576e6b659188a808b2a209b48c44d71024d8f34ca00eb66f6c7255c790f6f00cbaac174520749244882bf31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b74b42ee555ff4f7eec0c84fde19bd5fedeb4292553e0c86df8100a0dbfe900d30f64fbc8f34461989befa093e68180917c65a216616c59d71ee0be8e4301bb18df1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154fd70b91d1e4833a3276b9638309541df1ee33934b175fbc148604cb676b0c7551b75b84afad69e68851e3b1539677fb572c083184470a59b69398ece7b2d02cf51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0fb0c7884fb7d03b93afda3374335760944e4fb36bdcda6957e7aa007a1a8e5792cef666284b5e602f34d823cf12cf0481941597a2a228ad7d6f603f066a32b50d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85f896fbb1de05164072a9c5552c60bb7e947f325b706280232dea8e0850486acb02df7fb404ffcd525db94dddc93b7908037007ef491011d3b930630f77fd52a94a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae586c5ea5fa998b428e0123847cdf79517d72c67153f92aa58dfd21a3f6d3252ce14240db466bfa5349a34879eb0a85a465205708afd4fb02cc961c753d874dd189;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had6921a872e1d31bdfe956d75c541cbf73ce9c3d30d5dc7dbf41235d04f2edd4b3f81e640e864a3a80b16466a98556cb7b45ee566a83cf672081a68c817dd47be083;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ab9bb42c8ae9bbceec65999abc61df4ac14233f0f1bbf472606efd058e084385d410f2e966a45cc5166d5cc5a0c934bfbc1fc1306863dd071fd837a42f07d03a119;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3aca6bed999e21d25db85f53725753e1b1387c9db6071c3e1b7b341536080e587c6eb59be791766f7cb22cfc368b14d3f1b7139cb317947829381549c6ebfbc38319;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5297217fc2fb0c0de6b322d6d585cf3d3c1ade04bdfa568836178b7c642ead0e626610026f5c585171f362d35e099c24a60e540a14f46b5a09d01cec79cc5ff41d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d739d37c279de05dce38d348431bf38a45fde5c00605a3821c9eb5a9395e90de5a55bab9d218fef9833406b6f53936e350cee5ae6233dc33db3eeaba25a91ee3f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3755429151301b3477c24045d625a57ce9c7e82e85f5e547e4fe95e2fab79eaa6803477f64e7aa6374b7eb7a85a1ce110fb256ef7fc15318ce0960129e6bcc09abcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h563018dffa867835aab0e304b00d15e548e26b24d4c17917d6636b66475a5a410fba25cd485d4a9e7fa228188c00f860b78769ec146abc98d7709838e32b512a5327;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185e5a78d2f30452318123ee2b4b8b990d2342402baf6bf6da67c0d2d51d3953ec27bf9e9c69778474e9822e15cbfa4c8fcc7449af35c11744529c1fd657d2546155d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbeebd5c5fd9171c71f3306aaed99300bcc0950fb9a5bc0f9f774184d74aaa622da97694e35f6116cbf2e63d3975fb07f1ed1e74d46bbbcf20de8a5488076e1a508b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc0d92ee5326e67ef6bbf3cfde4ec3d1e176fc239e717cf9773d5286aa2de32c8f9a5b249e17d4c46752ba6a405cab6ec1566851fa83275663aafc872c40607e3e59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f297aa9ef456bc64436eac5458ff3c91ea83ffb24344844a4dc32a5d8488c5fa21d8e571f134147cf9d0f18f20d01bca3be9cea24c900560a3e7acb54680360a3a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101bc421c950eb94b22aa27b50de7cf4223410574c28adf1d2bdb17a6d5ed89fd19d85a7d8dbcf66de7b2393d5b8bb5a65de53db56615581ba42a66b52893a3509c6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c138eff1793fde215706152f364f534bf3cf89cd3afaf792919f37b19b5c3d7778e01582532945a858a413410aa60b478fceeab3f879f126d5e642f5001833afdb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93f38a1f085c37e2b41a2ec53886331862414b009db67f91fdec7a5b13458a02f65072474a97d6a2f4b80c8e1f46de48f7f78fc6a204676073521b7426c9f2935eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175582ffb236b76caa94af5fdaa29ac4c497bdc03b6628269121ad2e3af202a63073547a560ca551f465f91622cf81d47e8e3c07c11fe3b8d5999132f8d4692efa1c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c078e49532ce4fe288be8104d4ca5dcdd6877ffbe5f6716c1c4c1b2ed3f586dcd14ec872c8da4f042cede21ac8b12d7c810b7cd27d8974795281b58daba4429c36e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbab85ca380ae06e42917e542a34862af3f101ec36dbdc6fc05e64840de187b3bdb5882c8c6bd0b4f87e1cd56d63c717f358c72b4cef57539b450381789e43e20a3db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea103a5b3a48418a65e8b309886d6fa8d1f3203beea652be76e7f1891fcdac41e989ef0b6c5d2a10bda8ebf7288dd1d0fdf6cfbb7b1fe24dede45d24ba73ddd3c476;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98a9f0dd15c2f49f38f788ba9e29615f06d7b41fdb2076a51fae8798e26c241207ee2c6677d971449bf882d9a9bc2c77f6219e159cb6f881354377bdc6b98e53b468;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64f4dc2655b44418906d494aeb69c65de3a57ae95c4497e0e9c3e7ba5de0c3f58dc33160508c9782403b04963562e27fa47e9dcd538e92846b144d497f9527c77de2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4600f74c1b0f6e56bec4b691b57c8ccc02dd49382b2682cd71e6442be0a479791c04430c35b05cd7f064184cea5d997ff7701382f87bef408d8ec80ebf1e3775898f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafb124a2861e0156a35108b4446933a5038aec8b509846f766a649283e3766890335ab454775df9498ee3451272f8afc7086e2c6f6d83855eaa6f2096539323f8ec7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e2b628ed63e525155b64e6a52a02ad7ab012c6898407fd3b764838ade54abb421baf49cb4a103fb4e02153b8e0e510002356da236698dee6a19543183473b14806a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175216d2e9760cc75060b9e20c404df7cb317939eeb0f2192f217ff4d5c89bd4a98a2c597051a35600d94b40ba8b7e435d5097dbbec90ab1f44f0519e9b2678987a11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1504a79d489a4e06eac54cb7d891fd00a01710c7602693f9cb472cf4ef108f8751b0da79f95553c9ae7396137ceb0a32aaea9c550421bcc6bd76446c1863d18278eb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19cfe75e74c14f8c28a4a693a6e6f808c50cde4e23f228da0a9ea9c1caf9113e09b7e85d6b1651c0c98d6eabe93311d66e7072555b9b5a396cc563f7fe4219ae9d484;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1347d9917e04b8d1210dedaad9ad5de8cfeeae9dc85e8df73e3d3106ab610833d2fc4ef0eba4cbb21acb8d895969608241ec5e1c8e87c01fbaf1ab4e5a323e5231663;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e844d9e43efd317a93959939706fece7ed119f7e5d0a8d1236fa20b2d6374be529fd3505524162361a46af81d4178727d49291db578a30312160675542c8d19ef57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h483a63a8d3ecbb75581d21348641bb56064c122c98172d74e1bb54a5a134883b407bea9a62c0b303b9745b813ba62dcdec97fc31e0aa150b4938e8a4785c04ad25ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddd3d772030cde43f2546014a6f66b80b2bf1cf603ddb4aabb809ab8d4c8a4b28e7448197a210ff6ad5125e79ab7e54a0e1d0df172071165c1e0edb0f995af57ec62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1864b6f34293b627e16cea8862e786b3111220f42d7986cc137d467e631fd861c4fb49d3ee06893ebc8891d01df5d9a77914a6f0acfa0a94731f6992f9ec3d9360028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc96eaf7a87609fb3c67588b9b3f3235ea64e6c4b54fefbbe553a365bbff20f12884228ed6340037b2ba117627b722fc2c266380cf34e25e066abb1d9691d4ef502d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ac5d50209087196b678ab9531f92035b700b78ff2d6b66e782361f7a660e59ab089b425f3869004b469b07b85d2d2a5202e70af4224a01d835b0eb6edb8e35a4b82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1bced4832343d637b9a16ca19737b2a113f24d30bbf40aed28c5614b25dfce7dd02bb8b94b14d4c785615fdce530086a50a01461fbf048edfd2129581ae166fc10a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b0f2bf2d3ae01dcbfe15ec04bfbb3c705ff4e9cb28cf4fe49086a69611d119db28fbda47baa855a837cbbceaa8629ba5c37fcce143080619b641424326156a9e9d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bf4946aebfd97a27ab47f627f7a72463c14de28d715fd9035dd086a627e6578e6d7fdd4502cc95309cc7c4c3543472a54c4d9ab6619e980e7e793e064f10461487b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1118d53a8097bee50e755db77aa027afc4451b7666f7f4e9acd6817b8e14a02a7a0ca2ea8a2f7b3dcb48f4469016f068986e4e24a543b52f6c3bf833b3fc88fa52345;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c20cbd99897d8c800aa2bef50ec6b3a825cb7d7df2641bd24d3fb2dfea0aa77c7b3993e8350491c50ec57e11292dd62bac59c2a9bf2d330ccaa226e9d7568a703bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182dbd8130e22ca1fb579ebc319fd146067cccfb99ea995fb40e7730b32fcf072c78a22e5245c428fefab995e3866099805df9895d2c661e4df43ce8d8acbf2cf94ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132e38fdf220dae6611467ff78bf7f84d780e3fdec7a37fad26f0e87d5202d23eb7b149417c8a2d8dd24e6020647a3cbf57b291fa2ff5023eebab17691b81aba3aa30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e36c6dcd42a221708ba4e67d20fa9538306141614498f37447ef23e82b0af5650e942041480f4ea2e7e970a8ed452403aadc59928ffe750095439b3d57e11bbabff6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115c5cd18567e652e6cffc63d7506aebe25636ff3e0882df58a5925dcc067d82f2ce0c3c17c05cbf038a1cfdef344753b5b8f152d6a84e42f47323e39c67b38e73b4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d5eba618307b0b170eafd8d4a45f7fbcbe8401613ab700855609e8615f5a88faffa8449e1726b3d4c69de5ef3d25bd5075ff121486ae5de0417235022cadc90e0fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165ed85dabfaee3c82314fef26dc05060b62627c0361719033e1db7e413fbcd2a8f97f5befcae00811b0dca29bec914876283192c9037124e5d45a42b4341f57d9e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a8fb75c7aacdd3c08bffc17df6da499338638638d3f4b85beff478a44b43fffa8c8633cfa331eff4cd4925641efdec3cef48d7bb2c50bcad35329e6afb62e752b3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd14f452ee4b24803382036e39e6e341025c9a887041fc44845819dad164c5a0374489f6493b9c12a2d11711f01be78ff3dec12c86581d3b74017d0b5858ee6a2ef6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3a0428d86cb5a3e278be9a6c2560b392244de7319cf549959ac654f04600a5f90a1781d470dacd0e1f6501363c5a9d5080fc1362a1e10452ddcdf4ecb8c9cc56976;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8eabfa64be158a6cba704d0d7102a65668a7614c60ab4cd6b21342e29521f6f9a24bbdb7f5f814cd2233dbb6040a7b7c53d6571e57d3a7d5e23a61e0c9440e61dfd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc33fad55c155e40f8a381038a6e6b52dec13154b79e564bc6992924a0084c2e1a9154b9de7feb72a851f40291fd0bc08d8ee3efd9fdc46d433d21b33b5cc708c8d77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1193c9cc1caddf986bdade99adb7164b086cd2338115a208d0bdf7bb754ddfba5b65c2e95681dd0e06eb29625531e22513b2d0db3aab0ca075179dcf98796e35195c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h377ff644a2e241dd1748d12b5608f0e534e652eb46305b767aad469cdd0f07935aa4af29902596d88ae29d19b35a090ef47c0aead2f367bafa1425b189b928a10090;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd21a203001f60e205378b8e5cd11c2c5ae1c3b6d475e2be73d8238ca4ed8d64c6da96268f6c59f95f5780d52279d1178462655d91ab281b5acf7ca061dffc1bd38a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce6c646ab351a3ecd8875f446a5212ada7c814992685ffa5d71f12d86056d99cb04dfe17db0bd2d8bebae7a96810c7943b8d94e2445abf10c5c8a05a441da0e6b762;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b7321e4faea904a5e6a49ec6d874b67ac33e220e28ae3ba07f41f4237698943a6ea348d7d88c888f782eda694a994ce8cb45c4fa24cf96f7e32ee7c8a55ad0dadb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5b6353d551e2cf6d79548ae0ee91c57c164b4f303c3d1b81210dc649c4786c8d810eeb38fb97aa6eccc8bf0cfc1908660caffffc3ec1d0984ec9d38e4b384d5fbce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12012fdeced505f535ac8cdf005f5c3dc6a312ea0e801e1c94ee9febadd8972f2c454519354030559796131945b5dc4457fcbf4156fb009d283f029f38cad6c8bbc69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cffc631facc11acee5ee1702f5bf2c1a29a007a60dcb08559d2a210b38d0c504a41b4581cfc0eaf76733a59a377709ceb82ef61b5ea779e16f25a056b1af5ed084;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ba5803ce659abaeed2ed10c5032a88815cf8aa7097f47df3f76e759d1405b0c5076431037ec43521c64d7a20cb1a29f4c51270d834d15383e68b3bfd96a7c3cbf7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6d79c75da0e5d8ffe6914c8051112182b3aa59936e135340c5c12375d34b51eec6ec2620ad7b06c0b23877c9afacf4d31e85d7cd4b6f860dda9dc723490a88ffdf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb4ec32b4d2223afb9a8fc6581b70fc4f6c9591dd1bcfc8ee384dc4a6c632a844d9ec4024797076747e00e7cd7ec55c2419ee3bd42e3a7a50eb2741f7e8d9b1545c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1617ed46b5f83e8bd6d7a6a981c532ffebe642833a00cb63c8186afcbc65cb3fc5278be5853d3e4bf1832c1d05d0a85245ecb7197d21af906be56080cbb086103bddc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127908a664994bb9df714a929923c7b0ae4b1bce87883dbb4adeec15202da0ef00261137dd33e049755b6ba5fe4bde81daf5049e41a6babe85be91689b12af45f4959;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136b3b66dd5763c07bd9ab8c76ab9b3ef74a39b932512bbfc10a57066f9fac31d98628633c268c9f47d8209929a5c0b798438b6dd8a54676ef8490e06974d6160b0a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a24ffdfbb1ac446ee4bad1efb0c423fac9e1ed82adfbff42ad7eb80b532a1074c96c1fc51b3ca779a799d06e6ab5f1084d2905aa8611f5a7e7d591148e7a8eaf083a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b40efbd489ef343a57c70a0ffbecc6e3be7b66ef47e60425646d4259fbdefae6b369761bf33e7eb24e257a3269ed57700c1a6be5d03d26314b0238cb067b197153bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eca5b8b37c9c67bc384990aa27a0781af8c7d2081c62c767d5f0f2a85070aa9e87a54f7fb439a0104114947c179c44beda66334d5e0b21c2dbf1b0955f8c43116570;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1827dd0fb5d83f595d168f8e41622643fe62f1ea99818cd2e3dff2a10a9b8566fcabd0797a605c26d8bb29edf044ad743b3e6f91433cf06df811e9a3f41f33ac42572;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd49fbf4c038d979debf286087aa519bb235c4db7af0c86d50b866310dc0fbf96ba2c2e33248a9aa2fb1e21e7ab467ffd444a365cf6bfcdc75feb4d1219b5fb02cf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5b9f09561a04df00d47a811835bd95b4f57856bbd924dfe277fb24d1318da00440f72a3b68562ef6f3e937aa8fde1ff5dcd66c0c06cef984288be71ffecaa85e823;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8331bda41671e43631a697c053eb32ba666a7b84c36d18ba8f4eda2560bc9cee30db5afe521ea1b135773204ef4d4e5301d4f5b247107844349c587f5ca773d3fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70418dfe2068c328d8160f6edcfe7b26abc4156f67b80416e60cd5d1125f9ee970aac4289112dc4e4dfa23e0f0c507ee0b0deefc917af4102bd4ff29557b41f14cc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4a2b970baaeed4bc3e089221ba7afad39c614952ede203e5460577b9ecf2f07aac16f84dde59a63bad31be14be67493dff136b325496921bad711d571f70cf066c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h929acf1d05bc69b34bf609b5316972e5f0300b0732e3604c8cc87152dc743e2a838b116fb82ac1b97d96d7b2313c0876ea456bb317812f2ffdc2b9bea1f7caa74c52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a7f2e7bf92e15042c8fc3e3b124a7caa00f3e2cddfded18f0a4304c7d315e651a19209061edb0a364744745492a7ce28631d4fcd170eeada77e1c622486f06a7a06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdff0feae7fe2f7ac8b2c5af1e99d8395a943ffe5e53290f14f8b0ab530464c4dd6c7f2f43d2b07cba4fc4d234fef1b5189c323917adbf30577d2ee2275fbf0fe35be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ed86d65bc7db7c14f2570bf369bdc60d3113f0d5c3d82efb348e04cfb2746f4753c43c18fbf311e9d779d2cc7aeff7db9b8d56dcb00f0d847677e857c0de41272dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9b0a07bb0f8bd5de718a495dd05b01bb44111f44deaefc20e317baf2aeec549d44437186ae4e8a728d996e682c9721b92080c9a6c060bc7029438bf97c57cec2116;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78f8cbd0a335d65940ba74e74e53d5fe4255abb075b6aaf4217e884f1b8a59fa2467048b0145dee8a55fbf21cf0bf7309f49477591ed6b2975505512df2d3a2904f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26c5057706914ea842e21e5fc7a09a4de9d2d18e76a4b5804d7133847bb30bb137957edefc1851e62c0ab6561ec3101e61996647614076da5f6d41d46efdd5c64ca2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h728864bad6fabeaa2d8f629fc1a74834e6f38ec64934c3a4154aa60b192865fba4ab2da4254bc5180036fd953345e25025380717e463002f47a899136e334c8496c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1699d69cf176d546e0af2332b222760b5810611ac3234e9c30910c0b9faed25e34d090fbee4fe6e4baa0aa4276ccb3474233467248b8fc7207dd35925373617fbdd56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14119d6d8cec4d937dcba1897669b256bee0fe07d013d9645c3c546342f30306e285e760a7a628e384d19c14eee24994513cdbc417de490bce565567531210c810c79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a9ee8bd3f79349d4ab4e3689a655c022bf3bd76e2a7b7320008850e4fd27ad3dae807089c4ae24534d9b9d5d27125aefa23605799aaa274b6e33f394ecf8b3296f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67cdf360c8b131fcac6aace60e1e46e66478be7d99fb37da5747d277aed3658f717a5ec1a1e2684b8a3a97a5266d6c9c1f1e8764ea38acb55475d3133e6412555e74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134130b99ca2773cfd55a14046e27ff484bf602b992f2c1a1ca1ea7f1f6910a1eb3b06b6cf3c3773491a6bd014a1f809fe8a27ee491f43c2ef7bb6da7287e23df65fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1938e24c68c96bd866a9f78a7cc9f8a559d91d5e3285885c44f3fe63b88064839da8be30697ea8cb46d48745a042891cc589a710e0d68d50c6f02ef8da9fcbe6fc32b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82d1ed6f263d51575f620a9c4de7d796238fe9848574418354b68ea1c67a50c5b5a75f9402e142cab8040f1aa2327b1c538874056f3ba2ac22b224eca62ed11295d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b4e418e84f7f3c9624ede030b7c50ecd1850e20d94d8bac062f208f0d2d94aee3b36d72f8f0095e31a2b9cc90d5057a59bed66029672a31f944a2c25e6264a85777;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd2f10ac5a8209bdf91868883086f85c18f7d836a7ca138207c80d84ec9ddc7218a810e8ff219d7581929470e16ff93f9c4d80fac1d98356c331200c2033042a24b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf61a98e890b0aa86983ffd47ad2f8e177c1ee43eab25dc4b6522470cf162a7ec3b059daff63757fde1b15a007802709c518fe968cfe1739f74ab66d6521f665bbb1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fae16b36688aa173cc36ec5f992054196a7a9b6f49ec76715117f8f416b0305e29eab959df992111f3795a81dc469387e60bbfb764c76521076f6ea6aeb18fdf35dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28ba413635d31d51a8c7ca91471d98c8a7c69b29e77050b741c2a5a4620996b197bfd36245565446d54e37f02bd0cd9862766f7363b7daf5f286207a74571e506604;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193f8a94dc3b0ef6e632556c2a1411cc3fca810a17efe679220f78a103ec3fdbf2ff5e4e99570ca92d0517af05a09b511a6aa3e8e2c118d74f9f529ee8f1983c81287;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6954a4ee3cdddf09058519005fddb64ba10d37a6925cbb5912c6d263688293a72c6e6eec05caa8d67969f51b63cdd03e30f6104db528ceda4cd0e91ad2c10cf7190a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9ddbb0e6ebdeb8236cc0c9da75826be9c190fd8d49f439ea6011d8308d5c8ec52b88fcd500d3bab8351b9cb2b2f0b098469f2a36af6f2d51019ab8383a5eed7f27b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69a5ab82bffade8de1f710a35c49e6c2225faa28d821d610ea6ccbda35fe5afc90827d95cec00094a46869a2fffd92c65a4b257ee5d9e8969d364a722aaa45252327;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fce53f17906bfefa867cce628c69c2a4bc80a65aec3d8c080ec0c39790c6816b8be3fd02d63ef1bd5b33bf270860cb341ef19ff49f32cf8416533116b8d74c9a20a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab44b23a79204d27eb74a5b4a45879a3773eefa324f1e20440a76267ea5be319b0b20caed60c29f015b7a25eb54fc25adc0d1ce4d03b2c3512d9e818af45a6b6ff3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122233bc63c3302597bb3a0344a336e5716a322c0aeece69eb67a918bb15e4b6311ab19da3915f180f7ea500621cbf34d2578afe567a3281f46cd1024154329243711;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc536ee8fd82a79b29a8cd2cfa8dc2d9556ce96a692f06cebd1d5e66345601cf39b1f54a10ed9848f02bbe696c518fad4651008ac4231d19e4c477ed3fb5ec67bff86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda35a39b3d1723cbdd54efefbab151bf285e68b5f04953970d193babd79ee8e6ba13067cd0a3b5e1d45e2a8adf149fc5fd71adccb4dadd6ca0c839f16b5d20559501;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0ffd51cdbc11038234a09023b3967ce3301153c6b455ee332262e20da177f5073be0e833c9c913f2ae7c312652fd7198992478f7823c0a285bc78e401a6d4af97c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edff8abcd027c226bcf68200129f7781aa7c61afded02ad74cbabb0ab9909efc9de2fe52b6a69af0455c3b7d04e8ecc51b76fafcfedd14b4fa881d5822e5f861e70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb006ff8f185006b2517e01c95e17ad638fe7bbd5cd82a53920db19e6a88b2d5dd90ea3d86b932f71865bc5738d375e6eccf7f99734fb2c6887dc519d6119a765b253;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed944a1d5aaa4f22c95cb13537a93ef4e187be5a3c8f5f2103b7d621a6c9523b1c6c0b144c6977f0599df7bb2523f6d27f246d5fa98b2280cd4307981fc7b5a4db47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1785d8dc09aa8d78ef9d3b991dc1c73e389c9dcb18edc0d2a7c7368a5ec426448ac52e6de05aea99c1aaed465e05e65b87ea274750246aa25f0d6de336ab5496ded14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6063bd66a14a8cb81699963cd5ff253717e8420024b737be156fe5807447010d8e1b3ed1ee74288dac8459db46165de334c64c3497cdaa241e08702ae7779c6acce4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c27eda2ea6350dbf2922c73431df2f5b3cefd7d0b261f373c7dd7cbb6e755f613298cf4c475bfb079b0f75a3f4b86283a0eacdc2136700df35d32a92ca4b4c54e6c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f48b2fb59410c0ad009538dfe648a80f70eedc0b7913f8a29eb4ab00296826c12ae90b386582b6127a9ac8c28d608407f0f300ad16a9f57216f615574f5f2827cc87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3cadc24e7c00accf3fb8ada386eadddc442c5f6f3f364d67f34ea90403950c9588d831ec705d70ac61cde2820c3c255fe7fffa73f10ef120bd5b2d96993114f586fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d17784de1282ef9d11f9c3822b4a7148e4b72e8f728f1a0941584486e0051486a32ac7221765248bc7f05a5d0e85458dc64f7a3dce35cf9825aaea7ddcedcf9e89;
        #1
        $finish();
    end
endmodule
