module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70752840826fb987b79b6f6bb6fa359088f8eb20b31dea501;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93b90ce2f49eb9fee1ff67de8ba30bd9cc9fbe42e0cc95331;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcf3326d9124b0406e8f8b0f4185ecef3383e09af17c1a011;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haddc31d3cd83d98ecf9845e00a63252a95fa3259fd527e482;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb28e3f1dabdb0c452ba718a447ebf28086b485db9f083b14b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bbc498d591866da064aadf9153f7540e04f09648a133b238;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68ba6c612f61c34d3ce9da6b3a07a87fb8f45d3a35fc0a8cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92fb2df95af7370416349c416f1d86d21bf6b497002f6adb3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2e614a98398d9839f043f5953e05f4eb21de2ff54304f263;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28b48b0d38ab110de0bee859138e16e79d07be3f7d731e818;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h714f3c0522ac68a770b5f54f2ffa6b694e0e5ada82f9d95c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3e72313f486ab8ee85e8d695b1720cf781830be3fc75eab3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h755decbdbf445dbe9132b99607b7ee166d98c51fddb9f1f03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4127a7ba81e30afae9ae0ef548639047c83f8b52d566bbc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c0f8176368d9395a2a8ae383fe0cd598abbf8dbc921edfc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb09e0c52bd0bc6c75397b4c2768a44d3b6afb79c6baebcd41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8097c94d6be1b119e3a53ebe287b0680b0df9de159a3b21f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfef219d48fc0de4e6bec3e882168aa8e5889b1b2a04dbcc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bb320183b5431ec22c07c72ce8d0c9d324a1081852aca52d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h998f31a38c764fa41c8f2525165882b1287a079cbcb86488a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccd3995593b1c4a329f2aee15213ec90f2e38cd1cfe2b6b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf125b3e247b18e72c6bf14167a3c84ae7d9654b12ea916611;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b884d775baf38c135fc195c1f3c8c815fbe3c8ebb715f8f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf78338133c40cec034af8eff0d3bfaa50ab59caf0ff9224de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63994a5c519062c741278ce8707d197bd524c98202ffd1cfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0bd009d8f246febf4af7fdf4f9b0984836d87041bcc9ba88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54e7b10991aeadf3a79e027f6a78e299d30ba21b73ee90736;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f7949ecd102dcf68f536354c01fb408ef040a3081b3c8588;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h382185ed13f5b202550ff54053312c0826900dfbbbd8181cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h972346a87efc318fe752b007bb444e51c6597d2d0ecc1f970;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf1d40c79ee2f792432f85c4ebd785263a33abdfc743640d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47f528fa9a49740c2205273d8b37366dfc12f37d0bf75017f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haebe765a90ded18805e104379ce8801a21a723353e68c8264;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d0a78b1769e201e366c26682e7cf6dc10b4d155be5a7d0a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44302784697405ab7172a8968db6f119b6fc347570b06602;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h228302c31650e4808cb646cc155b758f6bbf0ae22d0bc1e05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd71453b98ba1ce3754f28eae95abeeb3fde1d3fda4537192c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45f467c35e7511fbb134ae4fdf8e7879e25965aaf3bc0b2a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha99e9be382dcbaf0a1f89366da14afcfb508fe18bc43cfba5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78ba1be3f2423583fc25ec1030bc0de974fca33eddc620fb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92c258efbe4fbe8e2c38e7161e85e2ad7c9e281a99ae3074;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h209640dd3b927242678485f042a1fb067d6b2da74138c80ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9788182f6938148c38e3139ebfb002bb72cbd987b2312e13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83bf4c12f86ac9d89446842f3757df84ff92a3544f555604c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc2f57321ca683cb616417958c2d9bf75186a998701b288fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aa60425455f3712ccb8f7f1b8b3cc8f8a6e0e02d9d3e85e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h760addb663d553d28c9353bba51088f4ba621d804c178829;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84471faa41414cc5433f2f4a831d1892d3a160095c896ea3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78ff340204e2648eadfbb9fc956903566a4df2f45f9c7246f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3891a8a4f6efd9884604f9a66ee690eb0007995412bce99a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2742df5fc7b64a259b009f6802deac354b35741a080d5e099;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6741d7c7a77ec3a067aa0ac7398199a4f54fab71f83537425;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51309cc9b0cb7d4dd0c85aec2cf0df0ca4b78ce3dc5e34e73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9be5d95408835a646821a687eb7bc8b7334af3d0e082a363c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h219241e9eaacd0d9c0f842ea3e5826e7fa7202be2915662ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h399d41a084b2ffafa283cf3b5cd2442c23aaa4c05ccc7a7c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaf7211c8a115740ed1b7ed787d6c15b7579c9ae32a52f8bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f57370abbe9b9c82539c53be2ef13d63b7779004e615c5a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha631b23abfe12f29c97ff561f4fb6e98ef8ee207a72b32c44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4144aa4b19d10f4076c10d0a3796a15550da000226c3c4b27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbbd8171341bc9eb726a94f0b006c39208185038a1d6f5cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcabcc0947f2b801c6f613daf8321f87aaa42902564c3db216;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a432cfe7edcc2e79ef757e4fee410e594bc630369af8e6a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha97e577850904efa20a8b7ebb93a2791ccb68d47ad04de89a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb170b61e36d212780f89615fe01b42b044e81434a633df450;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7e87c0e04875cea575c4d1d33c55ac4a08381b712a389e60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a34cc7426b192150449d7b0bdbc480ffea2d3456e810e6be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8edddc5ae0f6ce762f26ed795c4954e5a2ac21ecbe3e3472f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h126584f49f2c7d51d6036843561676cdef71f6ae5415ab62a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba58fb7965841ec073838903998724a6c2095876b2164a63e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d97849cc99b39112b647461661012f04720a817f22ffb237;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c19ef663ecabdecb47dd105aaede0a02a9f9462a03e7d47c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h200414c499dbf6d28f0831f111f26f348468dc10aed4a73ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fcb040490a7e6a4b5984b1f46f0aa1772d556963550e6972;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hace52593b15f310d4debd321288d545efc6dfa96b6f298aa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0bdf4aee477a6a25cd1a76411d3fe72196da3907f841951a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62704f80a52d12fb29a475b389eb3f270a2e34f30ed2d6960;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1d31545152f4883ef49a7e91bc9345b6b6155c8601196070;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h947d98114b9ebb12478145f96ef74519abea64bc8e74d49a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32ee0a6730eb3be97e6f4b45f4612a8affab1e43547490080;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96e56f78a6bdcae1629054d353706b75a054e0ee83d7aeacc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48ff6f1244e78da14225f5063f251357711e969e4f5a06d83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2036e4c7400c7757f4c537a1e4687c710bfb768a62cd087c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h515b7df3d1518c637db4735b5f35a7335e48c2966238851c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heeb720ab31954838d0b64b7f48f198f330bd412416bb86cf2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe535f7bcec5ff47c3a9c8eeca5b0840f3f00fcf60c2b8129;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd572ad0b588851a3c7af5b16f3251015afa5a1d4632c138c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc66db7745ccb1b8ef1d669573b103639ce8ced7b7b4bb93b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc56e022a954985a1143989430625c8fb3103ef2141e68eb25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf74c0257357522ec207a833270d130e2e4f67ce602bd50302;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4df35db154ba51552a046e8275d9dbd0bd88ff37d0be65b53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc85041fe29324a579dffeba6a6b6d04e7add48cf3183a2079;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h354a4a42dd0c8c5d33447b29341ea422b19e325ce559dc5ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4a38882391b80f0cbdf2cfc269e1ecdcfefdee932486f533;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e418676b326ef4e5012d2429a1381ccc483e1a367c19adb9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e2931cf2d8b5b924635e87b9bf75b12859f38f3949d622f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5ec0dba46747119fd3e02c97118f6f80d6c65e8ea46842c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99523e979f53fda0456ad2456da151e6e1853d119b8749d24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4fecb7571ac508e11ba283082eeaab20307525897af7d7a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf612ff034b879b1979197bf5dc4f336e81f19bad1c4192e72;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc261b28063dc7323d4a2c8fdae0cacb636a1f5cb914964a25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b3656e98dc662f92bffc28431cdfc515188ce474fa3fe78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h695d8be04cce42559e933090a8881794f767118ab2f1afa0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd86c54ddc94cda82d6aff8d37adb3fcedd9693546d90c41c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3abb8b3469c70efd8d4f1142123ca87db4512a6d90e388e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a21487ef32f3d6154fb0c3a651f6e41d3fa9597e77865b2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe455b745a2056e4e86309cbd8f7d2823b252425957954776;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he65d7aa0f725096771d87d969d8a8bd0ba1a76140fca49ced;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h195c25ab4f29a41fa72e4779d0558c034d3d65b6980151be0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18b4cf30615da2caf2590b500d6e0ea6d0546bf28a0b31ce4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae27a8a2fbd4bab91279aa3b1a6f0a3d3db875817695bd804;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25fb61500df97075022877c0c022f2c441ecbd899302356bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc547745fcd8263cdc7c5321c979a6e586c0046b60ccc33947;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e2c6abd10245507de0dd069dd71ca43a8fc7957296cb57d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h331f4656505d4cf9b172d4d1446f9beaca2ed8a15108dedaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h942a09d7e00f419f864cc9c29fa720649cec2c1f4a3864131;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2d5d344515d6aa16b3a1b6bbd4b05ba237c35f6aa636d999;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h242e35878e260d999545bc3daa084a4bd01eb4d561317f8d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52e965badace8a94a50cff631963b4be871a4ff781f4c4420;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h966cceff69206c048d43998fb2d3fffa93d6ab6854eb00e40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd556b3eb9e241c61c2453593a631963fb415f2cc6f9b84a9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e0222dedf3857a83674ea5fbf282bce79308d95b4b3e32cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had95206870a993b78942e2e3cd17888333c5bba4092b00078;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73c216cea3439fdb5f45f8e53c4de202e3122fa40ce878a41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73288f280a7f0a16919380150f1e15f873288215855708dab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d921cd8c0851650fd8474ccdc6b7412a269bf03eb339dfa6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h569434610a9100bee38f9667d0dd26f81d6ed813e599417ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0263214e3a0a201c099754eb5fe51c97c1e8927ea34906e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d582e007c8a5b50962de4a26771bff3311f1b7e644db3dcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb5384f75ab16289f3069243fa6700acabb34466d16d9318c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h393fecf914d29c89e8d35007bee19de0a39e27a1e74e64b7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff07d7e6ac5ad1b81d4a88bcc415b05118aefd62d64a66a45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82bfdc9214d907f23b8eab1de9c17fbafc3a9d1fa1616647b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73b092f956e291c376de818a2f276507411f8913d598cd4a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ed7770d3420f7dc2087b7ef8fa923ed479672ab923cb35eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11fbbf8d7a6ad52c21c781932383faad6a53b1551564a5b53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0f4ae14dae225169af88f398511047b6654b057e1177cc84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b21228234711f89785fb28a9b0e14a5a1c3947aa3a522c00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bbbf9b4e71a0021e20b3482204bc7f4e9e1c26557074bfb2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40bf64aa988b45dade59c8bab5d525bfbb6e22e0741003a53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e494172ee9398e38a4c79241a53000ea5865e6d63f8d5c31;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f50d1257cf9efd538cae1cc9e6bfe43f4f08d81a1c77aba8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89d22dfe12ff7ec18043a11ec39e5d4d65e6d5867398681;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29e4e9aefb785fb786c1aae79362c487692caada86cc018f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63d8d14646bfcff4c3989565ae6012e2d74d1faba77df869a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dd888dbd94738aa8ec420dc6b9dadf2f62b74ea8b2d9481f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbcb694148b4479dd1b067b79a9b8bffcf57208c1f6dc0142;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8835d6d331d72ac4121f61898784782214af917ebe08eb7b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8546b3e10adcf176d15217d6029edf4b14caa0e6a68bb7a43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c962dd6bd26189af4b02bf299e1046cf6944eab2f39ac02d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf63996af84f6b0be25e9e4a861ed0d656c8c90e10c3269f21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b268ea5863501a837f4dfd47b03aef510253ba554ad381f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1dbc8997e5f1e36c260ab78844eb15b099f7f1588d8f65d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha88bd4e2c9913b591e3363921b1d9e75ae8a95a54410d1ddd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h276d60d3186cf6c1203c161f8aa9ad581f540eebff0215061;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24314e4bfffbe41cf2169d8a94e2645dd63ecc4df93a1acd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfda366137e3e2cf8b18fe62fe695e044f7620a5fb54bdb2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58c1a1de8f9e56d621ccf86fca824986d3322e214fa2a880a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he13730b47c4b743b96a2532f2754f393e3b772aebb99482c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd40fd6c81a368c39a87f8e332e7ddf22a3f72a5c396ddb890;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5fe44692ec799ff5b75f73beb62d6336b584affe5a07a558;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7e4c68f45caf4ce38e777a1b6aeb49a969a4452fb04a35a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h972b80d7ba537c307955b6aa2be7b7055d0ec8b5ae9eb46bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3765ac2b59c0780088caf5d28689985977888141dad878105;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1027589a0cfc0eb15ed5ff6e413a13efa1fe37cc994004ace;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4492de605f083834b5c1351a6f8c8bf07726243537bcd83cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71a40d25fb0ae2a3e5a6bcc739b8cb6eb0b9a958df07123d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5351de533f2834d987200c515693fae68a63416f8daf8ec80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha45592ddcb29829ee89fe8b8843532015075e70e6f45cd8aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he746f0b059bf2f02651776cfef06fd2754e5cd8699e1e5198;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e657962b24a618aea2e2ae31048732de0d6b6ada78e3f8a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d4970242f2ee8ce4ba3492790ea8b6952022cfd523106e2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4cd60a9bbf4a05a5ea62b2dafc32e4d4d2159ec57dd11f81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dba075b81d9f0135d5bf9d14a719f3b6c63c1a3bc6e9aad0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2206025518c8d7c20283fa09015289437ccad3f07185b4d34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62b9a4eabd45fdf51841b3257af91aeed8016bba844c3c633;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71449aee8f0ed68744fcd14d6a51f8954c1d6cf36a3456e54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8184137918b0dd99bbf1a912338a1ac0f06f882864b9381a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd89edb2a2523232220590926c3f22f34fcbb76200a795c406;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95b8f750048c8d5a418ed561431df3f9b0df27f107b2a4442;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f6be3cb221ef15cc5671a2fd75e5ccd8589e74944dc26172;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he07746ffc649e010bb13295348ee1e182d23cfec7f48c8cc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8026b20af97e8fb47f746b1a51e18b70304905841ec5c195e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbce7a1f44a92fef285c9fe25bb48786f92591e4f76e80e79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45fd546a55829318d331a0dbf34625c07cdcdf25039f735e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h636d1acb8b5f2efc0a391394214ace79ae184a31d05f6719e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a5384bffe2bf1d17e864221fcf4d9b2c0f2a42438e2abc38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9da3dba2277b339bf8ef18a6aaf7b3789f78ebf46556371c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha90f0c02adaa0d6e89ecd22e53e199aa830cb85908372f026;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d5942ebf080d6d8c2dbfcc946b527d206e54700beadcd11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a91da371789051aa05819605c3c457fe7b9a73be00502f18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4107cdc73bdf5e0dae8cbd964af769f21a5662bb9f1e1c689;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf09ecd67e45bc869548da96a92972a5d3f440d1b957c1151a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8cd866a553d37d530a9d1d6b42c75da6505fff1dd91d42c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cb5e023146868189e183c8d47f6669090b5c219f0228231d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e8b6daa1c9b2654d06904fb22f1c08b40a10a283cfb6777a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5b8e3ed421dd4f9428faf6219b7964b5f9b18802482a0682;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h356cd393899ae245cbe8c5b64c748fea9c268785c51a681a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f25fbd4311757912637028e396afce282b5789963e053688;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dea1031e43b1becb9dba2f338b4ea9208eedb22eb0ce35e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h413a939d792271ac8162cd8a2a159ac7862b0ca20b6af5d36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb49e521eac511f935fb7142b94548c6382eff18991166a112;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h887f604b43ea76255bc8a3f03836a9f296c2bdf3118d22f12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5780499be761db023af452b0d600839b383e8621ddba884b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eb56f029d9cab6eef540791cc3c30c3d3997f88794ddf69b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c8dc509e10ad86555d1138d6e4a95095c9dafe710a9198e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7e738cec810c93431e092860e94094564a27f6244e14479a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1126c355ec02496bf1d08bf06a4f30af07ffd3d672164ce3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha97b2bf00abe04522c882c4d3b8a827cc60e1ce3f61b63a89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd793bda4dc2048e8c31f905af23da9b022c020a89ec8c4fc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d5fb074549018f5bf066f9f54c71ea012fc7477329e3a68d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5397956ebda25c9637bf7eefbd64ecb552da0f6b8add370da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33f1222b99c0bd86f22448a540a7963e3ab3ecbca10c87156;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8c1ee3645b5d022b8f60240a8ce8deb7bbf8f543178c0494;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h899de9baeb1c8bd4587484b0f5435204cb5a677f3a392c1ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb65d88d2ee16ec1343f4e239aaa751d172ea38c8dd6b0faa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c9cf7de6e915784c476d9e7336cb53fc4b48d750a935e325;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd730faa55a05403b07d323fee525f573aa7d587264e581507;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79fc70445b26df0fad10307b6a505c1b95b14d70862bae161;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95aef1eb7acb02b859e16e3d25b6f68e91f9d7e62cb30c49d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca2f1d295c1edaf3ee9a112fc49867500f5831cdbcf08eb98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb817912941784041e03edcbe4efc936b8bdac8c7b09e2b8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he744d06132fad8efe749955eb5102d55ee915c98e39570d99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he428f33d0d812f496b38cfbf1e7772a6c7009bb77b94ead41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf561cd1a094b4f829437350a1bb93f434655dbaa7aa9476;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40dee40e7b243b35ecedf33236df6c5976eb87c67293fb630;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56686627503789a5365f7d9864c294f964a66e552c73ce1db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h142b2995f746ed3509ce4c0f9f4d11f2cece252bfd1bf585f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60c6db3d3f79364e2bc1e3216238963dc8ddb847568da1bcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h661daf434f9637a4a749d2d5e3d15c4b2e474d2e8c8871853;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb37294a65f7d6e3b031fdb9f5d2cc590796a78e1eb0dd1fd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8eecd729d4133fe4a9371ae5b4e76b97e1368549a0944153a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a2b49d300e5b5ecfd32e4f7cbe8c1e66d618e6ca68667903;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcae1121138332e18f63cf23f453c3401600cf9117a1f719;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13ebab169dcc1806806d7763507cc136433da0ae21c715724;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98f1edca48713ae5481414c34995aa0c64dea0df7389359e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5c19b01255591fe7834665cce41044e013de9816d1c160d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ade492769cdbe37fd09bbd0ce5e2ba7f9b401e4e0ed763fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha53d7e3da9696e2db08160222832a9f24c0cf0d4ebad1543d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5710e4bd818880c7be36010b77ed0c065db71253e9c670361;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f5032ef6681f361c38c474af90a0bc68cdfc774748f789fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72c203d57242becece3e6ce6b4911ce1bd27b1791481bfb80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c2384379633f610c5312f57e9c249494c120eedb63a93a2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h343c510620b9e4ef9bee1d9a0bad328b5fb823d90aac30d8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h324379360cbb1d4e7a0e1be553a7a1f501a772c2d004205d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dec153f6f2d29671ba969d96e794b67617587ab84a382c94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bd15e7426d9c80d96f06f9b3386a7d4f112d45b83256583f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93c735930d9e80e4fdf051011b68af7383b71fee25cf354e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ec3f87fdbf6099dae540bc25f2b378a4af01352138bdfff6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96a53e15d087eebc64bfcba6cd4cb7169e1533133e071f27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he62db7a09d1d055f72291623e9d2aada28d77940d08f0db8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ceb3bcdadf0e2cca9ec444f001e7c6a2aaf2ae70691c3bd7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4e10e162d4e3bd911e0637f5edd43ee048a3662c05344b2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61739cdf793201264537b5b8a9081c1132a7694675cf95892;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6cef6936f15b4b98fac0527f01a2403906de430f90ef6626;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb8da71a0bc6170a5d40b7103dee76c63d097d7aa60b1abcd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde2987c47e987237d905331ac5a1e0815b53b44c6ff7acd46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d66c9e2670fb954435467cb13ee902319a9b7aa2b7ddbf0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h133107c08b04d289f2e09e3155e2be2e8b42a96dd79c4b408;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c2e7fe3afad51fce1c46bf957f9e30c64d051b85ff1f1bf7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a395f60afe1524dbee19abf12faab6ae8e6257e7d7b70550;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h229424301279342fe3f06db422e82d2630409062e26b29a76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d5b239c1531b32edfd503846def9ffb11f8798d6a594f502;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d66587b5b626dc3b36b94008c7d45c2416e3dedb1e023eaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0c3441224251d8a3e230bd7ae921c792deb43384be1ac546;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e4a761feab2437a86ca0a21afcbc90ed6520c411d1aef159;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c0dd6ec01df289ef48a2f45f6a73570a9eef85b6ac87524e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd8a1feccd762032d19629d0d571053b83ff6da191a70f939;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb806183a96d19b9bd0205db44907606574572db6ff90243e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h673b81daddf6d2b59d076a61931c96543e19e4bee78f2a722;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38231a767be257ca80022085e8c8a93bb4dccfd00710385e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58736365662f83323ab4751069f6a221ca5f697dfd6bdf9c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80ad887b2090b8b4112975b2dc18d7fabdf0a7dde37157f7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e3f8f0eb44df17b04fd439f9b0514d9e157c9c0da899ffde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ce3c5b7799a436f4e3c28bdc78bfbff2593fa90b994d5cbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h590589a2766a2df7a2f1eb522a40155550755aa480648d4c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8404c69d514cc37c477b396642407f15ab9323576c1e1663;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8898c92a77c44d24d0853d2c69618dfc8adf405988c2fc12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93d9f5f34c99765d09b44d2ef42822485b9dc0d9d062f5385;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had1a54c0a7623dbf8b6ad33290e1a97033fd3c5a072878a12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6ac411a9ac045c35c4a7ce9329aa384c596faa5037ef453c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb641e0a80ab793726cc2f331527a03bc9ace0f98854a5cb0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h409bc75f26efc61d0036dccc0d70304fc008ccdc4b028a0f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f906d78f158c6f254753d1ce9816d5466b56017220d94f96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8aca51a14a9f03323dd2049dd57fe3a0d1e503fa925214dc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb554b465a8a1f638c013b30cbf0f6847900efeabdd726f3d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd2939362dac7aec9452d3aad6e2bff907876e5009f947915;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fcce8f5f556ce32a9963b497061b11d60d45a63453a42f8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14985333d8d2901c3bcca56c0130d20508aa852465cd90f04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcca5ca25824ee04b2a6df9ed92fd072667d2d8b2be43f647c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h509d385870b16f762ea7fb005226b8a715cd88f899662a046;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f263c9ca3aa0998b4a954832519622f260923847ecb70ace;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d39988506a480083f5edc074471589396daad0788da6499d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4896ae46aa05ffe8f8ed61d6066bcca7f2277e4cf5f8736b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29f5d8f99de0c4c5c415ea4597a86560f435e97707d6f5c4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc744ca4856d3c9fb55a7deec9193b9d0a04df506acd1c8119;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h595296a436f4b56d17560d7e025a9dbcf04f668389b144fa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a8299eed25f786a785ef253ca988a1b950080c3a417e0f14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h457069a93214a4fa9d1be58007ab72174aeb8952e51763dd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd52ac570996fead188faa9845b1211200b9b2dbf4ed104481;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc225a92e39a4326127d61da761cd108ac2c1de183cd923f9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7790088d8c400e1529591b0756324ba9cb0eb332883330c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h505f843dd3360a956bfddd74307b8b332193ff7ed996d9a27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdef30ed43e83f174da1b8c6684565a6444f95ef6bc9925d22;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54b076ed51e26051f93de1a49b207c3d01eb73e80b8d0bdcc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he39d437cf1385e0b322bf8f72d91c4f6f55eba7d8812f758d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22b4c8c439cf21430aca6c74a1fdf0f7d19a507c95dc5d1b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdd6f34e6484a12df7cf39a2560a76bf8f87a0cda6b78c267;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61f3f21e369c2cef512b59b032d0570e8182d3979d75c2e07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h946c30c8825063acc9a2650ed0ec5507cef012dfcc003bcf5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h308b275a191ad36e65e19e3af0d0c4b98cbfb047ae8cb0dd2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8818615f2f3972d3ce3aca926c21b1fca489dbd1d0b50163;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12340def33374289e3dfb5af541395cbdc5830a2cc885ce8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96e910c32bf7ac1bc75f6853126eaa82095d345273efa5f40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc605a0732df02f76d69b4706501dde232eb1e3d51c0f22991;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f573ebd4030cf957c7408d43c2ebf7f991b6a4cbf3a392ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bd34a51b3ed89bbf48dfe880ba5270155fe050f28df836c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfae4a4b35dec709c1fde23351cd014cd095ea266cb4b9645;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8261cd58b4e1a7557062fd045d2958881d341977954c5c62d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b06488e146d6a3471104a8157624a27ab3dc3e75dbd051e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32db7c4d290a32e24ccd68eec78a39b04927e14b790ed489f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3b2038e5be9a213cd641262d9e71ab67fa9ef602adb79c64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7463b3c533a0435ff54d3df63697ed3260e2e53b293b92af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d0a2290b0fad87b75b7146374c27eff80f7b3a92ded00679;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h236f29b7770af7668082081c9bdf833acee05038b35176137;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a78c54923c4de2d4e19902a33ff2e25a748c3ecb629c2166;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84a4c1fcc36d8eecc9137eb709717917ab9ce42991eb84e5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7ca66b3f46ab3222f4f793df6074b82ca6e0350ae6ef99b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h883aa9d56fdd9a5baa8aee0066c82dba8bd988f9200b23c01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a63e1256b34ec7a31e68174215994a381c68a498f010ee2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66211bfe5352a41db31eaa3dd5634f66ca85b692ce809a582;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96cd97ba14bb885e081b86850ab237721f975c6558830a59e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe011cec6fa5ef24dfff2a746d3a70c356da68f5dafd1bf88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3257918d36de92b563133089a341ee986d5e4f86d95d337a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h810598925bdec9cce3dd595f4466bc9545dcd3e5e8d22ec95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24f5457d88dbea7f2dce43c37c02670196cd351842133e12c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b65fa9a09cec30e29ace095fdf9f8e74d9e9e89e524da856;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd232c4153a5f4bed332f21a495134ea595fa3568d2bf23531;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dbaac19cbd1fbfbf9c2711d97bfd26791fa82fa6486e7cb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h445abb8f0cbc661f34fc77b4f9c2be09dd624c5bbee90e287;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59e4d734ad29688dfcad2ce1b4c9f53a80e1fa31477c0eb43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed1e00fd2f0307a95c1194b7b4cece63ed061e68d38dacb77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb606e58902090856ad234d6e786d565a64a9d690599e55143;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7c00fa0ed652170c98fc4828971b0aa0577aeef9b69107ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h156b35e0729526ada63545e26eb0bc73d9b3ddc26921e7f3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a96464611832b1f7ce8aa8ac2a39e061a4027ed850b188c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d85be71fdc9222bf5c16bba03cfe045ee86b50b4745f9ad7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14c13b967649a9c581bf38a8f3991cc58c2abcec67df686bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc24c61cc6d7269f36f5727f25c2dcf2d6db6ab993bb76e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb761a14725451c9a75834abe38cb8fe89d0658af2d20bab00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h495e56329f159e46e346e268ed0f86ca2428aa34de169070e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ed76a5073ac7909d11163034e53fa9d3f48c4f17d6d8d30b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2d08cc835cd2cb02e045036320b43332f6ca093d51d89390;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h306bf79361a588611d652e61e94628ab40cd0ef5a198e2b1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5746660e4501c9deb2e7cba1c49b91a2efd74fa9293df2f24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9aba61f17d9d49cc941afe73f0827debc73f40bd593bb0fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc77f799a4808d32a6c397bc2efccdfe5e166e4e9f9d4673a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4437032f334ec9eab0e7770741f0c10bec5ca398399b7411;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2c3fe89c0c8c8b47fac7ec1ffa4c35919f6581ce8815879c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h793e6e0a7af4130dbb11046fcc4051c413ae40239fc6d6b8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46ceab62a7a6efdc11ba07c013fcc65b2772b357bd2921736;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58b1c0c0b2c6e5a0a894f33768f017daca3637494bcb249d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5e109df60dc41effdf4b8b76b35f2fb7c04b814877719eb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8021f370783d16ef52802015b3602acfc7b07f2fff8ec1d87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habc31e2796f008cebf766ea2c242c463f04f3db2b0ac68fe2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea3947a6c658f86720ca9ad461d662f6ef2ce8f3f7315ba67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbea38100662dfc7dd5456414d63fcf6012178321a2eb79c98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha535e0ad9ea9ae05f323ed39617d8ac759344cb1ed9546c3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dcf060be7168ad4dd8e768d114781e4ab44aa9c1b774a78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf83f6b5de082c03ae777fe7271a5884c77416e103afb16925;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he02060324c52e09b4e526426730c6b6d19141f6d74e07f46a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc326d125d9dc78217da20556ecf49798caed340d4c3b0f10c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a257b3d5532b9935ba397d6d8d1e832937928fe6d35f2867;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1828abb576b20c93262116bb65f89efc3f75fcdbe3cc98455;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34ead0277537603d36b6bb4f97b4d66ee7e1c71c75edd5f40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b51ed48166e293fb7aa1749cb6d907557c2afc60deb8fa50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9979abd26ad62e0e4f69811ec9baaf15de7849574a32f9d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc14e402633d881b2841d8b914fdac59783094816fb77c762f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e46c419dd06992b514b5d976ecc827793c7a2780a6756752;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99db04d3c4c57d264d6a052474aa6d20bbc2d5076dec89d59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5867bbf16652c963c8d95c85b8bcdb30554fcab0a5a7d6f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h370167ebf0fc22fc7c25c8bc69c243de8861195ce30a60756;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6b23ea9e3f0eb223a90f08e272e6587d0036169e1fd3d6cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25c4d8e69b826ea1b638436e607df79ab5f932a60ecce5da0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70fa07eaa1a8b70d29971caf72178d1864f13c2e8bbc6a170;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h675f13ea53dc67c7cf333db76933e8e070d73bb0eb0a8d44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4914e71f1f5267d256c3d6e0a88b27f3ba380d206bbb91831;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb18f0cd1a97cae0d7c2677c7c8f6a0fa49c9e7d7d7ab6d39e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2827cb0dc67dd6ba0f138e77a00eea5e9e85257a977877cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd50104fb0d55b2d4b910e1f0c20ea23aa96f60c191d1377d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62375092247fff5a8e3812c5005afb765f28d2a442bdfeb17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12c7a6eaf8104ea46bb3c4777ffce9cddfd94ff8ae55f825c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h552bf48f849d8a9c1c3d42686a3af2e3d0426e978aa828dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4956528e437ca5f72e4bb0a2d34e7ef666250c5c7066829ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bf5d7d62acf5aa58f3e463055c7aacb26ec4014aa6a4eb6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6923183df805b4f0bdd30c3ac62085893b23917ce3f507a16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31919fddfb7cf3c94f49087e160db7e3311b507b201214337;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h794ab08618a52fe23f379ecb5056c38cd76fbbbcc2bb59d43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5547a868d083af1d5f76947742014807cda8365918105ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc7dff8df7f7e38e0a6a9220b9438cac8e73807563fbb887d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f5a12871ee6992d4f02f53dd9f3f6ca0c3aebdeac9070df2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h304624f67221862216632712a504072280dd61a0dcf62d017;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h932db95455e27ee31f46ce6b5e85ada4765d4f90fe81ee0d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc05679d0bae23c04ea8453427f061a72c67a910cf0ef07d24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he08eec7d18e8dc485ac24aa23a9d3caf6f08f7903b303ac3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h607dbc8313ee5eb5c4bdd718cbf166168b89e3ba4ed5a44ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he06dd2b8643e440df9aa231860734ed870c43f5dd55b34b55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd3eb4666dbacaed8a99b3c24fb30b46b377754a9becdb5cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha74f71cd2caf23e6e3ed1b23f6c6ee4a6901106a9e01af9df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2281148debbb119eb790094879553558333d3683678a7cfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b69c272ac442527dc015d687667128dab2fc6bf0ad172ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8250291fd7ec13a8cec93e2599ff676d98835a9500fa80093;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha264c2832d806465083ddc4ac3a8fb800fb93285aab142dad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h787d8ad2c75235bd01ac2560a94009c980692d163a77fc13e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had1785a8cf9aec2cd2263842cd547998dd7e5267e42a74c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f7f0b4d19886d6d098d525a7b88018b40bd45b7203a7906b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fdb08564de823b4d4d1b64271a2d4f5167a96fb634f887fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h519834dbb3406378b4646bc6a3768495cdfeed065f5ebd231;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0a27caac1562df36e1d39210aad591b3d2ec5a809b3274b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h596b060e95951629134bbb3edcae5d91f9c1e00a8c6968f52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d70ee759c5f71728b6b11b0eb0c3e058c36c3ffbffed065;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62f0daf01f900f1526585ec9475b9f7bbeced668332dc60e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6c7d34d2540fc2741b087a60ffa750b7f40dd53d3fdbc9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e0c4d69576f35454036d250baeaeeb5aca97d33ae2c2f5ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99e0cf8efbcba899aaba325c6050eed0c5a827235dd4976d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9262bd0ade588e51bbbc4a214ff51fb68d1d2dd5e0ca290b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb26f68fc455b12b77bf2ca0383c48318d818a21edde6acbe3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75cde5ba7887fe36df741bc3ca8c70f37e5ae300eafd6c753;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbff66b4f63d81c477c7c370c8b5606508eace609a71b67a11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h151eee359307a7ce3a9bccda170b168ca0694ddec213a762d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b9ad62d481b1a0fd8f4c85fd60640e08e44f8a62147337ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ca07763bbe46a41ae38de531a65b3b73d6b7ddf078a1d39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ca7bc8734932f7b78dbff48046a3dc504f47777cdbb799e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9545dd647d5b8698730134dca359efa6dd36187d3e02a45e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2f214b6fc63063c998d882c2a8b152484a24160ad422e8b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2e6a6b74b9b6d8c77a4dc9d6f9bd40bad9514276643ca42f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37b87f6b9edb6d7e33c28da9afda474f662d60435aff923cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b7820dd1db79a4b91111e4d4c7ba9030c73bc55decdf6b4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c4c17a3aa2c0d92669d952ce4ddee7a349fdad13d3ef37a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc3d01ad8db03ff97b8c134b0429fe5d703c508d48a8c310f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7cb0740c5a76b3c1147a90c83b78628a365c96dc5082895b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfa384160420b02fe65d48294778c005499ef8a3dcdecdff2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c525679d2428b6fa182d99ee0e14a446a6692b6c013f9e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8a17b141c3633f10301d850ea65ef27ed70fb49a05542efb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78048e371b750472a5d022b13496adcc031f890f70ea54aac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c47738b614a55fe48071c8d1aac191080c3d60733761be5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a51e1a45175a9cdfba0aeeeb70bc9d006724285897d6a46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82c5b2e7b43ff1136872de5ec4b9605b429a3e2474798ff2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90183cb96aba560b0e79e49ba856dc79f028e0a0570acc0eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7aefd8c731bc1cbb0fbc63802100da329771c3cd25fec8e5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8c91c2fbb28daf5d086faa99297c03626a6fd0553adb461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53a1530976c6e6919adbb08252b3bbc3c4aab3bbf90158b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8af61e2b326863aed2560c443a13234728e3c1df7e2f41047;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfb62cff3f2085f760029ab6200083d2534c9cf7cc6c4285;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5062987e05bb5fc022d9b1f00adb33cbe1114ebd418f9e7a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a0573c218899218f02a69babb9425960b6b48b382d7aa9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5530b9c32322a346fc36fdefafe2938d36a6687bd1d615b37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha38bd4e2595b42b529eb17fe39218f0271f6556b81f496016;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h659732b0ac6e08d474785bba7156f282ef98c89f45d5d5b82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bfb33431147ab8ccae66409942f4deb8e57bd299b455be54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf368c57f81741b6f41dac9104767a8320c1309e2780924cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25373689114a5d6755fd13c8730e2ba8295ca0dbcd16f6794;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3c2130b448a653d6fa377cd4ed2dbda6047548b551b00be6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc76fdc85abef7ac5140c39ad97c3f227e1ef1fe337843b88d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5631eefd3c5e8aa117eee8eafbacedb0343918ece20636cee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42bf10cf4f3d5307f0d1f110d6f004a8e045c08152e6128b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbf52126279a23423aaa8a8268bef800b9f0c7e43af763230;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dc194217876b329df69ca57639e3ea94f68dd2f673874d94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee7bbd84030b95d92f75932936ad7c4d41e625b5adcbc2a04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96cd6c80e17c7071d027a07ae3f0d6dc9d7328595787f05fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc52d4c4f5baf117bf87ebe72ced3dfad646cee29a3dddddef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b1a2d4e803d6a38fa55113b25ee0084260f76459f31d298e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50278271f3e55f1968ff8f47de7395925fe0b1dced765aa87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf027d5e90687afc2ceb33ed91a3e02aea312235e651d95247;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4124607310e313b9d4bf8cccce89fb248d46605218d88291b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h767b0cd87142b32d6e5bf4c6f02bfcb66f0c7ac2639f22e7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebf640784166c1e2b7c555b7ab604baa605136276c5bf8a61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda659eeab5ac7d85f5959a3479aa577b37828a02f1cb61e04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c74c635f948f23d03961efa00f7218b0dd53bac996b43f38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23d9841d2fc07dc7974bc7a7f279601aaaab546ec74fab51d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60933a94b3580d27c3b718dd37da1143db5bb3b2e73362308;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae85c37bed9125554bf4c5413b1f6f464a20f83e34bbee09a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ecf17710512ddcbe831308a719b1d04c0efa1c994a53d656;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf96d6f83ad0a8566898108c9513d79f65c6742b3438cde98f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4323670cc6080499ed34504cff9d0626d153514e15e6fa4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a690a5e1ef4de9fbcbe319d77627d85c9fb214e2aa309888;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9abf91e676c821da44631e71e0c99c9f9ac94326ae9d4cad4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h434519c763c51be89c0acaba8efde365339852fed9ac5b0fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c4910039f1e51c0a1efe48d78067c0a631b34281b40102b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h210d62b51d6eaec268d62a0dd38b6d4beaae6face629f01a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha17008cc333b35886763a3694fe8daee4a3f93fbe2ba8591c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9834743d0dcb0e22455c444424aa0c0c6391e4b1643b5b08e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f2c666fbc487bcc4d809bdadd52295d8f9fc9cefacc5a610;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c8476e9689bbc346534e284b80e0c79fdab7bed071519a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h930ef7f2c8c28561493ef276b5f18879c94cf1252fcbcb671;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h237f9789a1ffff469b8f6f80712235aca8515aa53fd13b64d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefeb012baca606b11f4a9f576099549ab14ec4c62772242c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha03aba0bc7f44dc415b6d214810d718e1e45d6fa3349e6464;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd34b7f0356ac8fa6f2ba5ac1c00f9bdb64ad7bc05c112e299;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5178d3663be0e897d275b1bc51745b0da3fe00998a5f495f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca971126a47716149d5db96080bd504edb60ba5e87a7241f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had03add8949b3e8e6c9325b610748fb373218cd355f341ad0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68e0c436e2f61a325f5c0c3b45eba5360542ec2fa1455afcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4fa8a304619113293e0cd82f49b66e231fe6843be5e25b0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32e72bae289146167533812824cae29966631cfe43670f468;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa2490126ae5925f029333c669d4b4206cd25dd59b6fdc887;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ff34d57d6a1f369598f828827b81ab2a80090591c0f07513;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha91059625c008cebc30e71152cc0debd9da80c86436cca8b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h874fbcd714eab3b3eb609dbb072ac5bbc046960a66b20eb26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbabead03b004d756d25fe4755eb791c8efcc24b6e0cdcc84d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdf9265c6bce784ec84b8f1d11713344f6cb3b89043c9b38b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2aa7c62833f408949c7eb6f798e553994a8a253611c88db7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb80b2235c8360871aae92fbe3b54923af0cfce6d5cf2dc20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h305d68b9f65327b107f53c9dbcce918044a8c935a4a588b5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73a1be8808e8127c037b19496d2d612a3819b2ffc3358e5ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e34e83a4f661a16fbe3cdfb0b6cbd4095504e6a68f2e1a34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heffdcb7313a3c8d5bace2ca9a89bb4611265fb8fd9421a7b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb6abef0ceece2653acd798651d5bdb041634fb3024e65201;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17b4a650fd1f1e799daa624be8334b10756bf4159e6fe4058;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbfe367dbb32dc50046fc18723b142eeb0cf8c6c060bf821f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b029fd1d1d4d1684da3473f28f0455de7827345738bbd6e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb80880b615eda5a45571bee4ac8c3820870921e7aa1fda52c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ee85c0ff5214449ed1ebe9fcd96e088c9561c7338637471c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f5ff3bd172b6058f21f6a5bc26b053bc5b3a0c2df2bd767f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fc107ca5202daa983c1ac54e6952134eafa13e86b3f5bbc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a494e2c97df74645fa258e960c53a99d11dbd9e28a8012a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefca28c7a8e49ee1882c3b441c8768f8897adbbbe36f7364b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d7c93ca5c6ce644ce54d7668703b9c965d0656eeaba3a80f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38d6865b363b28f0d227c82f8c8f09ee9bc8bbbde9304dfd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa783f077f97d84c6b2713fc8d27eddfd34c3e53ea0afd624;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb00b0fe32b9a0b2ffa5882849499a801d0f65375918f10ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd273b014d2240b0d00f54766e8a9537a5c1385508721d5a3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ff34de0cc1c71b7b5cc17ad9a9cee6c48e11b80e093f3e9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf947071428e786b330471d87495e8d8984c6132d4059e60c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89fd9062dcbde92fff591f6e2558dd45ebb17f30284fd0a39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b8685ecd40a0d08bad1a3dbcb8cd2e16ccc5d48f29db7d7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe0f2c201c023f740f4e52aace3fe85755bf69ebcd914b452;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66acd47affae82ac20668d0e19ad242f3fd6abd5d2967e01d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c42c9f446390d44d9254185c76c7273eb4d41820615f5d55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf734bf1e89bc3e65af9fa4825f6e857eede78ec6960429cde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d0f81880c18e5a7d7419fbe2058bb976311388aee3512388;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6964db4a76f17011ca77acaa54f80981b80ab076cafd20225;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heafb8e88d68f93ada86c5279ec1c8a31ab3631777f40671ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95dfdab8cfc1a5ab47180b83c9fa7de53085c494deba0bda4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15d816f99b5d9ad3b4730b6b5697364eed5da026fc306876b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1966cce81fa42e725272cb78c0670e241c01207fd7452da0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h906aeeac3b674a2036af939842734b9599917f6e5f3b31b9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dead4fcc9a927278c63be674ea6a463196555cc095858d4d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd109d9ec71785f2a99a49efa6b6d51c5964b578d05ad2213;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb56546b9fb05d1da611be0c07cd8bcc779e7f3d502d957c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f2a7e35fed44d6ffd82db1c86594a12efc637db84f9dfb3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c2f88f0a95e87664c708479ba61ca2ecb1b709cab4a78a44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d783e8177da51aad6637929560c77f17835c181702daff52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha72a84b056a301def727a7609efb930206be6bd0393f009b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc89f969bba68c72feab43dba1bded4921db7b60a8c9431689;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd64fdff44c17231d254f2efe7cf4f5620962c63323824db01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf08747b65c9eb8f0ca4fb459bcbc370e2e0c3f7c3365c5f94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bcdd6436aa34a01617577b7635f10f3571f33b44bf0a9df5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa4682592f823a6e9524c134950e97419246bea4a601eac95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82f6656a412cb718600537aa33db361ec1ac07e997572b13c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8608ec64b74b26e66f0cf96ae285c8ef575a4dd57513c3fc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h521781c5bb82332a6c794604b4ef5adc3de839e7a37f8e753;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93f8b1cfe891758386a65b3d7da5e2f0a0ee87bc851eb75ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b0621016ac32ec15f552b3dd283e661becdc7206b9af8d92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf97d037345e8f77b49c9afd35f54f0c1af8bd9c3a33a254fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1df9225781b65d5213be4e080c6abd0dda1edec86bcea3059;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2aa754dc806e4704ad2ae3b0c25821b8bed48ea71d8394699;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb0fcffcd04931a7f0e1fb347cfa298a2eafb00c2a40b941;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec2cd179ae90011e06069e88aebb10d6f41039f26264cff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h807952e098eeb2636b8871d70902fcb7009df21ba1c17aaa4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9c2a918275946b1ace0383232e5ec3f6db279beea3fa55e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b281f0224ff9e16340b4a1ffa4e07886b2638760761615ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1978aa9a2540e3da1ababfb0feb72e92de5814617b6f8fbbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a6c870df08ce528201977f9153576ad6807282c4df191601;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h969983f12ef7d4dadfa0895728b23f84e7a97b90f80df3d97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce74e0434c2e578ad5835503c956721c92b96be97b37b2e67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71129d3e5c9c913229e3b1966189ef696b755cb44492011a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b02dafb7a1288ba3cbe811b01566783cedf66d0bcce6839f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he114855db0a735049ed4fcde2bd93e9d7a4c626488fce0adf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a96b731650ef5c21dbb65d331fef243606bb297661c4819f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9542cbce4845543b59f36577d26647944c3749124f7432b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e87fd31cb57dd7ca5867ae23b35a419aca9c55cc21b885e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h444ef65376405737fd6314b3ffcd2b6f9b8ed436db285c811;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59adf1f6a6a84ae1bf041edeac34b619d2b670c4a78954031;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3afa9a743748e6e515179a862c6325c6e411825e2a4dcb43f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24e30d2b2622034e4cd363f94f028d2117c398b4cd193284f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa4587455b6405ebff8332cf4484e6127dc0be7503cde3ed6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc961c5cf773fb66a45b8186044e43d210baa29e239689525b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b4a2d275fc4e0b2db30f6530361ed3fc934d4cd3af48ec52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78cc22cf9c4a7782979e0197e0a2a44e0a1ae6f8aefb006cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74c7b3f83514162efcd6811ac3a783eafa709dbf55b28a1dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14c805bba6cc71e1febb0778636b07e97ad254bcef3c38050;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf43b07e164a9c9baeca242afb9d12b7f53fcc5b4a0f638611;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha584d6bc4b881a3a8da208ac0edccb2319548eaf44b770288;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccb6f13fbb7f89bc145d9e27ff5398317171f5d68e355e483;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9cd51620c8c048ca2c092de1e0d2e44c00ada607a561ac01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he18ea6000d1482f7c96e3f370def6aa082eaaf9984bcc5924;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0171265082b793a9fe33bd802181a99d37424f73d0c266d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27dfe2d074dc79f7b0aaf3f0104d23f000349e15f8d08f2b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcb72653ac6e85fd56b0e6f115302b75a23f1857ba5f22e36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h679fd873f6d51761ed7d12c04ed5cd673205cffe9bd5bc925;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf043a20e87d71ea596b346f4b36c497d5a28b8b17daac6f5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e9eae0d0484b0e5e9a736b785d59847f463de4d97842b91b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72fbe8b265753719480e7f49cfeada7136eeda54327a193e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10615ff28701b72f2356af76c2c447c68050cbb971036cbc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10881df0d637b9a1b2245d7443b29a907f696e90d2a8a5c37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38cd975d5d965e57c7ce9958c097cf46c4b48e75ad1a1a1c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bcdb99b0386edeff04fe06b38ece9e9f3cfa1ef029dd8f3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf520d5aa349aeb0b23823f1e9a3777da7e2dc79b5f86ac868;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd52de91f22848e7f7dede4731b9edf62b466009b8bf2efe1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d0a153ba83ac5af02422d66fa372d87c5e50cbe519f9078d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf578757a0fe203e3d036b0c53204c9ad518789fd5642ff242;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39ffa4a3dd6b324279c36922c320a6e799fe00f01c03ca9cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h918791aab138da8589dbd10984605225a7ec818b59d0568a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebef38838eba834925545619f9b3373b8ea172b268dc0dfbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92c14bb27dd55b871d2d46d290d7130218165e952f9ae437e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h705cdc0fb06c9a733925dd0b21a00ec18aa55584a11c10a46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8172f9ba5b43391f346bfe33966ab4f50566c91d2c11aa534;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf173faa0a2dff558973186110291f09978f862d75bb864af4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee8fcbb6998ea9634a6ee2d3a7767a5a22a10a7237e1e9405;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2019544d3e139fe0c7e3e920d2e3fac1ae1271fdec3d1f727;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb282413c29e44a3dd7df9fa4ec1f7bcff56b9ef28f00f1a25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0f4f566d99375799c96d6a5996b903ceeb68d4ccd30bd805;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha075b5c3ec44bed0397d37bdf4b5aa3472de2ef339a4e2f83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9abbcdd292a484117f25a31a665ef4e50a813cfa10ab6a7ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab4689b2f8ad1460dca10f7b6d1b0381b2d7ec453bcb2f9e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d8798b561a62dfb41b0874ca5644eb8cf89c03ad990c47e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd88bad5434cab43c965c548778aa2118602fa947922de81e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf359175f936b42b5e9885e222a5d4d73cc276185b3457f7b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fb712aa02ebee2067e1d33d574713445f7e8bf738b8d5c16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9b903e619e97c68810b8bed8c290d5dd340171aa6738acf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb32e80130153b0144f55092ed281bbc5255aee22b0387b9ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f44ab1fdb729d962c192ddbde763c3908fdd152f497abf8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec6a5c74cf679cc34f2c1d29f99350eb5ab98872dbfe8a876;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f87a4fda873efe10252572c47ca9408faf42c7810c585132;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c3fce38b786886d26a61488cf3790d0954eda9c98e5974bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f2f80282127734e0d598da890cce2d7f62561f3fd35085e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77c7e5768488d60c77cc90e7115959e2074575b5064ac71b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dabcf3b2c7136501d2ab0cd38dcf3ca3d6145a5a6809ae03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h547e38675217f66d3e5fbc46c06d2a2834fb35513c109fe2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea9473832a79ca7875a13f8412917fdf1a1ca35d172e1404f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h460ed8c474b6dae001c9fa0299c9d2654fe6fa3ff69d0d404;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c28f48a35ac309363aec63a462a52d4f5d3e7b6dbf0d5dc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8825bd06cf301827fdebaf73c04d8d74d39eeacf09f30b7d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7894fe1de690fdcdd1f74a24cdc0b373e6355d9117bb4171d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2140ee86ab38187b055c55f0658d9a1cdf257d7d29dd4f409;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6d0e4f95063e4070fd3a31f1352548c5d78542880725fe4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafeae9b37331d8df1dbc4bb45fbfd9fe122132f656286efc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12d4fb38fb5c2f27dfc44ab31e1df8b593422dc359cce9738;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79cc729177cbbf9e40f2411c8b63ed0c1fa1f05388499c8e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ad5e8479ee33932c52d52993c55771fef11e27b5e0d9e294;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41a223fd526d165370fe46c4fb8f273f0de01dba11127837c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h685e4cb9e7646e19a1c1734277beacb99770e1b937747134e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e4751f4ec4728474b1a2f7a27ff824a30481c7d7fc84cdec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha42702cbbb19b216e1dfb52abfc552fd71089307db06eb601;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee0e0b7f71b92c0e7df06092640ec1aba63863e4ae371f12b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ba393ce45dff4947360c9c0c71f3069f876f9701747f29b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h598088238e75be858c13b9de2f403e236731dd01ed6d046ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h738e4518b778ff6160d6ca4928171e13f76029e35cc4915e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88976bb74d8ec018043ab4637d9aff0ca5789b2bc63fb934a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53b4720ac154ba7b7565f6499c059ac6232084fed65ccccd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe676b599768e102cb820b7a94063401d7c118d1fefe69a5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11243b1b2aecd41d8390aaf1460ca174bd71cc39d70c26a44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0f8f2857be04d2e4bc8add825f1159a6b93444b88be5886d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dd890623889ba434bd0f05df685aca6d9833c7cb91d620e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc760fd6c9c1d4bf206af8c270cee8dbeb36193c2c064f3050;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1434cd33b20cca43e2edf5d147ab1d013bcd9a281e2b2d19a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haccb7556cf1b2032e46624a7d4be334e82e13a84284aae3df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57ca08e720a309e39e890e21501b26edc3227ca957989aaba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f22545ae239130368d8a1c7830e40a3f4d4e1a32cf966aa1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h240dc9fb6e1494a99481d2ba86e9e24fd225fbd23608f01d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6133c16e2330667add5f2d015f2b4ac4facdb305ace568e7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc474259dcbc8f0e8ed339951ce05aecc80a9ac1d3277623b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17826fbd1711609a6495091932056241dfcffe2b565be411b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99fe88e357f7e85e59fa8eecd5a95333fbd62652f65b96a83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6fe2d807d0c73085c77beb71b6b211678f152ea1e38a782a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d252a14d75fa8d99e9753530f47a0ea4364051246a7e51ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75667da7ad00638d644b79116424185da161b51b0912f0407;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbde14d6e4f7b1c9fe3e78afd48d2d46d0bea3a31909f17318;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce114df77bb23b839334ded86f1d02435f77e203c5e38740b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa09154976d4b128b4666c2f1565662c456deab80833e29c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc7b112bbffefdce53f3363e30a43f74609e12cc8c3a5f8cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f3affd1e776b7b2a91c71cac56ba52a8a7903384677782ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h826892cb14b36700673f28cf83da9b9178fc81e4bda843fb9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha77c449bb50282cbe8a560d5cf2d20741b906d078453e3dab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4c389d34325ce13ad87b44ebe6cbf04c442a328684ecd4ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd729eca0e6c6212c0c3d0889fad281d2072a8d9b58ad832e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bb0f173bb1e14fa21d720c5176528d4ba1c352483eb3d51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb91281ba69d3bac87a6ed75f41cbd22bd51d1615f14d571b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e0b5c0183f00345cf93ca73b7ecc5940675b43d976504785;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf56d1949d539ffb97075a606c4c3a49118f2a924c072e4c2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc60260daaf25432daef7d845565affdbe113992772c217e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd2b9049df8c535ff1b0080269ceb90359fbe1f7d5435546c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4e2975d4fda2dd730360da1ede4fedacc0068a666ac61394;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6cdaa61fb14a664a5463a2607b846445fe0255825ebbabda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d089de49c395d493a8105084b278c9caf87ff88005ab2745;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26202ea51d65eefeab25c0012522f699af57445878088ee0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he955118b41a43b8e18df3c1c1def72092f694515483684be1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65228a71849103ab850fac2949e27ec649c9c7636dcc1f90b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94239c198805747867956538abc72187228da2ede7b388dbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46ae30b3f3e13b89f969726c9bbc3756ebbe9851da3137d68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1060b2d1b49113d3f98de7fa2e59e49de91ee333948e1fc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98ba8af0edbabc9a43a6198cd630e7149824f3f7d10bdc3e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18bba005d487eb9a056d2be3e097d7bb6b77dc3f28ec6e731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h879277157e8dae3d909eb0ef27789df5d16dbed91f511f1e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2713207dd23cfeb636a4b81c628248a51919564a429fd1e24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fba19cdd755fd9a662e5fb5fdd4da06d3455e2a0b9532ab2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9f1e28ab00b012a2b85aa9778d5acc32b61bb40cdf0294e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa50479ef626efd832091d29465c5f5914600feb39f3b41d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63f789e4363705a2ae049f49f017b98fb5d926099e1fe9878;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54db6c6cdd0d32eb027098e4c529fc10e689f63f4b0e1d2b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8b2b341dbdcb00f68f298bfdfa69b3076213e5eae0c7cd33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62bad0ac75c0a0d2e2a679e4545b03590f9c4f282345348c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6843601185809546aad2cabc1e2ff0297b9f889741ffc1bf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he391de0acba7aa619bb9691fe5df15d95919f66869aee4816;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc21ff1d3b0fb68274eb958dd7e1311aff945b2f83e7234091;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b1de936f08dd5434b172a2edff43e168890abb76d353a326;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95f4e6a66ef788d799c96d02d78a44dc5976a60215eaeaa6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h932c40fdd1757039221291e7aa3db5ecaabd0365011ba834b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cf708134563f1132567da4a4f4837eb62529445131bf76af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3454f8ee011b3daf46717943b73d0978bead9483a8fe42d6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc3c054e5df025a968c31e765c9d85e8f1e054be823d6fc73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24a0170723fe978ffb2b9073ec6344ac636f67793232cb652;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58c0c4307c0b9c900b1e5c20ca719a64a53429e667f3834ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f595536a4615c311f866feea69084ff1947a57f10a168134;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c922decef256dcf11e7af8bd53f345fd32384a231798d75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64cc217817db623922588aa73e93f4f44c342485eece28b1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67b5b1c5898876eb16509c81e7f45a4d31abe5754838d96f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7dcf383e60a51d47b990a42cf6d6ffb690f6a084cd2dc590;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3905af7d0c8fcdfc99270699583094bbde78b2d2789ac0d0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h660e98b4d73cce8890f382c43063e5cdb5cbd8c604f6fb33a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cc8d949fde8797649d7d02b29bc8e4686b0535fab70b8f11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h964d93573ffa8569bb0bac4431b5f03109c23dd5b49c9ef4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h229baab45c7edf4731e8694a64fe51d26a61907d5a080fc07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89fc6d546591abf2cb191d6876eaf5c897404981de8a17da4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21bcb1dde8abee15024bb9b637cf8cb931ba2bef098802bda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h122d433743ed8c8ca9c2f4b0f27be9c84448a3579e8160412;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ca64dddce933d0d1b25499829e2b05e5aae6766f05a5e6f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7316b9b65db91da6a25eb34ae648966c1d24db6a9af844a97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3b99836fc1cc9a0222e34694142643f9aacbb264b650b556;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8dbc3aba67ceb1b3d4f653d99e531d912887bf576de0c3f26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had8a22e0b9b5ddb6e7fe7b8df85a9780f9dd9d41abb023611;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h938449b3cc2da1002ca8e4d6d15c7592258798d75830e1322;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a12ac81f8ac4a032453d8e704175d30cbd7ad4e9c3c44cfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8adaf105c609fe7db82385b278be940b96ee5b8ed89d1ae2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d8b39af24ef9e543471f1428485680422660bbbe5de92f36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41e681441796744b2f549b18541284b1027b3a23d132d8c02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec5ad95eb68f002814e3043761cd04217a1e2fc15e04b48a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h910dc1771a9e11c345da423429937583e8a2c0069256cac5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf06a8fa7fc72c0f8de7b505bba143fcfb3909ae6c2dd31739;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h489ad3fcd5dedde156c9f476a39e4640c7e5bc14e84006a19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49c88f377c3bf19b3d1ce54784fb259e94728658fc9b15c89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a9f3a2887bfe98602a9c4cb3ac71491cec516ecb7b6b4fb4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fa0a4aefe935369261b2a12d0b5c6b66af2cfb43b840ee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7dc93669f7dcef8cd915858a94e44394adbe42f5e62a5407;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89043a42f0755c15e2295c8a37b5d183b65155228112a0135;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51c304894929fc50b667c9129406ec1ddcfce51aa12e3251a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc3540a2036eb1d4d5c3c4fd83d2db6173235820bec45e7a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5cf520fa193ea82cc04e4fb82dcad3aa3908ab6422e66b6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13fed5afb5b303c53357542d89c53a0373c1e6d9d7fd935a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ecfbae11b67958defcdbf66bb6009ac73d039348730f55ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8ba748cee7fafeff22cc91fa86f565a5a788336dcdd00661;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f57ec318b1db09d05afc80fcd2995c08dcecd79001dfd7ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha49ba501936668c722465ba5f1ce7afeb966d2231153ddc50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44e2b8c0e27118446da4633d0853876c8fcbaeeb8e51aeecd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40d29958442c9f262b53923dc5603a1f905c3b78f0cd86f25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he75ec4ecd090fcc2ea5002904d801276c9d537cee352db1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1a3fab00ef489f977433c40f3bb27686922975fda993d1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e057655aa5e1eb5fee1e5a5fd2e5e39599ada5b953c7865c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24b305fcad4d3641714188d5f278d7692cccdb589be33b0a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ff99841c09ff04df705d2036c804fcbff3d97f05d757f14d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b6bfd1fe1580e92245859d2d91ce64da9b6cda70738789;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88181126d5d58c1bb89e8fe87f49678f622b03e0e39f17c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacd95e51f03d8df7ef0dae8431c0c13ca735cc86db212a35b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89a43b3764c27391c3ac2cbfdbbe42948db88f74a3da2da36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca725a7141359c145852e47e9bc967f78bf73dbcd681f048;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53554e23a385c7262d5812b4c527ed0e30900a41f838d0a2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4849d309edec3ae460f5c08cfe1e433ecf78b6dff700ac982;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha93f6dad2f4ee1bb3dd711c7ffc7c40aa1bee12a86bcd6156;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10ed1cc9945dfd956470dbeab8d7711349018c6a1f068cb97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd123b1facd1a512957f23f6b6cb3e48572677de26b18f7e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e38954a63de734ecf44ec92343e41698d4f731a313784744;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdcc60fd2b050a057ef40efd38210a0dd9fc5882f73c896e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70e6fcdbac4752ad37db6abc92ae8c72413241f15ac3937c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he14bc18b4b0d4fcb26c307e822880a15972d49eb9bc591b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a6f8589ee5fe4136a081c0ccc83c676e18a964d89a48394d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b0a0f229586b3f2d74c8de5bb45491f7ebcc840ae131db3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6b42ddbb04edd9d64f986387b337053cef5819f8fe661987;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1ac9b9bdb0807ef6e58f4ff39cf50f6e060119694f800dec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fa96162547869ca3025dc7dfca733e748d97300dbb5f4547;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40355474b595f8a350587734a79f508c50ae5576bf2440089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h885b5ea11c7b2b0be94c8ac030e42540cd85aea791b17ea16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dc0262955f7df7efa4e76a813840dd38662e1b2a37d019a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14cbfd47e5d42dc5a4c61f541feb21dc14d2c2357b52f87db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb175a5e5dc9f3144ca33b498f6271b12569d8dc6199d7ace0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e2a3bc4209e94208b1f301fc08384628eb7a39e57b2498a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9373b41b49eec4f30a2ded543308adf7b2cd218e902c774ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b962afe60fb5bda32741421640da334aa6781966464b1caf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18cabc3a849d02f2485ed99b41502bc4580924a91c2abc1f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e327e2d3f7debc9e32db767e3bb8021d24be063620515697;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29d38dccc89bdfd1b1e7a1ae64a7dd0de78008692a89604a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb4bd4a251c4015f9dc0422743ff1c7a0fcbd5d4e0de17921;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7595368b3d8dbd1577037d67efe0432c6133a5f88c90d6e74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h993e588386aa9d63cb01eeef385b289a799637b1e2e5cc6f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd74c69db84317d4572b9217d744eb51f0a40a2406e94b6da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf132ae55788f9461dc0182fde398d827eddfd1a9364076c12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e8fcf355cdd11874b8b1ad41dc32c9f28a64730eb0adf5f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6dcf4cd5b15db0ca01e9004b66be50858a1c83da792a61b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbf4f6e7c8eeee204c407b6830b4a6a864833946279864b23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccbc4feb32e4b66c22c0568448a867f12120c393598f170fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd596e4450eb8a8554ff509159b58a644d0d7cbc1788dad328;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4419a9d0126ccf3032457a4def2ac32cbde82efa67fbdbc9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8d9033cc4447547ee519f88419c1a8c61229028ec79f8a80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf24ee1fbfc430f7f380d7d6ad7a89ddbb592c4db80597cfc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e3bc7f7a7ec1fb858f498ac9812829a4a5eca5ea808e922;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4821d53d424490ca100fd69abaefb0fcb39202fbb5f33d8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa0e3b7f6dc64c668c8b067c0df7bb33df5b92052079d9ba5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bfdc26860f0708413637c3eb6c52cf70aaeaae0bd78e3f39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h271362b08b0c5e8e843d5ed51a6fb1f59dc090e7d9987f2a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3988a9fcd3b0cb4a1c803d781a8cea72a8f3a498a1d152560;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d0c7fc6f9a0f1b2cfb7d1d14e9b3375bab945a87031920e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd92fc240aa7710ede228ae90762867eb845b3834f8bbf3739;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8982bf7ae2ca81eb1d8ce6d404e6f85f8e6abaa118d0c01ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4d2e956ebac488416f6c2482ba23d6b16725572ea6b4f10b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h909f0818a7433c13283e5f245634463d5174494ecae7fe3ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h422c3c7a8d1b9e73339251907fde9e95a495e49f9af06410a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24383c9e02afa786318426ea6631a9e55fd35570b4a68e893;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7406778aba2a8af4aa50aa3bb3a08b27d89fd5fa2ffe252e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9be10f3f33bd2e746cfd1528196c4d65a3cb0c2d6ea4cc297;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92c9c22a97988d38150b58539d6f9975fbb3ed15f35b19809;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1065bbe7dd3331933e3532ecd08c26d7bb1e5b1f67d182923;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf012aa7595512dbcc88496fa5e7140b685f8e9ee7bcb8c222;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f1e8dc0c624dcfe64726f0188fefbaa24e3a12a9ac30c2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ed64b9206620d9895908adf9c18633589cf5669abc48c46f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb8769cac5fbc39a728bb523d9f5fb84f0727dc6ee9c7b90b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb416abcb22be0654d9f5fb2d2df81e7d4111dcba7954ed12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6ee8255b4ff80df7551da52442abda0488294d5635c1d7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49a2ddd005614e19f809db4b56b8b92d99a50c2232cc3922;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he538513c62c1ccec937dcfc6acb709264a5d7a9d1ba74dfe0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50014e3f8dda47c97cb5a25ddf0c711e14828b95cc3608e4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc2b49bc148887628a8e2e224dbf6f277eb0c6e3a568de4ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4397eb44b35ea4209f1b99c5cd91da8e898496572f4f2ef4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbff367fca7db703f5b24af70a07606a0a1a6c1bf18bf88e89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h502853c3d71923ccc5a4bee8cb1578cf3208b08f9ac4792f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5635c7286758c7a844c37019ee97b5a34aedc3790525e5c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2284845bc646643387f06ed5d20b7327275e62b8053091d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a3fedee8f201f9518b53e5a448c377d7e7253b89e5a54dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac5a4d964058d57318cf5ff70de6b31b049a2fb0b854eb363;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b25971590b11045266729a6cdc17b44ea1c2fa15e9bedd06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf0f7a727be49b56ec6e2ec3104cfb8aa4c927e4fe3c61898;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31585866607d86d408d30002864ec4e5900de37c7506cebef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2ba30ebab7f3599cd54479cdd8501481f0c9492f4b1378ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75a514b5f5c8e018afb2f11e9e8ef0bb272c86e6c849457d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h783937530a2c36239018a149eb499c7e538e7ce558af4242;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h689128b9503b62f26280b824f3c6b6db0d2214eb582df52ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e92aa375ec6820a4ded9c276ec6082adb017b425085ca37c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57c1559e5e560b0fce4f263ed79b52a2faade6527e53225ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d4a674b931296f9fd31f47fc5c59f9b6f9e861ab8c99908e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he022972b03f4b070513d193e8adc13fff25e3ee46482773be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93662011db5ac95abc7acfd9b2fdc5a58a28a9fe7eb1c2f0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b25c7fee2cc584d6a8778e23a1576295128b072f1cb64a25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h476bdc5775e9cb12f632d12aeaf97de66d2baee6cd1c0d65a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h540fac289418479f21428a3dc09ea957f561d5e9f7e2a11f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd304ac5f50a131ef0cb1d0d0329cba03b7bf922bc9ae4aa16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2fd5102778d915e5dc7c0e1ae060a8289fd70182f9bf6098;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h273c37b9729270b01989017d0e8ac54c5bb8bddecedd569a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf82be83be645e9609673d74fe521ff46e3c256aed5347c60d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94df91a108a38f29bec296a6793af5525bbc83f10a573852a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f20554e61b39eec8502949bd5c99653154698afe380a9f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5524a8a67497dd2d74fe2126e86e14e4a6d75f97d588f5813;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee1fa166cdcc61e4f5494e4aaffa41014724e806a0e0e9b8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4541194c558c99bac1e21e4c35a84e2da83de88f47d110424;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75f01ce01f8ba9be1000d16d5b3065e5a85388cd71926e025;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf308bdb10dbfe71b76e7222c67e5a16bd5a4a82087032429;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97863f336512fc266366a28c15649eb42fa4d1f60cb00ce08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h163cee34f80f03af0c4a464eb0123b951ea5cc852fb7160b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3874fa62505a3b0835e4f4f7985a24ce8d8e5e3a5bc741210;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb77d18dd12aa1bf433b434dabb1d6ca19ab0009270bf91d4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5065dc81137db76b065052e27ae8a9817a3389316015c16a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb0bdbb4685b787db27c876c805b0d5ec30a8603752e7f3f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae19f8f17c2076969d3767d9a79279215e76f93e51a81e271;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4198985a441249946030cfe4940c7b6d850275e6d7b37bf9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90745d6e4265ea0dc74b955d515bf0b010766ef344718a5e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h994e1ec788fad1e116b19fab2bce7ff25031ac0eba71a2a76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had4db6a88de1059ba3832e310f329be3092f157ef345aea45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12c69cee2323b5928e342e804d094c371939fe42d1efcad95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h209b51ce1307f63873715daa8a0788a4bc843a65d2d2eeede;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d75c4458631c48afddb47a486f5d970c521b631ba2ae8936;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f6e54adfd82f4c79c1896219baf2a8fbeded2f016fe81e69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95c6f7619cf76d9f6e8f7ce04e54260f9ded57e568def435e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d423ed4306c4c5430174fa7539cd770650a69a73d6cc6b2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6428c3af9d520bef71a3c26c2138aa4068574f61b21ab52ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4833a4cf0c0247bad3d9666a31c62d8405d589b46a0435413;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49fdd218910d3556c8218e7e0d5cef9171b791949b5a79a8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a29ee1ef71f3e5f59a31aaef1439b3ba3f2206d3fd74c739;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a3039e2cb7408ca15cd99a69088ddfd97afff82b1d36356e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8be15556a20e844ed62e0cc853a7330132bc469a66f7e0654;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd87519525c37ba448756e02a3f9fef468b11cd542a57c58c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4431ebe5f8e4f1d01f98d9b7cb9748a35c7fd4f72cf07b445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f206a51fb58dcb1d3be802252ebb2867abb02d44e82cbfb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a9afc48a6c69f71ec34a19575513658ba2dd96e1bf7c508b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48005f8d8c87c68cf4af86719a9137ccf6b4c4460f1df8e6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h460e429cbe6a31e983ef8ea2073ad7dfbc0cbc09985dc9250;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78e57a72c9f8d4c99d38d77beb2a112f4b15c8fd42f81ed5e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ce888f96cc4161267230cb5a8c4b1e3a29fd0c2c200ad44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d90414f49d3975e8004a5f5e4c35fe866557623edc243880;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6098997474ca8eb166f8d84b2ecb395c655a779c6efe819d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h543df86a6ba32c004492eab8a3f914c3ca998f81d250fa13e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f66ed61cf6d182a3a594df9a5220dd6c0ccaa05aad9d37d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbaef73c2df5e18c0022285187ab51f1aaa9b3cb8b314945db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc1595a98cc082ff1b094b63702eb652557e8a6e0fc4d293a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h916aa99b68e48717dc04e7ff12cd9478ebf522a667fb66f02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c02a5acf8b1a3f7da6190e424deeb59d98c54f30fe5cdd54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2b5be30fdc669888512d875d276bba2e42d9e132d51ec1b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd20e131b521080775ac0999f8cb9104f62860435f3ee7f56e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h373c16735413f4c0a41a2d2564da2f49afcf7788305481718;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc0965a339bb581257cc5c01c56ceb0a1ebe700a9494ac953;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13193e5de53abc3e6e8c60f3c131111c4e32a2e556488bbde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63f67b9d3ec8c679fbc4f47d3e34471095f86911241599e55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c880901c56776882ec92a0d935d8f2457799b54e4f2a82a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf617b0b9cda85f95bbe1688d43c13a90d1e7a44088dc5b7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9096684169d441c0512aa23ff388d55fa27507e301daa4697;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b4d410672753979c64da798412092561ba01f77258c4d64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd1d1ce03815d161dc8545af9906f5a539f4b0808342fd94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h199d2bf9af2f473f6fa56e0174ec2c7d6b47a6b39092c9476;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a5b1c875d0ad2e5e9c3a4ce6533ce9d8416dce5acb1b67ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94d261e2bcc706f3c80fbf67cd65c63c49d8a089637718342;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0e4b26f1327084edbab5fddf587bdafbc50a48c23f5d64cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd39bac56ef7fbecb80059f0d3a88b7c94ccbadad47281c964;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h865ed313665cb828d260f0d134d759da588facd180113a71c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b7d7016349bc36385eeee52573eed1b2b02a57b378853aa1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b7f9ea78d43298fee1342017aabc66c02efccb1fc19831f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h345a093b07d167dbc498c5bec49c7987367b949e787cc31c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2453eb341c2919bc131f7abc559b0c040f3cc133293682912;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h345bacb6d182c08203314f0a58d1b64bd2c420e649590563;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9ce846f5f2fa820ca206e4802a915b1ac6f7821b3e980e8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcab6f656e8978bafdb4769897dbf8b05dd35765eae6f87b9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a4517cc631643626a262954c2752e53f2d6e64524005e193;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9781f7a29597aa92bdf2ab884b7d3563aa2176127a6af9958;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e4fd55f7dd9162291fa4068d2d628413f6ecf9fc78386ed2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe9b3f044eef1c945279f3acde1704434b92861ee8b288919;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h936b22a01d489297d852ce88b0880b7d7971680b702f854ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c5f722b6ccbf5b0b0735d0dd44c3a5bdb8558c3b9e8ae65f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb92fdf7a0633647cd35019a05704cec5a9b20b0838946ce25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1eb480981e6ce34402f5b1f1d7b3617002ea1d215a2c9616;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdefd4eb2ef073bf09df55ed3ddcacd19ce0eaacc0041400f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e944ab823f1e79d2fba64260db66ee68dbb393ad4c4f7489;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42aef939074cfd93bfc7acd46844a261893c477b2c29781a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf21e6619f77dda88e7547d18d294f648c882a48db4542f39d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3df367a69b09dca1bd62e4a04f7a2cc82562681fee133bbdd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd079af1ded7abc082bf00d60b004e8da687572ac462986b4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda9f9a212c34ebb723e014a14541f1c406502e2175b0e6a64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda2ba2d0c6def914f1b85a303d6b74713c8d53e5ad438064;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8c685c1f3da8638a8d55ed6fbb8574516052fbab6365d39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4535334bd187c55679a5e916cc6228393004a7bf6de8557;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd89ad3e0884e7715b4d6f2506016641bbeb573b05ccc4c396;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h427d86326f24cd22802b4392f75af16349e6330086737ebd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d4102adf69eea82344b92936f0235f2bc19c01a1c1a9de8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf12e20982a9fe35c8ed9826e1b603cf77ef040dc3a822c48f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h563b4d42c1a8eb1bed0decf6c754f70f5b485f0b17cf0f90b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3b13ec24032f1e472a6da4dab8431ce51770d424f224cbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84eec04a5677ed21d94579aded9acbd101d00c48df02361d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h182d0cb33631e83d9646d78150747019ff5901d3e96ea77d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd53b775d7fe774a9e235b1d97ee1771ac9b712437268e6ed4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haee630c7e8dc5b651e32893baea0a6df7d9981184a2c28e70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec131ad210f5708e1d091597b13a3e94b1987a7d2396b2a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h608eb55a9d647c09c5f5601fd434d4f400df9ebe3ce2748c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he35428e1ae5e56f0d95b2053265dc0b3683c4fcbce83fe86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa8754512a4757f29e40f7825e7bf3983194698c1fbefafcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2f0bb859908a99187809d52d789299af4ecb3aead85603ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3d8c28db6ef701bda16a6463b0819037a93ca81d29f8da11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74741c031245935432d537fd93d5c240cfbba07bdb363fb89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23c5a8b9b55eddff94e633bfa88f1c04d50249b05eaa105d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44878021ff5d005a32280ff5dd18b747140f249d747e7fcae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c865df8472003c92e1645641688407306d2fe052d8803178;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27f4749b4f194eea9e9734f7ca257eec3fb9c0423a25421e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d1aaca80b4d516fbdd2898b71dd0ca216bc67e10ef1def56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97266225430eb1d1211e63108396f04f79cee0fc40182f0fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f766f700f59dec7b4288dd4d3d92ba411c144b2fb10cc0d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heef8510ac5389c903dc94a93bc270be43bce913bdf37b4e26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefcf51f05a1048390ea4ca325ee6697c6d931681de93d7532;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab159d1747ec9d4a16c9d68d1ec88e57d2a96a8250d958b8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78dcf88d8c57ea88c37466025ea6fbf87c916a5426aff50e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c4048afd4e12add51679ae05b4b4eb734345ea9c7d91bdbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57aa1efd172c77900b38430d2b3165bbe1d31e4e7d321bbf8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd834f7a297d5d3a289773a00c727c08eb493b0c4319a9987c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d8a9178be43ab0d27523b72d6402ab7557d7abb034528d90;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2abd701f78f20bb1d3a9cea73a2dd235c31989bacc8afc777;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc1eed621d9e123cde949fcdc69371d9a8e9421596b4623dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h900b8a0419fbc145adbcba687ec1c8488a4d2b2d81d427e0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e8087abc316b319000427d51dd1d459ee6f90d864a65f681;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81f42ab583339a84ee76190ce4207bd81d4f0bea6f281cb1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74bfeedb86b9fad145654f92fdd9be34cf549e68af91d2c6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5ba98e6dc3ae9f99bd8faccd8cb19f5e856fd872817bbcfc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b278abee606cba2b8f15fdadd69aca2d88092fe77c4a6e6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f268e5bf75ae6783448dc3dd0a2a42fd53d2cb620ab36b00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd0f8bf32deda4a789647e3f26c57c24236598d1a022963ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17ed041d8b44eb12bf9ef312ebf59210cb7513428bfafba96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2173682e8472bab0f3ef8fec02fb00b5cab3ea1b27ed1113;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h330264a516c23a18aaab878eabc977ecc9d201d831517b145;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5ca16db0e32c0fe18c5cdad9ba8c1d23429341daecef6b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0412ed6ed1ec236e55ad5728223a56217e7070b07fc1be19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h774bcefbc7d242b6a4f1fd4f6d6552c729928695cdbe82d7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31335b2f6b075d48e1bf2c8251afd9aed72ae59d4061c296d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e568eceffab3f864de4c3f5258042d92ee5462f0d22cc151;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he920c6dc620ec4cabf908f67fc600fd486b544e2d582bea12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4948068ea7e8c5f44d27e97d9885c5f8e93151446a8751102;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16b4306363dbf7f046c5cbe68bb911f29e80b17def431e04d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1df476ceda0cd6c2c6a09b74d7aa5270aa743b5b9792d8a0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c7f5da246880e43cfe8e48c82bd4b69c9903f9cf147b255a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed15f2bea0d4129a2d830991b28e7ba3bdc5900b149fdda28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b258a21a422b59d39ba46db9e9f36c05aebbb1af2a14e1d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ced17fd648ab85a7b58fb4f618dc3cfb8fe4fe71ce9cadb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h479503b1ea2aa7267ef1ca267cbfdf414a75e13e864ba18ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ac91c78dfa0470a4d38a7d6eccd7deb1f6db08824b2b0c64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0d07e6a249555b2348fe0d9068b6d3a3df782f244b0533e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92fa25a539ebd742d3b1e1e69e474658c499095a8746ec31a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9db9eb7459ec980563ba498b22d1e68b58aaeee58f0ef0740;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h355b30f85329030e1d836c498c207f92bf2b86ec523204e0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc32763ebd8a8bb842e23870ca30f273da23573aea33bb5e31;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f2bd25c84ddd95a98d46ceb7e0f953c8e45e5e366b8f97f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb009836e15757ddaaaeb8dc5187357eeb5ff731f9552a6a14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3540b64011c1d7c7b000426347f48378b1c933dc65f3608c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64b023b6300f875df5a7299c32ce7ead5670529907ec32fdf;
        #1
        $finish();
    end
endmodule
