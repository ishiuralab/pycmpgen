module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    compressor_CLA16_32 compressor_CLA16_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
        src16 <= 16'h0;
        src17 <= 16'h0;
        src18 <= 16'h0;
        src19 <= 16'h0;
        src20 <= 16'h0;
        src21 <= 16'h0;
        src22 <= 16'h0;
        src23 <= 16'h0;
        src24 <= 16'h0;
        src25 <= 16'h0;
        src26 <= 16'h0;
        src27 <= 16'h0;
        src28 <= 16'h0;
        src29 <= 16'h0;
        src30 <= 16'h0;
        src31 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA16_32(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [0:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [0:0] comp_out34;
    wire [1:0] comp_out35;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[1], 1'h0, comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], 1'h0, 1'h0, 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      input wire [15:0] src16,
      input wire [15:0] src17,
      input wire [15:0] src18,
      input wire [15:0] src19,
      input wire [15:0] src20,
      input wire [15:0] src21,
      input wire [15:0] src22,
      input wire [15:0] src23,
      input wire [15:0] src24,
      input wire [15:0] src25,
      input wire [15:0] src26,
      input wire [15:0] src27,
      input wire [15:0] src28,
      input wire [15:0] src29,
      input wire [15:0] src30,
      input wire [15:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [0:0] dst34,
      output wire [1:0] dst35);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [15:0] stage0_16;
   wire [15:0] stage0_17;
   wire [15:0] stage0_18;
   wire [15:0] stage0_19;
   wire [15:0] stage0_20;
   wire [15:0] stage0_21;
   wire [15:0] stage0_22;
   wire [15:0] stage0_23;
   wire [15:0] stage0_24;
   wire [15:0] stage0_25;
   wire [15:0] stage0_26;
   wire [15:0] stage0_27;
   wire [15:0] stage0_28;
   wire [15:0] stage0_29;
   wire [15:0] stage0_30;
   wire [15:0] stage0_31;
   wire [6:0] stage1_0;
   wire [4:0] stage1_1;
   wire [8:0] stage1_2;
   wire [5:0] stage1_3;
   wire [5:0] stage1_4;
   wire [8:0] stage1_5;
   wire [10:0] stage1_6;
   wire [6:0] stage1_7;
   wire [5:0] stage1_8;
   wire [8:0] stage1_9;
   wire [5:0] stage1_10;
   wire [5:0] stage1_11;
   wire [10:0] stage1_12;
   wire [6:0] stage1_13;
   wire [6:0] stage1_14;
   wire [6:0] stage1_15;
   wire [9:0] stage1_16;
   wire [12:0] stage1_17;
   wire [5:0] stage1_18;
   wire [5:0] stage1_19;
   wire [5:0] stage1_20;
   wire [5:0] stage1_21;
   wire [8:0] stage1_22;
   wire [6:0] stage1_23;
   wire [6:0] stage1_24;
   wire [7:0] stage1_25;
   wire [10:0] stage1_26;
   wire [5:0] stage1_27;
   wire [7:0] stage1_28;
   wire [5:0] stage1_29;
   wire [11:0] stage1_30;
   wire [8:0] stage1_31;
   wire [2:0] stage1_32;
   wire [1:0] stage1_33;
   wire [0:0] stage1_34;
   wire [1:0] stage2_0;
   wire [1:0] stage2_1;
   wire [4:0] stage2_2;
   wire [1:0] stage2_3;
   wire [2:0] stage2_4;
   wire [5:0] stage2_5;
   wire [2:0] stage2_6;
   wire [2:0] stage2_7;
   wire [2:0] stage2_8;
   wire [5:0] stage2_9;
   wire [2:0] stage2_10;
   wire [1:0] stage2_11;
   wire [6:0] stage2_12;
   wire [3:0] stage2_13;
   wire [2:0] stage2_14;
   wire [1:0] stage2_15;
   wire [6:0] stage2_16;
   wire [4:0] stage2_17;
   wire [2:0] stage2_18;
   wire [5:0] stage2_19;
   wire [2:0] stage2_20;
   wire [2:0] stage2_21;
   wire [3:0] stage2_22;
   wire [1:0] stage2_23;
   wire [2:0] stage2_24;
   wire [6:0] stage2_25;
   wire [5:0] stage2_26;
   wire [1:0] stage2_27;
   wire [5:0] stage2_28;
   wire [4:0] stage2_29;
   wire [1:0] stage2_30;
   wire [5:0] stage2_31;
   wire [2:0] stage2_32;
   wire [1:0] stage2_33;
   wire [0:0] stage2_34;
   wire [0:0] stage2_35;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [1:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage3_21;
   wire [1:0] stage3_22;
   wire [1:0] stage3_23;
   wire [1:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [1:0] stage3_27;
   wire [1:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [1:0] stage3_31;
   wire [1:0] stage3_32;
   wire [1:0] stage3_33;
   wire [0:0] stage3_34;
   wire [1:0] stage3_35;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;
   assign dst20 = stage3_20;
   assign dst21 = stage3_21;
   assign dst22 = stage3_22;
   assign dst23 = stage3_23;
   assign dst24 = stage3_24;
   assign dst25 = stage3_25;
   assign dst26 = stage3_26;
   assign dst27 = stage3_27;
   assign dst28 = stage3_28;
   assign dst29 = stage3_29;
   assign dst30 = stage3_30;
   assign dst31 = stage3_31;
   assign dst32 = stage3_32;
   assign dst33 = stage3_33;
   assign dst34 = stage3_34;
   assign dst35 = stage3_35;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[0],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[1],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[2],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc615_5 gpc4 (
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage0_3[12]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[3],stage1_3[4],stage1_2[4]}
   );
   gpc1343_5 gpc5 (
      {stage0_3[13], stage0_3[14], stage0_3[15]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[4],stage1_3[5]}
   );
   gpc1406_5 gpc6 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[5]}
   );
   gpc606_5 gpc7 (
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage1_9[0],stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc615_5 gpc8 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13]},
      {stage0_6[5]},
      {stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12]},
      {stage1_9[1],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc615_5 gpc9 (
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10]},
      {stage0_7[13]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[3],stage1_7[4],stage1_6[5]}
   );
   gpc615_5 gpc10 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[3],stage1_8[4]}
   );
   gpc615_5 gpc11 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[1]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[4],stage1_8[5]}
   );
   gpc606_5 gpc12 (
      {stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[5]}
   );
   gpc606_5 gpc13 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[6]}
   );
   gpc615_5 gpc14 (
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], 1'b0},
      {stage0_11[12]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[2],stage1_12[4],stage1_11[4],stage1_10[5]}
   );
   gpc615_5 gpc15 (
      {stage0_11[13], stage0_11[14], stage0_11[15], 1'b0, 1'b0},
      {stage0_12[6]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[3],stage1_12[5],stage1_11[5]}
   );
   gpc1343_5 gpc16 (
      {stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9]},
      {stage0_14[0], stage0_14[1], stage0_14[2]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[1],stage1_14[2],stage1_13[4],stage1_12[6]}
   );
   gpc623_5 gpc17 (
      {stage0_12[10], stage0_12[11], stage0_12[12]},
      {stage0_13[10], stage0_13[11]},
      {stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8]},
      {stage1_16[1],stage1_15[2],stage1_14[3],stage1_13[5],stage1_12[7]}
   );
   gpc615_5 gpc18 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], 1'b0},
      {stage0_14[9]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[2],stage1_15[3],stage1_14[4],stage1_13[6]}
   );
   gpc1343_5 gpc19 (
      {stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10]},
      {stage0_16[0], stage0_16[1], stage0_16[2]},
      {stage0_17[0]},
      {stage1_18[0],stage1_17[1],stage1_16[3],stage1_15[4],stage1_14[5]}
   );
   gpc1343_5 gpc20 (
      {stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage0_15[11], stage0_15[12], stage0_15[13], stage0_15[14]},
      {stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage0_17[1]},
      {stage1_18[1],stage1_17[2],stage1_16[4],stage1_15[5],stage1_14[6]}
   );
   gpc606_5 gpc21 (
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[3],stage1_16[5]}
   );
   gpc606_5 gpc22 (
      {stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[4]}
   );
   gpc615_5 gpc23 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10]},
      {stage0_19[6]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[1],stage1_20[2],stage1_19[2],stage1_18[4]}
   );
   gpc615_5 gpc24 (
      {stage0_18[11], stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15]},
      {stage0_19[7]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[2],stage1_20[3],stage1_19[3],stage1_18[5]}
   );
   gpc1343_5 gpc25 (
      {stage0_19[8], stage0_19[9], stage0_19[10]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15]},
      {stage0_21[0], stage0_21[1], stage0_21[2]},
      {stage0_22[0]},
      {stage1_23[0],stage1_22[2],stage1_21[3],stage1_20[4],stage1_19[4]}
   );
   gpc615_5 gpc26 (
      {stage0_19[11], stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15]},
      {1'b0},
      {stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7], stage0_21[8]},
      {stage1_23[1],stage1_22[3],stage1_21[4],stage1_20[5],stage1_19[5]}
   );
   gpc207_4 gpc27 (
      {stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[0], stage0_23[1]},
      {stage1_24[0],stage1_23[2],stage1_22[4],stage1_21[5]}
   );
   gpc2135_5 gpc28 (
      {stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage0_23[2], stage0_23[3], stage0_23[4]},
      {stage0_24[0]},
      {stage0_25[0], stage0_25[1]},
      {stage1_26[0],stage1_25[0],stage1_24[1],stage1_23[3],stage1_22[5]}
   );
   gpc1163_5 gpc29 (
      {stage0_22[6], stage0_22[7], stage0_22[8]},
      {stage0_23[5], stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10]},
      {stage0_24[1]},
      {stage0_25[2]},
      {stage1_26[1],stage1_25[1],stage1_24[2],stage1_23[4],stage1_22[6]}
   );
   gpc606_5 gpc30 (
      {stage0_22[9], stage0_22[10], stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6], stage0_24[7]},
      {stage1_26[2],stage1_25[2],stage1_24[3],stage1_23[5],stage1_22[7]}
   );
   gpc615_5 gpc31 (
      {stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage0_24[8]},
      {stage0_25[3], stage0_25[4], stage0_25[5], stage0_25[6], stage0_25[7], stage0_25[8]},
      {stage1_27[0],stage1_26[3],stage1_25[3],stage1_24[4],stage1_23[6]}
   );
   gpc606_5 gpc32 (
      {stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12], stage0_24[13], stage0_24[14]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[4],stage1_25[4],stage1_24[5]}
   );
   gpc1415_5 gpc33 (
      {stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13]},
      {stage0_26[6]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3]},
      {stage0_28[0]},
      {stage1_29[0],stage1_28[1],stage1_27[2],stage1_26[5],stage1_25[5]}
   );
   gpc615_5 gpc34 (
      {stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage0_27[4]},
      {stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5], stage0_28[6]},
      {stage1_30[0],stage1_29[1],stage1_28[2],stage1_27[3],stage1_26[6]}
   );
   gpc606_5 gpc35 (
      {stage0_27[5], stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[2],stage1_28[3],stage1_27[4]}
   );
   gpc615_5 gpc36 (
      {stage0_27[11], stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15]},
      {stage0_28[7]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[2],stage1_29[3],stage1_28[4],stage1_27[5]}
   );
   gpc606_5 gpc37 (
      {stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[3],stage1_29[4],stage1_28[5]}
   );
   gpc615_5 gpc38 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], 1'b0},
      {stage0_30[6]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[1],stage1_31[3],stage1_30[4],stage1_29[5]}
   );
   gpc1163_5 gpc39 (
      {stage0_30[7], stage0_30[8], stage0_30[9]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {1'b0},
      {1'b0},
      {stage1_34[0],stage1_33[1],stage1_32[2],stage1_31[4],stage1_30[5]}
   );
   gpc1_1 gpc40 (
      {stage0_0[11]},
      {stage1_0[2]}
   );
   gpc1_1 gpc41 (
      {stage0_0[12]},
      {stage1_0[3]}
   );
   gpc1_1 gpc42 (
      {stage0_0[13]},
      {stage1_0[4]}
   );
   gpc1_1 gpc43 (
      {stage0_0[14]},
      {stage1_0[5]}
   );
   gpc1_1 gpc44 (
      {stage0_0[15]},
      {stage1_0[6]}
   );
   gpc1_1 gpc45 (
      {stage0_1[15]},
      {stage1_1[4]}
   );
   gpc1_1 gpc46 (
      {stage0_2[12]},
      {stage1_2[5]}
   );
   gpc1_1 gpc47 (
      {stage0_2[13]},
      {stage1_2[6]}
   );
   gpc1_1 gpc48 (
      {stage0_2[14]},
      {stage1_2[7]}
   );
   gpc1_1 gpc49 (
      {stage0_2[15]},
      {stage1_2[8]}
   );
   gpc1_1 gpc50 (
      {stage0_5[14]},
      {stage1_5[7]}
   );
   gpc1_1 gpc51 (
      {stage0_5[15]},
      {stage1_5[8]}
   );
   gpc1_1 gpc52 (
      {stage0_6[11]},
      {stage1_6[6]}
   );
   gpc1_1 gpc53 (
      {stage0_6[12]},
      {stage1_6[7]}
   );
   gpc1_1 gpc54 (
      {stage0_6[13]},
      {stage1_6[8]}
   );
   gpc1_1 gpc55 (
      {stage0_6[14]},
      {stage1_6[9]}
   );
   gpc1_1 gpc56 (
      {stage0_6[15]},
      {stage1_6[10]}
   );
   gpc1_1 gpc57 (
      {stage0_7[14]},
      {stage1_7[5]}
   );
   gpc1_1 gpc58 (
      {stage0_7[15]},
      {stage1_7[6]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[7]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[8]}
   );
   gpc1_1 gpc61 (
      {stage0_12[13]},
      {stage1_12[8]}
   );
   gpc1_1 gpc62 (
      {stage0_12[14]},
      {stage1_12[9]}
   );
   gpc1_1 gpc63 (
      {stage0_12[15]},
      {stage1_12[10]}
   );
   gpc1_1 gpc64 (
      {stage0_15[15]},
      {stage1_15[6]}
   );
   gpc1_1 gpc65 (
      {stage0_16[12]},
      {stage1_16[6]}
   );
   gpc1_1 gpc66 (
      {stage0_16[13]},
      {stage1_16[7]}
   );
   gpc1_1 gpc67 (
      {stage0_16[14]},
      {stage1_16[8]}
   );
   gpc1_1 gpc68 (
      {stage0_16[15]},
      {stage1_16[9]}
   );
   gpc1_1 gpc69 (
      {stage0_17[8]},
      {stage1_17[5]}
   );
   gpc1_1 gpc70 (
      {stage0_17[9]},
      {stage1_17[6]}
   );
   gpc1_1 gpc71 (
      {stage0_17[10]},
      {stage1_17[7]}
   );
   gpc1_1 gpc72 (
      {stage0_17[11]},
      {stage1_17[8]}
   );
   gpc1_1 gpc73 (
      {stage0_17[12]},
      {stage1_17[9]}
   );
   gpc1_1 gpc74 (
      {stage0_17[13]},
      {stage1_17[10]}
   );
   gpc1_1 gpc75 (
      {stage0_17[14]},
      {stage1_17[11]}
   );
   gpc1_1 gpc76 (
      {stage0_17[15]},
      {stage1_17[12]}
   );
   gpc1_1 gpc77 (
      {stage0_22[15]},
      {stage1_22[8]}
   );
   gpc1_1 gpc78 (
      {stage0_24[15]},
      {stage1_24[6]}
   );
   gpc1_1 gpc79 (
      {stage0_25[14]},
      {stage1_25[6]}
   );
   gpc1_1 gpc80 (
      {stage0_25[15]},
      {stage1_25[7]}
   );
   gpc1_1 gpc81 (
      {stage0_26[12]},
      {stage1_26[7]}
   );
   gpc1_1 gpc82 (
      {stage0_26[13]},
      {stage1_26[8]}
   );
   gpc1_1 gpc83 (
      {stage0_26[14]},
      {stage1_26[9]}
   );
   gpc1_1 gpc84 (
      {stage0_26[15]},
      {stage1_26[10]}
   );
   gpc1_1 gpc85 (
      {stage0_28[14]},
      {stage1_28[6]}
   );
   gpc1_1 gpc86 (
      {stage0_28[15]},
      {stage1_28[7]}
   );
   gpc1_1 gpc87 (
      {stage0_30[10]},
      {stage1_30[6]}
   );
   gpc1_1 gpc88 (
      {stage0_30[11]},
      {stage1_30[7]}
   );
   gpc1_1 gpc89 (
      {stage0_30[12]},
      {stage1_30[8]}
   );
   gpc1_1 gpc90 (
      {stage0_30[13]},
      {stage1_30[9]}
   );
   gpc1_1 gpc91 (
      {stage0_30[14]},
      {stage1_30[10]}
   );
   gpc1_1 gpc92 (
      {stage0_30[15]},
      {stage1_30[11]}
   );
   gpc1_1 gpc93 (
      {stage0_31[12]},
      {stage1_31[5]}
   );
   gpc1_1 gpc94 (
      {stage0_31[13]},
      {stage1_31[6]}
   );
   gpc1_1 gpc95 (
      {stage0_31[14]},
      {stage1_31[7]}
   );
   gpc1_1 gpc96 (
      {stage0_31[15]},
      {stage1_31[8]}
   );
   gpc606_5 gpc97 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc98 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], 1'b0},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc99 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc100 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc615_5 gpc101 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[2],stage2_6[2]}
   );
   gpc606_5 gpc102 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1],stage2_9[2]}
   );
   gpc606_5 gpc103 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[2]}
   );
   gpc606_5 gpc104 (
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[2]}
   );
   gpc117_4 gpc105 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage1_15[6]},
      {stage1_16[0]},
      {stage2_17[1],stage2_16[1],stage2_15[1],stage2_14[2]}
   );
   gpc1163_5 gpc106 (
      {stage1_16[1], stage1_16[2], stage1_16[3]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_18[0]},
      {stage1_19[0]},
      {stage2_20[0],stage2_19[0],stage2_18[0],stage2_17[2],stage2_16[2]}
   );
   gpc1163_5 gpc107 (
      {stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_18[1]},
      {stage1_19[1]},
      {stage2_20[1],stage2_19[1],stage2_18[1],stage2_17[3],stage2_16[3]}
   );
   gpc615_5 gpc108 (
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], 1'b0},
      {stage1_19[2]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[2]}
   );
   gpc1163_5 gpc109 (
      {stage1_21[0], stage1_21[1], stage1_21[2]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_23[0]},
      {stage1_24[0]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[1]}
   );
   gpc623_5 gpc110 (
      {stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_22[6], stage1_22[7]},
      {stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5], stage1_23[6]},
      {stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2],stage2_21[2]}
   );
   gpc606_5 gpc111 (
      {stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[0],stage2_26[0],stage2_25[2],stage2_24[2]}
   );
   gpc615_5 gpc112 (
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4]},
      {stage1_26[6]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[1],stage2_27[1],stage2_26[1],stage2_25[3]}
   );
   gpc615_5 gpc113 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4]},
      {stage1_29[0]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[0],stage2_30[0],stage2_29[1],stage2_28[2]}
   );
   gpc1163_5 gpc114 (
      {stage1_29[1], stage1_29[2], stage1_29[3]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_31[0]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[1],stage2_31[1],stage2_30[1],stage2_29[2]}
   );
   gpc1325_5 gpc115 (
      {stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage1_32[1], stage1_32[2]},
      {stage1_33[0], stage1_33[1], 1'b0},
      {stage1_34[0]},
      {stage2_35[0],stage2_34[0],stage2_33[1],stage2_32[2],stage2_31[2]}
   );
   gpc1_1 gpc116 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc117 (
      {stage1_2[6]},
      {stage2_2[2]}
   );
   gpc1_1 gpc118 (
      {stage1_2[7]},
      {stage2_2[3]}
   );
   gpc1_1 gpc119 (
      {stage1_2[8]},
      {stage2_2[4]}
   );
   gpc1_1 gpc120 (
      {stage1_5[6]},
      {stage2_5[3]}
   );
   gpc1_1 gpc121 (
      {stage1_5[7]},
      {stage2_5[4]}
   );
   gpc1_1 gpc122 (
      {stage1_5[8]},
      {stage2_5[5]}
   );
   gpc1_1 gpc123 (
      {stage1_9[6]},
      {stage2_9[3]}
   );
   gpc1_1 gpc124 (
      {stage1_9[7]},
      {stage2_9[4]}
   );
   gpc1_1 gpc125 (
      {stage1_9[8]},
      {stage2_9[5]}
   );
   gpc1_1 gpc126 (
      {stage1_12[6]},
      {stage2_12[2]}
   );
   gpc1_1 gpc127 (
      {stage1_12[7]},
      {stage2_12[3]}
   );
   gpc1_1 gpc128 (
      {stage1_12[8]},
      {stage2_12[4]}
   );
   gpc1_1 gpc129 (
      {stage1_12[9]},
      {stage2_12[5]}
   );
   gpc1_1 gpc130 (
      {stage1_12[10]},
      {stage2_12[6]}
   );
   gpc1_1 gpc131 (
      {stage1_13[6]},
      {stage2_13[3]}
   );
   gpc1_1 gpc132 (
      {stage1_16[7]},
      {stage2_16[4]}
   );
   gpc1_1 gpc133 (
      {stage1_16[8]},
      {stage2_16[5]}
   );
   gpc1_1 gpc134 (
      {stage1_16[9]},
      {stage2_16[6]}
   );
   gpc1_1 gpc135 (
      {stage1_17[12]},
      {stage2_17[4]}
   );
   gpc1_1 gpc136 (
      {stage1_19[3]},
      {stage2_19[3]}
   );
   gpc1_1 gpc137 (
      {stage1_19[4]},
      {stage2_19[4]}
   );
   gpc1_1 gpc138 (
      {stage1_19[5]},
      {stage2_19[5]}
   );
   gpc1_1 gpc139 (
      {stage1_22[8]},
      {stage2_22[3]}
   );
   gpc1_1 gpc140 (
      {stage1_25[5]},
      {stage2_25[4]}
   );
   gpc1_1 gpc141 (
      {stage1_25[6]},
      {stage2_25[5]}
   );
   gpc1_1 gpc142 (
      {stage1_25[7]},
      {stage2_25[6]}
   );
   gpc1_1 gpc143 (
      {stage1_26[7]},
      {stage2_26[2]}
   );
   gpc1_1 gpc144 (
      {stage1_26[8]},
      {stage2_26[3]}
   );
   gpc1_1 gpc145 (
      {stage1_26[9]},
      {stage2_26[4]}
   );
   gpc1_1 gpc146 (
      {stage1_26[10]},
      {stage2_26[5]}
   );
   gpc1_1 gpc147 (
      {stage1_28[5]},
      {stage2_28[3]}
   );
   gpc1_1 gpc148 (
      {stage1_28[6]},
      {stage2_28[4]}
   );
   gpc1_1 gpc149 (
      {stage1_28[7]},
      {stage2_28[5]}
   );
   gpc1_1 gpc150 (
      {stage1_29[4]},
      {stage2_29[3]}
   );
   gpc1_1 gpc151 (
      {stage1_29[5]},
      {stage2_29[4]}
   );
   gpc1_1 gpc152 (
      {stage1_31[6]},
      {stage2_31[3]}
   );
   gpc1_1 gpc153 (
      {stage1_31[7]},
      {stage2_31[4]}
   );
   gpc1_1 gpc154 (
      {stage1_31[8]},
      {stage2_31[5]}
   );
   gpc1325_5 gpc155 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[0], stage2_3[1]},
      {stage2_4[0], stage2_4[1], stage2_4[2]},
      {stage2_5[0]},
      {stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0]}
   );
   gpc2135_5 gpc156 (
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc615_5 gpc157 (
      {stage2_7[1], stage2_7[2], 1'b0, 1'b0, 1'b0},
      {stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[1],stage3_8[1],stage3_7[1]}
   );
   gpc623_5 gpc158 (
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0], stage2_11[1]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[1]}
   );
   gpc135_4 gpc159 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[0],stage3_14[1],stage3_13[1]}
   );
   gpc207_4 gpc160 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[1]}
   );
   gpc615_5 gpc161 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4]},
      {stage2_18[2]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[1],stage3_17[1]}
   );
   gpc1343_5 gpc162 (
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0], stage2_21[1], stage2_21[2], 1'b0},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage3_24[0],stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[1]}
   );
   gpc1163_5 gpc163 (
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_26[0]},
      {stage2_27[0]},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1]}
   );
   gpc615_5 gpc164 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage2_27[1]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1]}
   );
   gpc2135_5 gpc165 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4]},
      {stage2_30[0], stage2_30[1], 1'b0},
      {stage2_31[0]},
      {stage2_32[0], stage2_32[1]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[1]}
   );
   gpc1325_5 gpc166 (
      {stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_32[2], 1'b0},
      {stage2_33[0], stage2_33[1], 1'b0},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[0],stage3_33[1],stage3_32[1],stage3_31[1]}
   );
   gpc1_1 gpc167 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc168 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc169 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc170 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc171 (
      {stage2_12[6]},
      {stage3_12[1]}
   );
   gpc1_1 gpc172 (
      {stage2_15[1]},
      {stage3_15[1]}
   );
   gpc1_1 gpc173 (
      {stage2_22[3]},
      {stage3_22[1]}
   );
   gpc1_1 gpc174 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc175 (
      {stage2_25[6]},
      {stage3_25[1]}
   );
   gpc1_1 gpc176 (
      {stage2_35[0]},
      {stage3_35[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor_CLA16_32 compressor_CLA16_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc62dbd0348bc254188efb178470fd3502cccf8f2bb1b89f00dd0de0c8c1d9b19ab46ee90e96d984a5e4e174bf78d9b96de27380cf778564641d71fd5b464f4cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h42d5d98c562e012fd01990c0057a8c5b9818084328ac3c34abb8fac7a0dfbe0e10627d5a50e94f9cc09d5bfb1675d563bd62ac1e17b90859ca7d8c0b22ebc393;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h219f55018b93b5fae0c31fc55791aefe4a4b5941838b67bb94e998174e5749c6855896cf8b8f713bd69aa3e891c2afdb9da5a0a04a04554f9ac6d7b94fc5bb02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb4d41c98438507d513e04c6788fe8425f82753a58b4e77265e7ee2358e04c0e5d8ebce06a974b59ce0eb1dc9c792e5ec274c5af04117b9e44ee776112f7355d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7ec5cc28f3201ddaa38af17aaf011cfb9871da2f5cea8f6004f1928f012a65f08b323f95e34b90be3e13b514c49b9e503182697d30c34553e3b4ec233c975c29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hea2d70c2933c314152492e8d3f1aa617b43b060fd21c787019923ebcab2fb7cc71dc0b818fbebbdede54a8c5b28968f6b2d5cb6367f6e5839eb13799acfdb0ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1d96e8401ac888670b2b4b3d62c3b7c03124ca708278f43471969ca63f15788bf6226fdb25ec42f53408113101815710d0c140b06692a1632531ed3dd0dcf5b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h77832542737c5b635e5cb2daa4113355d1f2a3293639f8a8c82fe8e00f5bf4a1cf56cec52b05059e402d5ba0c43c05a190fa26a0f2567546fd59b32a96bbdacb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h30a0ccc68463534de4a3c6fbcd95fd8c5f4bd2e8116ca9f1e1ee23e6edbe92b3c4f4927d3f4f06dcb3ef935d053069cd7d05cd9b677976bd46097b397a8eb316;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd1595581b312f5dd27ea9fa6ead1e85ab9535ac6ea93527b576d2490988a5bbb8f7a87815b6b39996f27fa32321edc4f2e7037704f356a215761496b30046adb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h859804d53c61f067fe8df64f875864b7b8c3f3b0c955aef00726b0ab1fccf1746e2672f486c89f697a2685603056717b906ea5fe39c2ff40534058b4f845c0d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf44fa86496dd923c85f78032e9d4aa56f80ed5d0de9f563af2dbc8a431243b41a549a1717d164707988c0726b122007ccfcf059044fab2a5d29e641a20cc1c48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h87a4affc0001cad6fe81118cc743c878ef71d14aedb7a7900d4b7e7979048803133345fd9ef621e835641a5c9657cb12c72290089a7d9582e573ece34df7cadf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h358619b3afc50655defda46df0361b1c3e051f25155a5a5b1fd0600cd6f8787dfa5480ed5171d6585494c8957cb64cfafed951da246e95ee3137f70186d2bbce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5d6d7f1e7951f56668540d12bc7f3e5800a01dfe303f39c8b85b29be73269eed8cb7f1002059a1960f926010b89592414c8825a7acd3917bac082c7189f3199e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h16d107274b6b5e980aeb010ae2628935e2c1b5c9f1021efacd8f3bc4371446f472f34d478d4468174a06b1581de9f7510fb62ca8f39d85241783829fe8d02ee9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5dbc4ba437df53ff83591a2be9bfc2f2b2b9c8b49ef4758698ae26214f3c9817c041f9caa6d6b8819c4803e34c76e26ec3658aada899edd119046e7e53d1be08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1a92356400ca1af5943925f6f9faace47a47aa287de5d08d9be2d6e03976db1f0993f9f23c17159c5304c7602ee8a72471b0edead0bb456683d6f7e1787e00d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h174e1e2db3ff7c6524ae36b35bcada9196dfa8cd1e7493e0bd3120bc9cd73d578c01e490a79238255857616fb9c033e90aab9d9edeffd4d30ff21bc0b78be105;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h97e4be8951e6e7dfbf5901e5b50ba0f47dcd819d1ba60061015d17b2dd1b9a45e38a5a4b6af664e12af12c70845b8bf0deb66d384427cf67bb718008ddddd714;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3c517155677547cc1fa00b8f7a9ccf9a9a200a6765861c22bc1c08b4774025fb0a8a6d48b3f441565db5be172c76382ab5f74bac0b9bc88b73e4caaf002a9eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3753f2cbc55ce0262ce6c228f16f6c2c5520b6d001155686bb0169fa373ee1d5b7233f380a4fde41330a77c5a56e6f2af3487674b851d96fe5f8e123c78591c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h43f10a52e3938413c1db959566e6d282211b4cfc49beebf49b15929d9fd48fa6f7b05ce795eede551d2a313c04a5416fea60267ba330c15b7f2066c5b9cb3205;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h22a7c95bf906f7ac1acfac9307c53af977a4068d2269e6775013564aba140ba5a44c6e86d5f6d5c8a2476aa5b704f6be19e58256c10f1e0af3bf0a22d443ac94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf566dc5f759d6e5d9b8bd764d8a8a0964be198f154b6fd8089f5936642e8ffa3d77a83ccef27180706a819135a96c3fd0ce4a3f54beb99d08b256f5d334edda8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcd4a3bdd5f18e95efdf1cdbf51bda00cd73281b1378e6c491018bfdfe715012c438ea59ebb03a05fbf1ac5b71c0dfbb0209149bb0f653c6255fab7b50f8b2340;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h532220621cb94b8b3176ab85c8f08db1ad34e993763338ccfe04c25baadd8b17e3674ba9fe5a527ee8ba34bc183797c202d9b334524a241415c25583defee71f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb451f776ab99bdd06cd76a7d88bf652ab056e02ce9ed9c79d83080c88d28b675d8a032f3b0152442197fefdbb83ccd33737b097a31607005399bcab01c12aefe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2dba877d8a96d2de8311acb50be04b8209018662ca44db00cba1a8a7655f94b466d63fcf26d748ccb761b71cf74d61b13395ff72d379b5273797c9ad7ce7ca7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h383132f4aee2cd9383a316d8f0c428bd097511d2085eb3092885e3371d08c5a8c134f04f9590d05ee6cc24f7ccaa2114f81df96acca2d9444d8dc57f3b20c79e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h11fbd0366392748096e312cf2dbeb4bffad3dbbe7c92e22436a52545771e3a57ea24a98b2231e937b464a35e540e0490c48773dc321067e3702bf488f94422f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h16ec168ba64b6e265ebbafca2ec8fb64346251075cd8d9ddc572a597cb8b419a62e59396ddc7f2a57e5bb8a8adc4baad1e26708ca24b09510b5e14f894492caa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4dd73354339314ea1d4fd4176addced64e0a3a515080582c048a73211c88f0ab159b4d551df436261dd22f7572ae8f27e206cf8117be83012db9d03cdd27e805;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h36144d175f68b7ab07cc8712492a96cbd49ca602c6df65c62203f71e0e858a9399386d6273b31ed65cd62bc8de60b3b593ebbcba938b81e24b1875a2d3d9207;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he3e31ee9e446f8487ede50c5b782003dc1e49ab7c432d324b6108227efa347c5714dfe514b3b72832a528cd5c621155dd001c47c022f680a4e4e633662a077ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2bfb8dfe882e0eabdd2e6af0417825df4aace04469981b1a5d5ef1c227aa462444da622bee2d7ebed5b9af6b83f3daae58a29ee43bfeddc1d1f20e42d0032c53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5cfaf89fd0b88f8c5d6a5d84fc95f8fdb72e13612501cb1e65745906e729f194ad11888767e0ba3acda654bfdaa18fb2792437e95312106eea694e9d346d7b55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h40f4bd90546d3ef00afc810ea066fab65a5d3069dc39ed0b21514ddb64bedc6b3ee0a12d3ff45f645675f32bbedcd03e6524be38cb4cdd19249da3b52c9da870;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4d5d95473c2bf497697c9d5d1396da5a562a3119491628cbf3548a918f91c33f7bf773bfeeb773704bab61e33c3dc98e4a87b382f1a17220f82f5708f44d9c4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd71128f44320bda778abf92ce4e077f4e90fe805213ebadc4006b3567d1e281f14562c851ac0172c5661bc58e747a1978a891b8000ccca9330576c0f91b76caf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'heeb00107bdd535623828da6d06d629014b70f70b71b985f6c06c28fc4ba86e2c49611a61b2da7100c1da3db8018dcdcdea343c6db3802f3da0a0efcd1ef4b0a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h54f4e953d1dd635ff0c221113267d36d6a3db0e3dd562f50b5f786e6c6cbf4eeb206d96937a161cd57fed21ca523bad1932f63c98e153d820f8f47a6f06d19e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h12dd371122d037418adaac1607361ec909bda83d0b11ff71c8f80a264628057310041e96dd37ea58d76ac8db4c07620c19362d169859cdec390d02d63e48d753;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc634087840da7784fe752bf6f75d7ff17bcf16c79bd093d3a88b60bc7c1f465360252af9263444455ca945ec2a81f6c8f3d294d7fcd4921f70571434b23d619;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h136bf50464a6f6461804a7f9e91b03abb2327a42c184b6445769046793d7ac6b27f56dff6fcb95af966d9b1de28fc8d70a8e61e01ba8544cdceffcfbc80bd453;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcb41cd641908405b7cff884025f0a89c20f0de5db547988710dfb4d3940e10943f228b109354420c7ffdd118990e9234cd15f9e7badb5d00d6f506e973f553b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1593232fc9cb2fd218768331556f8b27b0913597f7b1f270c80829e7604a754b4f87e50d28d2a3fd885ede927e244d5f35f1e6a0b8322cc72439d9dfae8b10e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h83e2be12fc611bbc4c38642ab9760e55f672af915b45683b3afaadf68887c93b54141d4a77bb8b0046bb1ce871ef8e8f8153860ecbed20194910b030728dcc5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7fb700353143d3dfb260200b3cb533b080322b5eb5cf053ffd52ba7716a7b48cad3016041bea59e618fab0b7cc36b8d494a7c710b2b4e1575e9fbb04a208ea1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h44e8435bbffa49e8120d6f6c1ca33140da8bcbd724c7c4c7ab251124c947e8ec91807c95131d041c835e2156110b46b711a8905db81f66b97e89d2599b443056;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha8fd135271980dbd745be075a6de17606ad3408af907161dd7398e7419ff3be238e025e95cb0f5144b4845dfbd6b8b4ff938dc619f080ad1286eef1a47f73292;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hee28b6801e03bd9cb670bc2c802a6404a970d92efa6cea2f58650d280a07819f8b3ee9a0b804f1e5cf46a0fdc34f29c22fff129751540344e0caad0d6b9365a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1e3118c8b64e7708113faf8b8d7285674d7da63718dc692ec88a61aed9a76c6cfdb8825494c5cc003e147b44f1c1442d016fd0b597571316ef1dca2f69e219d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h11fb85b518414a841ed34c066c20d7cd1d7eb10f86c6def5f7a683e91e888392d1abeff89fbd926842539e7b3a4be96c62bcf6536762f9aa303708cdfef1f99e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7e4b9171c25767918e8cb16ffe329b2be3963cfb08e09896d93242f44216d380970dcaf697987795fc89133dc3a9ccee4dd8aee05ab29d3b9201187cd215fa39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfad28b53fa1ccfb2e8553d1cd04366cdb7e9124d77ddf09b33260e74e7ba4122d638f9e49285ac8c17934d916d5bfc4629cb18a58b46f6b3ff0136df2de9776c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4bc4cb987490ba4fbc470aa64506fe53106fd4d0ee2a12a98c0ff28f76481361601870c327f0de751cf871a195da80e08d7e128f0861e4f4c6d885c04c09aa1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1831cee11a493787d52e143de8c717dc600b88e44570dc224de2c50915f13cbc79ea64cf17b266abc78489934e93f4437b6fb1829760688e872be0b5a6b48304;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3b2f76fcad53893c53f8a7ff21a60c597abf4e903eb6b3edc82009c9d04cb2cbdfa3bba5ca4e40a43dad9f3da8263a7c6896c7fc0de3df1b37742a4ef82a6868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hef3afd88bfaf4777458130ddc6ec271a9b70feee5fd563094225101f3e8cc3fbf66dad8779c949fc1db98bed2940609e87c55199833f5505fb892a68297db086;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hda6cfeed4fa6e2bbf13e9b0e7e6f1efa640ba5d4f693bc3f22961a8357d80a8e27ab96ed270f1a28d546e0a006d903ea6411168e3ea5d7867f28bde19761943d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5f98261fdb449d1f2d88a90bc8f4c715026d3e8745db450b03fa381de839bb3d428f887a0ddbbb753440bdbeba0b5c4161cc8c3f2df42c28618e13158d3e4511;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb1d37a436bd86e1eefd895d49645cfe45494fe60d2277e655fcbb0c9acd228c6a0549ba9fb0506bcb4d49be88e0368b6c52b17f5f3e672c93e7ee26274836540;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1f8e30ea82cbab14d0f5003d3746a70680f61054cb85c86dc82be8d76365588db33d7ed5307bdac3e545d1f7927da48240abdf00b450339f98c924b3550a233;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2f9b83370ad3d593cdee9e79514ad066e62b63786a6a9e7d3a58bb7dd57b8c78d5c50117e00bf2a660ff8b712d8b4b2b3f15612a2de1cb561451aa76a8427607;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h60aeb637a5ee8491384b18ca8c825fbfa512237fff7fdfe3e674cdfb94d7531d6176b8ff6a8be5000f5aa271e6567af5f7f67f3059f4535b8ce9ae76b4129fb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7d02693abbaaef45b89d1fc6cccc6766a5f390677d6bb32cf3cfe34b798612980c16d2495cd658b04695a3783e6f852a7e31623d81de019307fad6366bcc7151;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb66a2a48c067326212e95c6ba833e448f9cb5220aba05de508b6e927cb88e8510d570f37233493b0e94a4c1b475037e6890718f035c0ee1d777c393f88637af9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h20cdc073e708f7048b326f2ebff0a26a0e0fb6708381691c26151a7b93580fc8a9a4c80352ff19789bfc78bfa1bb9fd9fa3be9232d292f9e0273b838fe9cc538;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb04dfe69ae97c0b33b27524cb20974f984dbb992d1515eaa6179be02f53f2a6506f1f9dffbe6481a4601f1583554f9d5d6cabe1ab9ac98d018e232673854aa2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9f61694959370e86485ade560632365f33618a5d82650ff6235044c75e871c0a92360cfa26093a01560c7c1928ebc6b31e2d4efb0fdc8fc386db6ae30e47ff5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h24bf42e7d84ef0c221a0eb23245f78eeb3608408eccaff25ac37ea15e6b1e606f73a5dd45b8f7f815a5e52e11374c4fe9af1a3c141d5c488f156618fe21373a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h13ac5f042bbedb2f2a940abfe5ed5758cc666feef1fdd88f272bd9c5b2d51f03f97ea80c24f2f4733a571c421e84c54f6289162557edeab65a61318137673a70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3886e5c7e2cb2161d4717c472507943d58b67a8719c6f0957f6b59ac16b73d0493b7a589afc3df77c7e43b135f1d35e1c1f891e93cd87e9f41d287156cd8eae7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc18fd7583745fdbe4cc02e84b79df798d72f81e84cbca48cbba6d7e22fd42c00c307d900e2954ac34f3a1c7621af0db5bc888a6e3e1b56f33a114e95e101d806;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha12490b885649d0f0e4514d1b971717bfc8dd0a9e230da2fa04e19876f0fa30a23ecdf09a871632863ecadd66401587eb0357e6c311a1056d1ab9989863fe6a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3c97a7f964da0bdf095eb59e62d0be7c649d6f324aeb3e2c52e40dad36ab375535763099627c25a4455fbf6177cb107f66bb088f79c3a3d990a0683cce836f36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'heb0e9d8e14c5d8957b5a3ff2fbaaeb17dbeaa86cf6156391afed30a45874dab480eac1bedcfc0f71ced6047d76cc702784060e72fc96baa6eecfda0290e210c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he9bfc3808af9a525b1fad89406967c7d7cf095aa8eb8b84f23d1fc86f1d167ae48b918147267ac0ed3bec52a83be8d23b849616ad1def5932dda54188a6d7836;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf0f38ad6792c61eec9c6c12023a6d4ec8b19abf630e0356127e8f7051265f62ab519c4c08f2c33da0824a90a82e9bf5f86da8458a9efa757832327cd397d7a2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he68180bddabc6babf33a16b7cd21d9817858e44a7dfea27bab7dd1bfd9ba91867a2e9b7794acb7fc7f1204f3f9052c3e0a1bb1e72ae563a1b9217cb01a308a88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h249e6e9138f2563a35de7f66279174ba279d5ba10b836b94d65d3e71726d6185067c308763e89500a3ddcae2f1d0bb827e1812edcc5af23e33d0a3da2d4c0785;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfe57c0fee57f8215ac4ace05790e808db21e88f4f51ee3ef46e2f406a2fc19037a9c6bd14ac2995ff58f208d35073983d40a816fee49bf2445dddbc2119f407f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1d9b523df76eb54295d099a62220f2a1a2c21458ebca83aa67cf59535c5ca79c34a746bbcf8e7ac1331d8cd93dd5e501e468ea6a04ebde25fcb9a631fb3066cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h198a53907601df1a72334b179acac372b43983a167f138734d68bda6dd4c3d407a88768a70bf47c26b5e885ca8f1cd3887bf56bb509f7b0b194cc71acc00d59d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he019ac2731bfe777c6a6187c917e81d23b86d6860309c81c397a629ce17fcc5ad3b67db9d9959132a8a68afbca12fde87f915971f4a466c04cf6b1934da0301a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h523350a97c31ceb504c2b61851724441bb57afc30ed8a54092b1379cdf21ca9b4c0c03fbe32a556534824a38ea17de180eebb1702d0a9ee149f5f9577d42bb87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3656da2c33635b38210d75be6998b6ab19c9a96796ebc1a9e46ecdec9809a47a76ebc48ebba72604622c28110e543755565c2126f300b8624cd692eeaa1fd69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h17ff5459c30db54082ee463eba4c8c86e38aa528a7bb2481123060b7e92fe0043a94da831d426764c830a88cb5bae664d33c6c1093614fc72fe0e60ec3cea32a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1466cbab624ac0161e58517a853a100c2b70eac1302d93d53ecf9b2af962dface46a89e4d4dde1d2b917211422c632b1e3fc739e2981bb641b1c6a213509a9fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6520bfec57c3888ae16638d1dffb7b7fe7e4574281df595a91f1138365145e8e04d35a7b491504a7042ca10d48bd21d5e582a91fee21a409477b2b83e4ecc0e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h91649d977c5eed8e4030b0221c4d44f960be96a8474623be858e313013e8599f60412b364d782aac4dd93eab32027b34d05d505f624b0e5a3edbc85f95f6ce14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha52ad0b7d8d5200c814431ef2fb398ca2275e9826bf598d3bae2d56ad9723cb15f1bacf0723815c8464567971955f7df9d7076b70daadaf6af7f7a80b78b3f9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8a8f7d9a09b86175252bedc85864b6cc1354dafa0f58e009c88a453aabf6774578ae2ed6b3bf4a24c17de1984ddbf5036f134ac33cb182d1d43098e9f8c807e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb8897dfebbae468e3ca53f67f3eb4784bcc505d92467ccaf895f5462adf8f69db3c34860ae82a6f97435248577443f3f1281fb24b8bbe15f59d1eb7ee9dbcf50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha69fe47c0df8074ff74e81f573a7b5799b4e8c826c51896737d47db4d85a944931628a003c7f64975ba38a19de07188848c97cbe6e7ead1d40e33b46423388b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h485473c904afdfb981e23db28d13b0128c97111d1e22b727756c81e18c2f286d756c42f7b4f403d44ea199d90ffaeb1806ff765a3a47784657f905286a4aec7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha1b948c0db49f121095c9049b88963275fe6f922f185497ac2dd1186fa5d5dcdf4c24931d7a195d06fa397caea61e75671c5cc17670c0b53e86ca78e6a183552;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h109d6947bfc60e6bba471a31edaf05a661301dbaf0f1911270e33dadd705be19e04a2bb811665ccb032ac069d7ad4cdcd55df43efe299380c4c82e0c6adf9cf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdc377e6eb8a80de741acdd4b10347cd1213b3f2bdf6e2307eb076e9c8f3fb4350e99b2aedbb18d883a0174c979eddeb8a8a2648b1f0adf440a312989f6c64c35;
        #1
        $finish();
    end
endmodule
