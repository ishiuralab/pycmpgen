module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed2f6222225f3f68cdb3b9c122f687e37c162e094d26e9691;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28e5948c7f948ad956b1a746751aad7107dd43cbe9afcf5c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38af546cac6477684d00884441e1078734c98b19abc6baa4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33872774cb7dae54ba04896adfe579d7e69175e8b509285f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde00da574ff74d699b89927fb93791f281b94a0521c25dfdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb76c16fef75c930d5324b124c2773bebf15e11c97ed86a32e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0d5bcb79f4ff72def5074204f8f6a8f4c2fe2c157ddf0bb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89997519baf52e4b41bb2259cf6b8e2a6c3bcf393bdf301f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53048ff2b15b99e9dd6d7b0591d31f98a8b16711c24f74d40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8e4a2f8422e31d24846baa3e3736419a2fdb2d889b519907;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41ab390da5fcf94f4edf6e9920a837b046c2ee2eb5c12124d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf19d702952dc6c0cc7184df3561772f423e1f1a20ed7357a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0f3d50ccba5a9390368f4be7dff31e4016edf376a24100ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8552ae01df2f5d50929cdc0c6122c5ba09063fed38edcd560;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a3e138361d8959aa5dcfd4b233310532b51cba2de9ceb1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22f2d797dd0a2b6520e54d6aede6661025b427f933b8eac48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5260f1336d853d795ef99d9f3ddb6f7faccd982027dede8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d63cfa04ced01e020fd59a40e085535149f89a509d101770;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31cdc80600bb1f36ea21381a80322b30be27b8dad180e1428;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf645b83fc54b368cbdc9bbba41833674e0f28d05679f24abe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d095b1caeebb6ed6a742de9e9a8a57523d9cb128e52c3d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb42c7642c3badcc07b0f4868d064935112963d90a538f0da3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62c02307954f819129a78448aa3cd149eebb8bb93250606fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81946fe3ff9fc0571894caeaa14ce2a4f88d96d894b476492;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35e4587679fffc94299b8b23d8a856d2a3044b4cf030bc59d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28e8c9d189a3cb92d431b55c853fed40e63def5c76356aa42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84225b79eb0b8ebbfd7c47cca8000ec0358cfc2f147a87ab0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h642edb3c59856a30da9f9ff7c510c514f46b692352a561897;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37e5d9563b1a33cd34ec64f250cddcf2932136a26bde048f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hceb77a33153ce8f18b743a63dd4f8d8d8249dc9913baea167;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h101ba146236a5521b7479ac466f73860b56ee0b1bad51e406;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b72ceebb932d56ed54b6eb5b21fe5ed0a0658591b5054612;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb40c7e05d471c5c526c25ea9be82f46539f68bdf628765b3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1636b02a7e9cdde73c7927349837b8a682d60793b9ba3d7c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbfa0a5f79501cdbe8a860a19e67f546818bb734ff6f4cd8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc4d52fb9a2e3ce54ad214c6a7289608362dee564701662ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha078f56fc23ea8932c9f35b2e8219f835b2de9c0a1d21611c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c5773d03279e9a64e7dcb09069dd720013bb8866bad66bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d2d7c75c9b00598f3715363fdb3d7056b1b9114e31b53b63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff4cd7a649e942286f7b60dc922b3d222caca548f158a2992;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha36a078d516454d0c59bc02f8fbfdf855ed35a882051f8581;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4b46eef9f9721f5087758f9c3fb9afa784f1df7e7c5ce0f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ae16d38a4d9f29bbde30c9c404d71ab9bfdfb3f44d09f68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcec8b219f3b5f6eaf863ddd6c3e1c0851393bbe420f64cf52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eed06ed3ea710b2bd584ed997a4056b89a9d43aa1ec5ff3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64c29cd34fb2d5783c0caecd87be901e1e4eb9f679c1c3559;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h746beb104129dd2d51962a8f8299376f27da6c1ad7fa85700;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93f26a8570488cdbfd57484104f65a8a9c814a8131e65f173;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5f51f0c1e1a7cb4eaf8824b7cbe6ee7be4da5d369c888bc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25a93c41a9875b956ebb34f02f1962255394d34d78fc3cc40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4fe02a9c2b7b5946cc3dac872b6f13a253e483d2544894b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd16548e9da21c98860652ae0f62a8a4e869e76f8893481aa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33ec0cf9df413720991218cfea50c5896d8c7db212f33a249;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7122cc13afd28b83246f02052a6ce942518646db8b0b03be6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dad26607d128536aa6eed431954db72c5a7eac5b955d3ee4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57bbdabc47cf33be5070831a90b620d937e09064da285c09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fcf2ff3fcf9c580d3cfe3e0c94d12715e3e0f21f3775a3a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haad1fee66ddf14b7d328904f6dc2bac492821d3ee1cc0b3d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6380d78f118e75838e8e16024f9251708e63d4802af4bc4e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9a3ee6252246d82f7bf4778c168c03208a8c83d52845aec5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h218f3dbc886d1dd2b899d06f6ddab894e90df9a29cfbf5ee3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b4a7ff44d5825dfedd1e61deab9ebc50331ff6cff0a8a189;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f240ffa5caa088695d873d58844db5d4ec523b47636c5a1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cccccdf93d45fcc0dea6dc135ecafa540344fe06e2873cbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fcfdd5d6f5dd147fd9b5d25139b0acf5f6ef2c7c70c82433;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a8b75fd766091d8cf5826670e741f9b8815f1ec583b6c92b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb04f8d8cab587e70f363409ba27692668cdb524ed2c03208;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a82e5935fca4a53dfab31318a39c38071c49bdcc23af9e49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec23f0188360f6194cde0663a806b2f626ade0a2095425c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65dcab3edfd4043fc04488e175d6d8b95fb8cedc252d4f53c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h943f3a511547886231219ee0362f0066805c7c1e67452a1bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80f7a032c2ccad1667bb5e07c20bb12c70b8785a2597818fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd133883374113a6c8e6c3aad12a69ceda278bd96e57161c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdbce13dcf47a6d59daecc2f3d13550d7cd371c395fe8025a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff775891d7d06163fb74a8ffff2f06d479ae60379ccd5ed5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95b295ee55c354f9f4afbed65a0c02d1bdd3f0c300601c6f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c663d03783f4b7a1f1e81b7d6a30038d6b5f9e3ca131c564;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87511cb3414bf4b2d38237509331b094bee98b6f6b96ae7c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h439098dde86102f098984f89f99be9fb653c273c40eb251b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h635dbafbe0a394e451161d0fb8e6966e0456c88b93322b006;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c12e22b5f2996ea6e039f8c517c1a034fcc59673ba2f7593;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7edc022be4b1d25b5578e5b8b330dbb14888274712836893c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91a36633ce8b580c7607dedea61cc8fd42bcddc251a0b77ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha05602bd19611f49593714f68dda02a6e1c4fb3e0969f37ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26338d6e57c260f7a5ead69dd93c879c1004ed3536982a084;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habfd1f5c04214a802ca3d0c6b08d7197a2cf5697eac998ffa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d2cf4fdbbd021c3d60127007f761683c8da7a3cbf3e91e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf35a99eec7c4a366b621b237c2ee53a446b9f43f0bbcb4718;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4239b8b171cc8dedfce73f42699f12cc75c69ec8b33dbacc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e59b7c5eaba679af92c9f211d9cfb799d05705da53ddfc76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c12d85d491ed05ad249ab8390d900e93d4fddcabeff3ae29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb75dbd5c9d7424a5fc2009d3ae737d7f47722a709a4337fd8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12c5854f74426f9aebf4255526174e347d1a25b9617909ba4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h208f0d11e72a229f70df2089666967731503147d242e2e5e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4042985b41f51796f1487d72040a96b62a44e9c5352d51b8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd523d4ffd7e999ef0f0950abf7c92b61854ad7badcc353164;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cd5d2c82f2d7f88bb09251f79a13ea8f07d83ac65d54ff9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf576a3e09426fc4ad68fbdb3b6350393b481055bf0dec7fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec8806db3344e83da49887a30b4665ac356f15b1cf68b6dbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc51af55ff7b6d6d89588551103232664e6fc20c6c53ae6ca6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h880c579551950c207ccc5e5b543313389bd76a0bdb80f4d1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6602dc13b8a917073b55aec450cf50b3fc78d09922680fab2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h411b8a212f9a811cfeba1afc0b7554ffb67fb07a0dd6afa22;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habc93876d24404c89eeec6d6bfe0cc7ca83c250350fe57a1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb60090effc7917def3b40f46f28f4a2bd878d9408cb1a0ecd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93494b40527ebd82823cd3598325f647de9eca959fd3875ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf339d6e2758cc8fd59fa61c09a24ea8c342e689bc03959293;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2dfffff4cc411f310278fb8bd697debd470616582229f1c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h773d5e67f359af3d5f45f3203121af26e5c7e8565642f95e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd4ed01420936f653122c7e6c8aa52bbfd0f4f87ae63a3504;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68f83abb982543a3204f588a37d736fe8845d6a0fc914f35b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b57cf2aed8c4e5eda5d791e8cfe44914d50bffd030d973e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf05633d7ce45f30c0f28d61fda0dd2f685f43e4a542769f03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bda165697430e89eb56a50d3df4fac3260280050c669ac8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28c96b47b2957049d5a1e9b2182cd111548c0f0f51e713187;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h666989bcf144635a1bb6a1aa312ffb1cec4bb1cbc20ed9dae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he84a8f5214e47a10082e50dd5759ff7be54de62c3a24eff9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fb46d79df23e02ef011dfa1edeec1cd7180f31e6263f3417;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he014692ff1ea457192015e24ae4e4c000153036832e9e48fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h957f95d8df25dad921b4f2efe2348e5e83db9a5786249de3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57fd99a82bbf0b9bf8fca92d2f47d2584628a452cee78d2a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69f8e040e3c006b2fe442b4c677e8a5ff7a2acd7947b3701b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4d670f7208d33f7fda4df6926abdde3301779fb440dd9f66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebda5be31514336904794cdd8041b3e66512a45136f34b90d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa8fd8a28877f977bdca79a8af177ca0d1175fbf45a77b807;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h460cbf2db0df4048ed54b78c381566c955b06781baa6bfd92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6b0c679a1913f22a3a0537bb8ac4e4fa53ec49037b2e26f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f707bfe46767fe5bd2aefc07954dff86b93b72509f27784e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7de8256c8168f335fa88327a57c5b2fdc951184d785fcd382;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf04003ff5293487709ee13c837aa7aabc9cb28690ef52596d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3c8b2d717504218470b3f73891fe1bc280cb48143d21abd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84243b15a37691bcf9b8190ee510432b4777d21527b923d20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e26cb5e120b7a46ea8dcab699b13990580c268781f76cffc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfac50a8c4d35ee5cce95ea1eb739de7c470f0f604419c6ebb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1bd24bd4de75c60c55b828dd70b3e5af0b06f91a3cb9be69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h958b722c6ddaa748efeea5329a360b5d00f9a4a4970fd0b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fc636d96b40de87a648338caf37e225ad143e18bb0a84409;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d945299e402f91a50729950d6f0c688f9e3950955eb714e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf50532607f1ffdba16db28b6f5a809f911f21e40776a6e1bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97a93fee7a8edc5b8bc5b6c98c2d987aab6148f35457f2ead;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c393c6ef684ba7cf7e2c687314509795c494f8b09b723d84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f1e3ee92abdb8e8adf50b45fdd38c5e724db1e24b6ccccf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe83a4ecbe95b406d7166dea578be3275be4657dbd9dca7bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cc2b3489adc38f0d35a1e9d2dd9f8a0a5eeec6831cd4176;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95c4dfc6666ee1203d7b34d77994bb36017a33506a6ac1cad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc917d5e2585f49e8b05af4c6591716dec3e90ad5a6f2cdd8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81b5f64a4b00111638e45a43d84c307f3f30075f3d9143172;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca239c682df819a3e4940d1b70dbca35384d4f8620102074c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he276583517c09c07026cacf7f34af63ae947e1ff333d3039f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0d272c6e0fc5a2a1ad1a65aeeec39c508fa352f997376dbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf14c2a89a73ac070a07d0d5431103382cd2a4266d98ed527d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc57828804e937ba8bdbcdcd2db9c57ff1caf53811c484b9d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f736eb6f1b506c8fe10df82d32be7e8a8161feba39b80256;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h628dc4361d9c1fee0937ef7d0a1bfc6a445749a68e76e6c4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21754d31c2cf66cef0b318c3edb1c0a718569b029bd463341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h178559e727bd952e455fda2c89b19c2a3ae480b316237e632;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2b55f36924cd95dbbb423f91b7e3356bd956abad259a2e0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd95030c270c7970f1ee4d393053046404cc380f0927bc724b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4bf1368af3f63d70f001f6b21b358803f7979caef8445edb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd213bbeab075a107cf780f004d0caaca48963d17a5e7239f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fb1ae11492e829aff448e4f22c35cbc3c14ebca59966b954;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b966a826e419c104fc1b78583a0d9dcd4e49d0f06a509202;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec0ed728b080082de06aa7a23c1ccbfe891fd2be9cd87c34b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac5fd44c79874f3aed9b91fd6f5e2c6d30eec935f791fabc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6e92fbf64aac1c8bdf768cab8111b62769dc3cf14a97c48d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a5c4809eb2a910c472a66dca30979aa1f52ce4ae676b1f64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a10e933cca6aed5fbabadbf2437b635bafdd7f737935be24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3ad6563840fe377139a32092daa04c873c5789379f65835e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65bedc93dff63f9b257f715da0ef0294644935c9420e8c543;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbdbb2dc089f75964330eebcf0a6afafaf0a6886ac85fe71c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63f62c9ee45634518429f0b1ce1ac5503a6cc8999611f3ed7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cdb0cd3c1ec65bb7f56859a8c4f513084654a5588dd5d9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf0dbef28f7ef2b6010ca5abdef2760bd9a0d71893818e319;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93a2ebc7fd8829f3e90f240eba62311e30287ca88d7ff87f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c3da6f81ac30e9d4acc88b3ee8a44f0720d1ae7c23fabfe3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fcb3e68f9543f228e5aedf677d2013caf8880114c952c906;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfb0beba46f62202ff0a26362d47a7c2aca7483e3b934ba8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5911636ac0d8aff1755f7ffcaac62fdca74e92452ccd6363f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bc3066d9772d37a4a8ee984bb8f6af51c7ac4357d12695e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63568a9e393016fc2adb9873a5bc2f0cefb4ecfddbf40a957;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b387e731838abaf1d7278e25d266e914e5423856226b862a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30e9bd19e75efbecd32ae9e8c8e44048b154e150a5e0e59cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h918f6cc1183339e7608306e60ed0705d686e6488fb3e915a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73b400765dd04d99e4086302223b5b58a38ec63cd8b4a5ea9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h682b6564ff2154d9b2e62c0c48adcd98d3c710433202d1ee2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c1cb2224241d11fe6fd5c1403e0e43e3d5b398c03d98660a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9510eadef8ae579cdb0d13e62f71806ede3de0fd21a46d96e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85c12f358aa2ef9495554e6be7258a085902fc2c5325427bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b97542db49d061d4d8268630b1f6b681f9a437faa378fe11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2ef57f0974bb6cfaf4b1b9f128abdbcb2f898b83cc7f559b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2149d0122e1a08b21caa48df30e1bc8dbb0c06f5bc09c339f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7eaf8ff875f17ce25d680f7b92fa460e6e0008bfe72343e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3692274429e5805cff0fa38dae9c13b0328d2e95baabf718;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ddf877ee319132536c25080e25fa2b283d77ea946816e894;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbb3617279cb23f5e982f33a299450f50b11ea9d2fc7fa56a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb89931eb87f4727a0664c44cfebcedabc358b856134107c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c34c73c30b2862ad83d8c629fabcdb4b45951f969f87cd01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a31ee2ae5a9c338056d70721e94939f271b3d272a654ac2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha95a253c9362d6c0c9becac2af5b0c59f6e851cc3f32a63a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae47a13bffeaf3a1e85d48e47e62586bf96a53dc3acb8f598;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38b86028d7ff45ad1746c21ca60ccc852718eff242fcda2a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h622b8be4a8fdd724786385b168c56992216509e20dc3c8d78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedad4a1b578b6dadfedc87b1898ac80dba57e35dadea57afc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e6e0bc6f35a27418afb2558908c4a216292a8e248696d08b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92fa0fdb241e103176d54fe3f2ee4e830c8ed307b5b18d94b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc816163740cfa9048c78b09b7847d09a3a1ad48031248612;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50306167fca9fbe010104fede13f58b16070cdaf5662df9b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h512a8aba458bd5340f96664059aacfd86a48434c397d65f45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h785160e9701117e14e3afb898e078afc6959f1485ca5163ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb43f0ef0d0deb69eff52680d3ac1dcccda1c90b7c7c919337;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h271e4165b9ff3cb6e94eee3711d8bb2ae0862252ae0d6268d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h291f1c4be115decfa846940e4b6c2808a0039fd8ff6946d3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5b6748ef9323455231b1f2d8acf351092c2deaf7e4b43fd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb547b06edf55a427a3a3468e3894e65261a25eb7ec3813b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc668998f42b75291ebda0f94c85c356a840373ec2df4e116b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4337d6acd771dd8950aa098df5dbfbd7cca657a42ec0d5479;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63ed91ea29113646ca2852b6d65fce3a2883d785b8bf01e48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5c381e24a79f5e01db6c031f86ce9801ed1fbfbdc1d3d682;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdca9097f46e8f4af6a353dda3fc715ded2590ff2a1f1ec135;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34e755a05edb5e609b1b8069ca1916c8e51f2d643543d324c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h110d48035a61f6995623212718ded18940b743e889035abb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3939a0fc49d4b26a0e86f0e8a12feb00c434400580be1a69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c3d6ae2ad466ad5550090cab4850f38f8060c09eecfb1545;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he03a5cea05d088242fb8ed4869a1412a332819aa5e588431b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f58b6d1aa2c1051a3eb2637f09965990a9c38d754d355b84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dee329e8058b713b53b2cc4a22132f0d3de9b4e269255a08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc69e105550faf645aa196501d3bbcf52ff9682325a526cc74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ac0ce66297b38c9282e764de98889fad97cbe66fc3e0b902;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a52712ee8337565fbbfcd666721fcf13ae3fc7ab35dc91eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4becc6ba5fde45ac58b38db3e32910814864fb381ba1e6b50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8ce658bb016e00d54f1a73f11a369089c9725ce41516d9f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22b80d7410ac7b4d4968a44f68f6218e9151129a0e1d76bd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b4dd923ae4839ca6398a87222a4d9f33df8e20a1cb961b88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7541fc198933a40e0b7104ea7498260f4e74b9e18244c602e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e4c47eb67b04f10888dfcf575e59eaf034612b9e957552b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed1e009312c025b7889589a021dd8f3cae7665c33aabe2bce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b335136a18eb88b4bfe99d48a433924bdac908c7142aa566;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb67d7dcc09815195df3f8f22ac49f5472ed492e04c71ae63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0016c4da74fe24e6f786a345a0e66d8fe4659fe18959f6be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96848d6c2a118bc61d47f6e828c4e7f8bb661d7da31c07da0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h441915b651622c44dcb00641b686140a09ed8771648caaf1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h423c67d8aa2fa8b1b5b158fbf223a4a1fd25dfdf056020bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d50ea11a1aab474f32063fbec12ab4b67764e4b2ae11a14f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h401cb5f54981511e5b05ee00423b75ab35462df5041006878;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb2b8a0a4e3d3d0c868e550d03383fd7afaecf8ff73fbd88c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58e9868cf148e99d10eb5c73c72312436fd94edc69f92426b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3990201160510224dcb4f4a77ef06b7816da9ffd01b31925d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb09d7d15c7d9f1a8cc8ead385a7f7218e6b52b802be8b5193;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h720cb738e3e1e5456ff2deecfb233b1b5a1c7dfa5a16410b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf763ab1c1760e67a54bab3714b3616965f60f16a3637488b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ed80ee514ce79e73fd516cccabb288790b74c713bbe8119a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heea0608a985dcc9adefd5523b5eb7a60da781ad637bee3f6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5af35f053670a003558046cd90de94e7d2c526d55eec7b5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3a2e542bb8c3a1fa3a50303de3e150d45c4c9db2d9888790;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf99b466f30493c59610e80018ae6bdc4075a1e3d86761ea8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75a3b7fc38a8bde43e172e469d5291534f49d37b81a864d70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dcea6be13c0db30db36ab07bf05f362c8af4befe63b67beb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7af8bf9c1f17b9550f7f20eae49b119a955dd61cdc9692102;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdab8b2dde5cd84b48d003fcf75dee62b5341fd704c4c394d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57918e29699834e981ef1ac0bc027288a73fa6115be3572d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe6106b26b5e1f6ee9bc31cba9ba27478b116adbc21a75479;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78adffcb0703f1ff49b0d316c86095433ed6a7a824fbeaa61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d84c6c69bf6e4b5195b53019bcbd35f408f43e9ad814e04d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f557a6c4d392cb9396209a1b8e29f9554866ab9743439f8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdde7f785534527b0204e06e75e9a35f8f18a91d7f6ec691b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hced84581d3b073f554fbcdae8636ff0c23bde5ab9ac09e474;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6db7302cc2df0440e04ef0c6465c9c5106ff0f02da03f31b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3088c7aa0d5ff66a8223f1e05613aa07c46957ee2c42c699;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h890956d606f7913e4223cd6419ffe5071ab8fed6521d038e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34a15d38d425ad83c9086537507ded43909a35088f7062b69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4148a4247d2ff7c382665bed7a98543f92b4918cc8e56c2b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c540f02a7589db014301a5237a584cf7bd2b8cf01e06bc7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2ec16db9ebc5ebee41a0835a9ed0ea24e2eaa14f3bfefe9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfa5282b928c0cfb66c4962d21f6c5e462021d79b803ba7bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf41ca030f4e75c5ecd17298b37467fdc8e767b3c25bc210d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8e9be0bf4f5d3a0959daa7e324f604828f84520dfba8e1f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h649ae93134f5c129cc61f221fe9da06e494357f74bb6924df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h803ac107d4bd7579ceb5e5129c1f323e5e69f6d0a62112536;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62684436e1e145e383badbf4817b9a9168a8775adbfdaa535;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f3a848e872507b878e3ceec82b6c8f1244ff862c3ed18c9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63108a6f4fa3c29f9b8bc79825014fb5a96b2f2c14292e0f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16b1a542a5a5089e9c1abd9c97d08a404c64945849cb82ad5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2d1144f5b134069963db19c219470f866a5a0aa2778fd5a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68d64f39709f51c99a969ecba95b0148529008aed45ce8873;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50eb38c2728e42e9e2c007dad4a8fed9466424cbd72c8ca18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7382adb452007ded7c54dee5a6a394750ff2452b1dc922378;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e5cfb38ea7e887b596b7fce6c2e8e980cd9055753c17e296;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd61968801b47bc6123fb019806a85f8ad5a78656b8c5fcfcc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf14c930a817dcdd1f6c08e93f7e58226a5d0682af9d2437d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda374b5fe5b80ab1be75eefd2371cd53af3ff6e354396c464;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h669ea6863e8f9f48bc022914d7f7d3e1f29f9e5bb14b76cd2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7ac65d267097f0d6617697bb41cb62cd9f484425afa4a3b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83931eb6f7ef37d5f7051a3903abe9d4b55a57d3a82a97cac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77442a893c3fcb05b0a9fc6707c9e8559e27d99e212ef248;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd37a3a266d002c172802efaeac266b16063ef5f402f0d5b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b76f9b0bc6dcfd0462fd32aa734cff0d9a7e977f8b36193;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd98d04f098ae9901631c315ef576681384c098078bbea72d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27e4774f9d0356162705057478d4218034edae0c52bd775f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab82a982fe2b6693b2b0f9fed389c50f5ed8b1798468e66f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60b02720f5ed7e09ad38c7284dcbca7d8082e0a5c29023cc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf7c9b8c76dd6447bc06d093017f2c835c0e24d32a77473c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8945d0d467441ca0e26056c1ec7bad3b5b6eaf373724548be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69122621c79dfae32237dde9400e6f120c1a2eb0ff6e02458;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65ddf74bff2fd5ef594c57a70db071864da51b57556a2db94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e7877d22bc4254208e612b6f3d624010c0aac4240dfe7218;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3863fab45f51a2d1251ae00a94b52f0156a89b9b4c77d8f47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ee69b141b0b85783273af95e1cbaf97b750540d315dffd49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79bf3e8d2a070d3f3c8ba871af730c683d5073c8051434e79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd929ed998a587a0450634c65f9b4c2095543fa9c5c0a7fccc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb409f47139fbe827d5b926092384a134d7409263b9fbd765;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f52959af30f7edd108a1b32f54cddf2d6e3dacf89540b027;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ada6d53f22fbbdd8bb5837269e4fd2481717239ab918bce8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5089a13b623105ac57c4ac3b07add7fd7a6ac7af4b9132743;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7a24e814d8fa1cd3f99910fa8a214fcfb9ab6708bea0d519;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1f6079a4410a02049eb46a8ea7e0285da1b8994157afd9e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he195c94bcb1bd097a740efa04d9de9e2a2d0d7a515bb1afe7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d9c3f770eb502d6e0f3deb07f3df6ccba048893781dda681;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6321bf00b24e845ac4f50d7306382cdf9ce02034a36fa95e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4490fa24879f165b5b505d1f338cda9d4a32fb39e2f2958c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd20fd9e18f083e2124689e09a881d80d3559995fe4be45a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98eadd39aa81987b8598d42aaef7b64bef062a6c2a712a259;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h478353acf55b7d1935bcc511989fae905fb75257a40881a84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77fa80d7690ad0b3e94932b0456d6c5aba53758f3de11a62c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19acc4425d726632ea663ec2f210fbe807e19a06e16dd85f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbb1f07dd8331363c686afd7112e713e466d9b3c73bde56b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h606c6b92d0d6ccd2baf682823f48e2c73027ffaad7b700c68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20238e32caff79f6eab1d00b6aeca81942994bf2784b5b54a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4da2faeaadab13977fdf2204a109dbcca8b1b7a40b15572d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5da80ef3b9aa8242b671649a9711f97a70015b8219cdd69ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5996ff81239f9de069569ee9d10a116da8e2c0032fcad65d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h383bc9a44844c505cd51e92e4d8141f8240ce115927759d62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h648d07da1a3e10a9666ccf6866601bd6791b6150cc3d51245;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a42ffa5b9389c925d1a499835b082a5d6cd60b3003e1781;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60acdb1e10aead51e870ad551ba9eab140160fefc131c2755;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a7dfd3e5f0cf97e1bc5fee78dc19092dea994fc325a59fd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2105ff7600781fe4f1d62eb24f29a7fbedd5030395e48b705;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5728468791cf50a51abbeb30646755e895ce0084d6cb580af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43fd1e8e6a7207033ac795816bb3ce326d20467fc2280b04a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf513da39997428cb32b606b26c2059d4c64ee1fb27b193e77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7cb1bbfaf1c3612d03a7e5eb68939108683fa828c18fa1f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde096807b5547e651919e96cf027f1efd638a8fc0f8f9e2c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dd439e89cf7e768b7b64c104cdce3fd24f982b8186fcc8e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfeaeef89467a159ead8ab82ba43e9aca0e9c2afd812fc19d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2471023a1d4e362973e043085fe3650e16c5ac34e9be5ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ede02c7f1f803252f31789749bc79e086434134e17f46523;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f97c5b0a4b6c45e9864ea0b77bb70fe34e4944d35f5c459f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha595405383321294b3b9cf335be619c0445d23c66c400d00d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48979dfb7a000525f1cebd50f7508407fea9a677ccb6bac93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bf064611fdf6b99cede75cc33236357ceecdabc2fb5bd105;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d716f2d5a4ad0c76ab8da9c6271184f3b5d9f2d62b4d8ab6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h712a1b3105b417f6a1114e4d57128eb6ff8796a50941b7e32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb89d99c3feae9301f41d07cc9a290712191a3a9c7af1e18c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3f27b6cffb13d868a8b9a710cce87f56067a01b1f31c147;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d069f1b937b869e3a20628ce8932073fdf4dd1169c70bf4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26cfde60566bb80ee148cd5efd0a11747a30a5fed12f9a284;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2305500c1e4935c006fda5f8686a4ad3c14d372d69bfa29d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbf901742229ebf8c698dc005f506e04db09979f608dcfb26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h507f3a270e2c77f7915fe31f97f2dc6f502fbfb43681aa4ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac853385c88ab64ced9b7c51ebd64287d841ecf42f9d295d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba18dfa57c0ba5f7241cbb9d4665151fe53a1a795ed75a481;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c92fa73e6af6fd5a833892c947bd1d909e7c9d5501e549f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ccaa9a03d1f179a85fe128457e22788c6274e5de5efbc843;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9324e4abddab0201bcfe49d5886ca98efe6078f0f064d087f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee200a4d2eb42af8cea3d371fc555c31433a45d368736a3f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee842864299b25dd3ac96972bb1833601a6c428137f317d67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6197c642a9eec921c9f4cad6df8aed1e69e491abdb838f8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32ae873b62a7d60390b6da3aef486cf36bb804b45f22d4086;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30b7a7a716095b6b17679362b6b5993a33e74b86f9e29febd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2199df3fe3067da9b08a5fe1d4cae2fde821646b8b4f0545;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfc363db974dcad831096fbd05d38b7a3dd77550ae3eeac96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb751ba24d70cb4f128866ff23498e4b63a0b58d53aa6793ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cc316afa9876fac503af78acb697dd3d592614949af67b82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc01c9ec2d2a1d40442bb4b264d5709880c1ffafc36f0a4b44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he836d29a0eeb1df97d09301ccf257f5cf3da323871cc57512;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9470c5293ad853f6022804f8021d522823f2d7de78a43fe2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa034c820913a797add5c886b5bf183cb3d73a7f0c585975b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37bdaa61bf089f59d18ba3c85388d240d029c7a3796d104c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88bb08f87c05555ce3943e18769c76e313f0eacd601986cc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c7b7dd7a72be7cbdbf68fc1805a5fe7cb5b1d0ffdfa58bbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe43ca4a6e8d813de15788f543d948a5cbc81fd4838047b5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h418e968101559627fea53cdeaada5c1193ff546c7ff63657c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h276d9fa2d42b2f854235c9007138a1f14c2a7494e90c18d89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf829303d14fcaec00ed451b4bd1745dcd95908f8de3e37152;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81f4f213d0f156fab070e7720aec29d30c36fec4bc695ee61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha069b0ca86b70ce705427a700151206507f591c2cb383c684;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c6850ae1a7cc29f92fdc9e5ce678270411ae8768b5cef932;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e190ab4bcaaee684ad6519d716ddb96bb5b4790936bebe2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42dc41f1d8017d823a42658dc53c29a878696704446b42c98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe23ee69e4f16514e55ebeb93e11653baa5aeeb126719eedd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e66ca37072639779a058785ed57191622ad8a7e28b4faff0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4195f2b27754a200dabaf40c32ce9b12feca6472c44f019c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6436f5b0f76da53b88da611fc51f1026950b8daa5dc602a6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc55349316dc9c261369d8704e6377077157b10d0a858fd6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h542b42841e8d14606bea398fb92e378f473f8699c2f6b92fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4db61e42cbb4985284b48ba2d127969c5a079ca9eb319cf54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94139c0bb5fee5bf8a1245535433d7bea40b936a1612ff211;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa854d8975a04ba3ca9ff07cdf82563973b0e31a0c81c2122;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61878f2e4aa441f52888daedbf91540edeb0d9cc5d0f4096a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaaf5fba7985d719b51c6da23af75d8fab6389f251b918248;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9317968f0f8ed81d3b78460f62fa5620b4cde5de993f1be78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7d3e3123c23540ed225c7e07f2e4c0ae26ec5baadf968147;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94fc2d1598bd3c5b9282aee393539ef4a7ee6972d4f55600a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58efb9a5d09dcdc62066f03b88a9a98af525286c6aa7fc93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1727a517d960c5d3398692e6d3b32d8391369b0830b7d590b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7498dfabe32c86c56db08ed32f7272ab8f3473b4d7d517e78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b579e24b58e830ce4f10638d038cc0c7dbed2fa100b4a89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e8b39e46a73f869cc09717f0411f86368e8f13863ffa0534;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4508bedd22464150650cb2ada95a44c69ab443325a71fbd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b2c1031f00b4c12dd759d789809e128fb68dc6c9a8cef248;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he55607aa8bc5a8e99c1113af9277a6fbf1a8fca366c7d0ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7134bff669b71bbd79fee2edd0658fc3b6d45247d9aee3534;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h608d79a0a188c426f00f230d459827bf1e92903960353aaa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ec6854bba2d03a9d80b692c65a48ccc509b8b2d98213e89d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he225343abc158641ac4e7d4f48ea34441d032e1f7247f24f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd801e43ce978c4b9bd7bd053abda421aff19aba22d7cd44ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1234655905a8caaee6c904ae657fd48ff0d01a21367e5ecaa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fdaca7722bf1721218010f590d054e886d5935120360e9b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1fa547069dbc393d58f65bada772290a004459dc462fff2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebaf8a98062a255e98750ee83b4503ba2fdf7a1276d90c703;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a8c0245c312c56ccc9bd026d0c7a950c8e68954d583bb231;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a33c3412de44ef9f07b07bbc4ee078ca1fe7c5bca6f0eb70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47e856697d6beafd650be1f13c7d547f8b41f04fca7df7912;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53dd32104878ca772c6386784a64452867639217eb8a0e9c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16e791cf4903e19e451dc50e08364c8d8e9e729d0cbfcfeef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30bb46dd5a82acdcff487b7c1e1b52a0e02873a3e6eb60bad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b8e5b123cb19d561e39787a807e8847a8a2780767b22624f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heca9a4056f3b7d9f1837cd3d810fbda0e6c4c803220302bca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h267f0ec34acda200791c0b55fb498744ce1ce48d32f91872f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef49e80957177768a5e19f1ae780052419ed15953202bee45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc9469e5c7d95996d5732aab78183eabe4e5e2ae0730e8888;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10e7e3732eb278c7969183232fcb0057d82554b99e898b685;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac0812978dc5545adaae310db505d358e419cc7ebaf58d5ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haeebc3d2e4e2a1c4b3b07009b34631c3f68b5699049fdda40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33138708a29a2b098d163042131bce2c909fca1db378b3368;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ea086ea494078df7f924c35d36565b8d927129388f00ec0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb62ac65c08d401e2d54a8acb8fff5f196b064a5c3fa532147;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52f5488e2a3b5d29e7acdf8a1b0182cfaebd1e15898e70982;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha13a1a42c305c642d6068c07eafe3e0bd5cb286bcaed858f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded2e199d3cabbd8d783ef6f0da8708cee498d62dcac0ecb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15e1cb97b2532858d10ac32479f68403bc734cd3e253631fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5da1554e84c040ac6d0569c43309ed14b89c535f92225c4a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3202404047942e933e91eacbba7880bb03f8040f87e95a02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa7fe27c9cf1851b8281a975d5066e84ad6587f5512b3ae7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b0254be9002f3207342fdf0a9958e6361592fa4c306640ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h707d2da66dbd4e6219e132911c28b5a6eb2c051f333c59ee5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he034c79315b2b8e8b9fdb5cdd7b7654e35342a60ad11d5885;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha157d2d7ff29c369b71ae8dde2d6ab1efe8539d834a0773d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c5518dfaf513e27e8dfb87d4595c99e046b9cca65b23456;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf509162e8cf942adde8ea0890ae537eebdc13c1f98423dfc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb2988fe8af391ee9014f4c7076548e3ccff48fd856d3bbf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h382a7b73f52b0eab11afe6821d22c6c466e526df1616c282a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h596e59d5b4862ba928c83adfe4972ca5ee878c6c0de169302;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57f7d7175d81f92796f7f8e08749d9e38c1043a3de4ca2abf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h131205a8d21b07082c09a7127c9c4ad361c390dff84030c07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94f01b10a644a62d523623c73d56f349edcf5e51f94784f7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf56c8be3b03ee77a939b4f04d4b4c9c388263d59829aa10d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fd8d3057e0b0ab4c7f20be670339566d03d64f23722dace7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f3fb08c0bf6eee4221779675d3a0f63a3a96c91a6258d43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fca37109641410092780365b955ade2bb669e33aca407860;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd5ec52e23a83d5e1fddf4ed39e061d20dc57340de99f31f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cc764559836ef25c80c4444cc264f776c6ebbf3a2e6a4c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cf3153e424e6fbe6135e68530eb4da4b1b1b0264f1da3d63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha960bde50eb253c27cb06f3c96b894832b7cbff5c7ce73886;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0e4bbcf9a314506fd097fece71eb6f8bcb7efe9217a9227;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d6e8ab5d8ebaf545fb48c2505b060ee66db0223f4e44d39a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h496134cc0e4b8ae90c080b751ff80599332a237a2ff472ee9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4a6a8b6dcc4a31cdbb8b02f90ea40b9b4b1265a57c5350bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h652174c5ad0cbf3ee0345b90946ed4b5f7f6df0a93bec03ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2af7c074612bceb7bca2aac930cb33416c5ff3cf1723dff7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c79474a5d1941c08a9dee589a0586f1249ab2b95b8034aba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h933086d0c3fc0088431bd5e86cd3bf12f804de72e00d7a773;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f0cac3dcea06a738ee40fcdf66faa196d566630d7d4c7802;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h429e1dbe3040891aa5e83f6e9dc1a58593d5938f70041e257;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he69bf2ab0771c161bcb69f980f82f49e53708e460d9b43036;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebd473e4600c81c87516178a3a30a723c15a0c414f9c42b2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38be30f89798e70a8e2b154b474685477c19e0e92c6ea9b0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95a6dee235da3e987031dd2f4361e20b7b2e5583d29a1c158;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16a8badb490b5b042f59bccb4aa0d4f1b55140178805b0560;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34ca08cbbd13b865be0d00168cb1c65b6e53cb30f08f1103d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7dd12b08aa04d22bc4c9d3f9381051874b90c48dbfa4977e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79b87d3a068ec7d099d5d35ab57f92d68f6b25aca43507bd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f440d2842eb719b5d0f8471f191ff005b3f01cc85efa2a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f2d506950451a33b12a6ec058d73ed1f87d7cc498f743aa6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h563e159bb856e6dc2ddbc2b64260cfecde8b0481f8e72ef17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b0a32879be83c4b43e252ad70c8efb38a750ba7a9d8ef40a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e545bf547593634af4d6bca9919c19958616051e28db919d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea16865c53d721a1cc6f86f69011a264b59af705b9fe0218c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd541cb37197ecd9e9bf9c4a5c2ec7d5398b7b42e40e20b60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c955e3f8fbfa76d38f9ace34ad551cf3d0fc6d927e6170d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99e601849ac5385c43e9165de167ea80aa2967b900b6dc694;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba4eb2f83a27eb9c5836888bbfb20258fc368b9707c623010;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heba5964b0f0dcf02a797192109314a2df60f64c304cf7269d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9688d02700967b8b7d73aa581264b191d1b3a19e84d22a322;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6925fb86ad64722dc9043058adc4812f4cd59a44fbd235ef3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0531ba88c17ea3bd97eeae9ad1f9693b912843b6111aeec0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bbd2ed4f21bb34d42fbacfe824e49debe53440e0eb2eb3b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1351d9e2d891b488f6470668996ab01d64881b6a5c7630c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9627221049e26f726891b59645de986ad39465354dc9c1708;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf8c4c1ca95ab695a57eafe6e341382bac1690a211cca48fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha30a5c1457c0368c4e22861883ee8a1a89796080ecfeb3bef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he09e64b7cfdf6caa0868bfb9b87104fb6cd9f5d9e80733e2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6f1e7a1052afd9005e54eb546dc18e41fa597d1643eaa507;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d03e36ecbf1ea713a4459340f63b8255213638c40b2a31e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc33c22ed19a6e13b06c0a99bed87ffef0826a4c3743beb702;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b02a538d7ab28efc4784df9c29e40554cd655b7dd9191be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98f0863c7db51e0e40453d721b90bb3580a56344ef482f3e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70963c81565650542cd3fbbf240ced37675376ad7f35276b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1376273a7c1e03a901fed8814596cd87739de5cdceac08a50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h815d58ac76cc5fb7ad3f299b607bc20e1f6a3bc571106aa4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17723cd61ec731ca4d2868a89161ad99381c7fad121fee807;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebf859ba42786a99dae9e1b42ea64ee3837ea5ee8faa54197;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29cf2feafed23652ccd621de52774450caec0b6a6665b779b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f685c420ada59d7186364725e15b45c276de5640d20319ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53e2797840802e3d40bc8089e845a9eb06882b8241808ff81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfc2958cdc415449271002dd27b2490cdad17b15d3ac4ff41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51f9bf045b186e38a767b534fff7ca6c45abbdb3d90af2208;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b6a9b3c37de23c4f20b3dc81538e66b58987cbe164bcd613;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc434ca17869e9c3cae3c0cab053a08244e020304c69c6c0cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e0a4c5744a6724f5545b02e1069c1da6c50c0f338277f712;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9967d55ce0b1d37064c44776a99d53bcdcce7b57fad9abd07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h813562d8a7612d1aa9fed41f2d0fb38b8b37161d0dd6fcd1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb337c947e25112760b8a0a418933936fe56ab5328d9f33fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76a35e5c36a14b279d569d2ff2b4d40d6f0371f3ecfe9f164;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c168be38598f9816ee55ef01ce05a5f00d59bb17fa748f90;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fb92fc9799ca755a548f2f2791f0956c7aa3a43264c14b08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4946c1b6b044c692907bb67d37a5cc06e72d26d6461257fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he41e7d6c9ce3df3bcf381878cbf35e9fcdd9cd72a2ecc37a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70cb7514219c087f3c9180db677b01fe3c51b76aa2234ada6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9776c8f8b376d3068393163b41720648397f34b82af9778a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dcef4c62023eaec28c5900fb14b703395270990beedb97a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65afcbb2cb7d1fc3b2570d2c53f347f08cbe4edec7a08f42f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he53a889e1c193c4b20cdd85cb12cc30180dd4ec733fdb9657;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h582fca5a952052965e15e2706d96f651687958304a11d52dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h528b062f2c6edd7d46474ccfb1cbc4b96dc01e33dc944f948;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecaf99acd14bb5b3c1db2307f5a159ab4ed0cb20e49ae702e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76944358f5e02f88eaa7f48c44b751726a1ac0a723dd1318a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e375ba4e84504ae8e2cf9c23bd0f54f6df2bbafeb34d3f41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h424d23c5e0897877be2f1480d311335120ca2797219d8aaae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90d25f69340477c1f0622713a4f38e011a38ee94ff096e8b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66d265f6abbddc6a2c7b50f3e417588e0d5ceca3859c6372f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6cf1f0411deb9bc7aeecdeeb2081c4a66211dc996c178001;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d30847fd0b6d436017c916e67e269621733ff97c4ccbe6c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he17c63ab5a597d6a735d41876a5db183842821a690c313de4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52d910ad8eb76accd4d5393ba43305c46838956784cf7f6d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5637bcdecfb2eb723948788d475ff9ff6c5275494675a0f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb52dce56d9893159996621cfa38a83c67173f182776a11e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81e9a9e497b37e18ac3a2612270e6215b709a7435e93fb96b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4317ce9b0be21f24d63a7a44af7bec886ccb633df82fe89d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9edef200d09506bcf13da176b3293250494c9aa50c2f15146;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b826a57e15352c865cc883481e79f282c96216870c5544f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa455106ab9e55bec8d435226233fc900af05df3c5e8ac07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65c4a842e1a9e3a4d60e467afa7fc27367cc9f2def8696f57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha12f223542684fbac15d5f268a540b51902cc883348e06daa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd81d8bc985b0f7cb2cc61ef852d285bc1f6684dbea25f1d5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8d6943ef383e2f9a96277263d205afe3aada3bed853aef26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h405d74dfa41f1800c38888a47ac361deac1d7e9cf47a03b43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94782e7f1c7483c598c829c41a418994f052250c2a1195d88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4da7af9eb61642ac3afa71f8d43dd54de64980b47bdf0fd6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h514d20e77abc061a615854431c9d727d95a6ee67bdec58368;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e636006b29b9fa39b3ee43ff84ac1ce78c506b6c7ac3971c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb76da2e662478cb775c47e15016dab880611a352c30695f92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd0aac038b9ef7123017e82defb4b9715a157a4af67d5d8ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec6b1c944644936f57d6a80c131b73cd60fd9eac32ce28bb4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2eb190351543fa73d4ab8a0a4dd83ec5a16c860aec474305d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c135758795edc68befc610b091d07e9c9a973a0d836327d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b45de3bf3ffb4c038b22c23917e71ed43ad334857a5b6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc325afb27255f21637410dd01549650874330414fae67fa6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3c175a5f6e186d1b58dd53383e2249f69f329ae5b72d5374;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0a68a8426ec6e13924d16f194ee9ab8f41786daec9380f47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded299a5ac12b0bf55eaa3f1ba9135ede50fb081c71cab1e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf576e9b700bfc6dc302d9d0f43ef3cefb9f248d91a9cb62fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f68df517e24eec994994b934f6d19739efaffb2a80b629e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f61865c0ed3f3865ee075a99d3db69427b85fd8e9a907c9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1312da92259964360155f8e653276ea7b51b4d39f37b78025;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha93ef08cb751c873ee10eb73014b0c12dfe39e42c12df7b6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3214ce52f959d7058191222236ed19916f90cf242040ea19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41793f429bbde61e9e1ae55efa678a7407bc62c88cc898eef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb5c756f47c6e7413937b4b661f1dbe9aa218d266811f8eea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfe6d9ee0b4daa9d97b793addb59cb240533fbe89efc92610;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d94d510b7d8b7d0a1bf1abf63f4c0e6472a410d8d9fe5166;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7dcc33d4e3ebd24978716faf1e5e9dbc7431507beb58e988;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47015c89a4025d3992b0e704ef09dfd37e5e185735d37b478;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he687e856723c73f7090b026e4a3d12b03e0b7b39b5c2d44e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47b676480742d39509865ba664966c17243c438cd262b574f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d7df1abeabdec028d8eb6a62474eaab1507fc1302085c1e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff55212eaf90395e5c2a05ca86d1f551105b1772b689f7aa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cd404468425d752e0379f6fa5f2a4126dcde9ac37abfae06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a138f363d3393953252742eb7cebd50a5be38f6b05d82b00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5786027ef1c0f1a4b43ac0e56c46fb5a0314489d3ffc357e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b88192ef68f3626101d00ae2b1d8e6dabac3a90858bcb942;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3c06c7eeddc61893e52a6397e5852ffe42bba35e038c7c94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23b1a3936948bf953714ec67714dc856e9b582d09f8b61725;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcbd40c50aaee8704224f2ca2fa15c738632670a51c91515c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85428c73b750493713972747ae6ebf8797e2c2ef9b0174e3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87f08ab818c86be2e910e3dac7f359d21ddd6cc62dd98f9e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h896792607f9a80b9bfe902d2867ec113d677abe356c63aa11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f2367573473e9cef8d64031a98e3b8b35f729d444b4da1c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c22a8cc8adbca9a95fd551f6011558c9831b6b68d0393be3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbec5035a1735d903f152682cff5ca07a9ce5dbfc05c635641;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde3fad668dc6c8531282aa69bb584198f538d23efc5175a3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he98feaf5a78371c04242479c53e21a5f428cdbf313acaeb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4993fcaa73ab0f1935eb89c2f0aa8d04d1c65cc0b24cffd03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffd83dcebad52713eed85febf0b6458e3e3f933aba2e5e77d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3561a14933ba5e5edb753104f4745102916ea6aaf21c90a80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc27e3434d626ee026a32ea5a0a923c5c7638ed5dfcab6857;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64905fff0c44463ba9135c62591778e9969e7bdad70add56f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8594f2b9a7469bb4540e24d4d62f794afdd4ad38576553440;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1297c924d9dfd29c5c232cb61b00d162d73aa9ac0f432b86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7be416aa3fbe75be8797939d7d8a2e4cb328fd8ae8e8400a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha25aef1810087a0939793185f2b760b44d4fff52bff02880f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5ce5d2061d9af6344fea25532b80d70d8f975e5684d90c5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45ba5daed65fe57871a5dc42b51b1da41195abfa904913045;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31bbf73a124bcffe62be8664b03c458e9865e962f382c3722;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h110106e899d54cb23e164f757300da567fa785d7628bd7390;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f3b4dc99207c9df29c345567ecbea97917e3a1cc5bba714f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea0110682d8fe6898c793cf8379c2753589d7ef4939273ef0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bd0b1bd81ed961c3dcef68f7d96fe65548bfac9a361c56b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd01747e18733fed519988ad89cdbbee000b0029b5d5e950a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12e6ae956a22d249df9ddb3643b54f622b203469085c7b26a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e386a44688907b7f9766c5b39e7dc3124a7dc8acf9f95cc9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea6cabeec4e08815e22df08089d4f144266169d4075adaf96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd113ec5f76cdd9e815ed0aa5e19cebe5943f4c23d34629bde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdddc10de278cd4b20a780ce7c245fed227d3fe0d99a4954e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2ef0d7d012107e16930975e802bc76229c8d8335ebb67a79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fd01d80b49e1e8f240bb59fb13a687ea6c065fe33b3d1c35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ed22ba80cb4a3cc5690b119dd4922c941943e7a4a4b6e2f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h293b619a78190a32f10390300be7ddc8f29ca38c542218e64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h800943b771787a3333d5e16ec4e40ce9b4f2daced5ae8937a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9685e61a3b5179d0bf92f23ab3580e65b25bf87d132c7504;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd90046904c3336e79d0f7e266a639ac233eda970769f3df6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dbbf8a89de13fd6e5087328818c873b475577a56e89988f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h756ce260eb1c70fde56322cefddd6dd3d1511b9dd0005d72d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb630e92b4ae95b522545d13ff31c7c3cca207baac7891bfa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fb810d41ac3945f83c2c758392081a9becd11df471011e81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2074580bdb6352cf4c7235341796d96bd6d0e8e4aae33532d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd9376a5cdf1113087c6807791395a02bb780f769bdfce5ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7395d2cc6fc6fd1f38a9b75e44bfac6162616e50ba716a3a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc10b34c3e6c7f98f8831b7b777ea574d20b2da07376231fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he12a5e1a290d7a10c21e111235c5512c86aa2a7c1aa5e3ef3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda6bdfa222ef73c8cddb5ed915bd39c8b8ecd469a07ea6e00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7809c180799c0126f16007f33d161140e21c210999676e57d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cb004636850aa8f475a84537946a917be58c0ef1eac75c67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f4f368a7fc154087028e0695503380325716e98e39117ffa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h917f103c44eb0b644241bcebfacd45d34ea7914f03a978b2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he607f7379f29718c7e3409b3e431a123dd39f205d4ec179a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2ad97958500584682b3d04435ce5f0f1d628f53af432965b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5343927cf2cf548b8fd883a6d00ce44562e0541768c039f75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32896cf824972614ea47cf519c0651d2d78b3e9c2ad143e19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27110081ab879711f719361fae89fd6f9f7befe59a7b9f450;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcdc4f235cdc0480037be5ef49cedfec3cac02f00de11edf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc79196332ed71ef2fffe1e3ab5772e57c7d04b00043cb59c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e1c6245c31f2e7496de4298eb58cdbb087edb3b05d668ccc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc7f114a6f36d5acd64c3e2cfda3ede75d61084abfa7d35c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h986a01140238218d568165c30c4a166651266a947718e488c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h312fefabbc6068dc8ac748f9afce00e0092e631f48b6bb8e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32b64fffb0b97f38596543c829e83165c671cc1ac970588a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbeefdcfbd0e9b95237fbdbea772cd8be815fe996b9b0ba97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5ac50b387c7643bb26dc42a475d319e49ab18a53976184b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9aa3d64fcfa87f131df20bc8570e88914b7ecb01ab9a6647;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96d268e430826759b4444f4fcc5c1a9f6372ff5b62874628b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1d88e6beae3595d3ec1c1f802a38754b51c9368479b60b7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfb61753039bf0c6bf013dbf34198c620cf332e60a0ad04d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd76afadb4c7dcc1bbc26847127ae34306a25f9e9d692e2fa5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfde92aad481d070c82b9b66c5bb0ac00ecacb4113fc150663;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a14ee24538db1a2cc2deddd14aed4d5806bb3f2cc3ef6b5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h933d4971d37d8d7895d652af2d4ba0d286bb508c14593b275;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbb67c9cec74f25b519a549e41bae520608fd837fbe626ddb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15873a9b3f0304c28670da49438697a0e13ad5c9c7bec9593;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57960c7df13433268460d67f154afdee5e0aa540ccec83434;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h140116bc106b5474e262b2c75158e168daaba703f4c1559df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dd6cdd5f348a211da1356ba443e6664d08120ff05e32cbfa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4418bc9a4194faae2c4ce66be57219e92594b43bc162bef1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9682fed19ffe86967754ca9c70721d19a57b6ff97d15ec1e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h657a9c1cc51d640f6815c9f68858b8f40854614e78231d3f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d5d16e55871d635b90cf9c1dcfc59dbe4763b01c02a7cdb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b3ffd5072f9f72fa2bb0a9e3a61040beb5ab5beefcc14dd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3a21ec5c59e8ed0b2f7ece46af6d2474a1785e6f81e7c77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75041ffafb36d6b174e294a629d7ed09c0ff2340e77c58b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h235a5330658e5d01ddd3fa9b321d97eb27bb4f483b1d64866;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cdf120604b2a05fde9c6d0d373afa9f1723a7e7365e4289c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2a61ed0bc1240f1f1764be99f13f577a4380c9fc93b8c661;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14474ef41138b2abae01552d5039a11979c2278527f608f1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fbb2b56375806b7b3355f072b69ab4ba06bbe9c6d38fcdbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86690f0a31d5c2a2a157e157463c4921104ecfbc618821122;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83cb683e5746026c65c08560c6b350c6d222d5fac61848c9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc00dd0710c6903461b18fab56fe916dea417a94560cbf57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65078f2f393c23cd88bf63a8d88aac4c11c3acab51bf8bcdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a02b76e97b3758e1d47ea17873b3898660c58b0c02861e95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa342a2d7fd692a9da0cf721b138808ddc5d59974c192e02e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a78e47b61beb1671449c441c2e9c43c24387c3fff5c5fffe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83c6cf13d1ebf93a0e5ad427bfe920d21f6438444d46082e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1227075f27b4c7538b0a0b100d658f30e77fe8fcffd5b2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd864f291f0ed159f46d09a68dca8d1a99b2759005189feaa1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf570a4c2d8a280c189be394f464e04d67d0f09afa151823f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44b944a269fdaa7cb1cc526410789d58e22d07fee1051b435;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ded3e63b7823db8e6b7574113580f4e979120f893c2aada9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e15bea6f8638604a99410c3b6ecbef93b7e2f764d76dcfbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21f1c7f9649f4a8a3d70677711e1bf3423517fa470f53c4cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c7864d99ed7faa15cf3a070bebec547123467d0179f369f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9e654bb82f7813a5889e006baa8e3c9ed4073d7ba1b53582;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h810b88afed89aa32ca8249eff7c5cabcc58c37fa4929f21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h825795f670b4c4d3a8525cc3be92f0dcc2f3664d97b223490;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebc991bce6cf9fd0cf95bf0afa8ff47a202b91d6e6588639d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2f9c3bfdb278304d4474e4805eccb90a564ac9ad20e995f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h228aeb495e1531cea2bcdd385df9fd7c9bec712e1475ecadc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he61a1788b9acf49c2a9d1b33f69c1a442b48618795c7f5a92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33aa6919ed9bace2247fae7fc5a7c01bbdd2eedb47a699aef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ded57f044743f68c1903c5f51fd2524e1f8df81fdbf8570f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c44470e48a4c0b1d6c2f7bdfd9197791db67ac4ad668f9b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc943ffd621752009e014ceec89bf63d44838a70b31056bdf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f7343984f031e3f4ca3a326ac1a526d0c52255a09ce3cd39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha03809a294477031f83d04e4c457948ec3c9e92a7191586da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a12e08440670554983b7c6107cbcd91557459926604581c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda5234f27ee143f995dc40b32f2d493ba82254aa08e9b0451;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b4dc4061971584f17450d586267f95dadee227ca8d184348;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1e97a7377ef813933db30d9d5aea29a46ccdb633882f209e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cc2ac806fe023a71a2df5076fb20303d32c87193d5ae3cd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcea6ba1bc3cfc3286826ac363016141c2ea58495b1dc8973;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2687003263f5af1546e58bd93b09c2167d0b8bde33ffdf71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b71445de7d01186b7bd553dc663932a731b5b81b01ce97a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heeaeaab0d616226b7ae6591902c6f3415f4c655acc876b56e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h916c12798c4cf3ee0dc4446bddbc103a44607a6a54820220c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde8f4294d69d9852b2d2a17ab0da9c584f987d222d5c07d33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d78f022116a1577ad919c7bb953e9ba2c2eaa8814ec2bc1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e4f1b3ada430cc12dcbc7c30bc601dc0c48b6b79ec09eb2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e075095f3cdc6b52e3e36c48f2063fbb46ae2a6c5fcef09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba4f5200c7f4f689c0204de92104336ad8cbd6741b953435f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha14a20210bc1913a6db82846dc26def9c85d71f62fd24fa18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6841b5c1d756302b37ace0932a2a66293056156277132aae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbff7f916b2944456b63d341bc1d52f3c61182a91527c33111;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha52a1cd24ce45761cf387367da5661e1761645f3f152d79f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haea197fd34f74e65ac1ba593e868c612eee9eb326b9b2219b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb953a29c22574f756cf1c484147489218e951c9c4e6fffad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha65378762686857a4a18ddb79c168e88099ccb7fc0536a865;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d561d251f897e6d970ef99e95d5aa153d7fbb44ea77f75bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95d2ea7d15b44d4476df19bdd6a5d3ff4c83e328452c4bf2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79503e76176cfe7fb3b1c35e1a5f352530eeddce4a33acce3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5b1ee1be14dd6ee5ddbf2901c4b95e35401480049729a37d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f19a71365c594075b26b5c8db7f13d310ccc7d26801944f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e18ea69d04c35decc687b7259c0170286261b5b1109223bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f8c2e25cdd4cdc083403e175f7f30dbc46eca82632fc6b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf07e59e7181b9e1d47ad68d126433a54ad946de8145f02cf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eabf36be4b2a256b03100645909d448ca670b5034598fd2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfce3b3b9cb4298a79bffdec4fa1b7f8f51a380fc359cc6f1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef18375fe0295b65fbb17c7fe0ab16b0c6a6f8f7a5cc49ccc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he08f7ff0b039df6b37ea2b3be3df0e90f3537a7fb0d06a064;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7236b49e6087c0d3ce6e2c4a073fb439cc0ec6031e19faca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4f04219353ca23ac80239ec4e550d50afd4c2c77729f8126;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ad0c03c736a8f41ca791af4a93a287623e63a60b717b25c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b7c05d9bc8babd10d53bf54ae886da62c794f381fbd39e92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h703e0d696e79f9b02bbeffc45fb5156e5187bd83e5a557598;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb62f68ce351022d9ff6e5cf15c4d770516535721308e45463;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c922f0ab0aa7fed9d068436ef18efc033fa86a1dd9c8577f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c5e1290f6fe8ff42f8797bc786610ad29063fe4782738226;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1d3e6c3961d397023ffdab2c315a1049e5c491c549d28252;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedff0443494ee708025d28293cabf8171659e9543d66b0c35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h952b32bd8d36e3ddb90321c7468d6e6d2672fa06a303b17e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he222d7708d8864c485d201cffcf2dcf15618f16cfe6ce2f59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafa2293e95fa088c18f58638c81caffe535c3d4c9ce1a9ddb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf17ec58196979be917a9212aa0d3d045088daad71a6094c82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he939deb6938f6cf8ca595d823f31962fd466b54dfe26009e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9887fee0ca955b4dd9c62d8205d2ba76649daacf157ef994;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9b8695527c9f8bf0ca3dde67969464eb6195d584d2f7329b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3970a1ef07eb97851aeb41d542c6765cbc00e4eac5ab589a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71a1994a5d929570a390a9050d5c56962a5383e6825299dd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc42fbad8d3cfe50475028741af19b9d503e66d7c8a92d331;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb206b756b49916fb0e10d8e7ef59a2e47e04f727f258c0e1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h479f20678fdc54ffdc71cfc5810b05147d36aed3e63c69220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfaec5d47741ec79b01344aa0086b82a93d69530fdda1b0092;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfcc36b7cc1ad58b238229e5a0514eb4852d499ac7da47387;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ce7c08c848250d54d2bac173b6c888796bb040def91802db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb1e6b48e09cd614a11a3a6d36a57788b62da05395da37a6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8f54f912f4a4320b371c5bd599773772bcfef8df6f749972;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f693c2432061952079a614591eb2be907008bc16f60f3551;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd41dc02e3bc08fa30f5241642f0994d05e24cd9f8c5c4dd78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22f1db4eb829f11690ca68fa91b4e57e0d73fd72edd477b5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb4767819275eaedc87816bc0d54c43132a1f90d229f8a791;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h322e840390de43a6e144938146b9888f4de81f543608944aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe8ddad930350f97449a6102bec666f47909c8894748c42ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bf95194e077b50a31818e1e0dbbbe970dd35ca6883745fd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fb4e8476daa0380fefeb21daa50e4ce1cc75960d50c03edc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h147e2379a925277886520595869e2ecd31e291dc15255ff25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h287eb1e6e9964d3e953dda0cf883ff2ae801288ed96586843;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h594916e02abf8feb0d72615f3265bafb7aa1f42ac97081c10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5d1bb81b83afda3177d6118e734ed8e4ccc9ececd60faafb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7a1b02ff9e4fcb81bad3a7d51b19116ac5220c25e6c4a92a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf74677ec9d8afafeca3319d682d97f35b69d1a663888374aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha478da79157d4cb1eebb72553f08d2fd37f0f71249a4ffa0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf996ed92e15ecc2dd51911bda5f591edc6baf30e68a0c4c4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46085cc29b52ae48f3850a0fbcffb0f44ce51f9199e1caa10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h324a18cdf81af49c516a640153ba8d269eee974bfa8fddb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9d0d65e2f95c410e0c3c96b878e64df36f237118968f9e0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c458e55b6dd0d34e18a4c59a00d993db902ecb9d56c7f0eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78c594bd924087270664a203ac127c6462a734a15d872b52d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ddfcaf5cf2b6db2a1e4a489c8595d98751bc076b4f5873d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h116776914be351721cb4fd2d160c0700a8bef0bb6dd3fbe60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2596474b5143362126759753a99581000a1b3fbcc9ad25220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bf1b5437a83b241f40ab662025cdd8bd1c40fe7ee26bbe8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4043a85e34213825f8ecf132655e90793fe1b193c07d57830;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he36d2c18c40516fc2c97cbb2f59f40e9f1c84e5438ec07094;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb0ce621900be2b23d3624260e7408b43344f2e6586c318cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea69452a3e4bb93d74b9e96a33caff19a4c1cd75089a1ed4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75a0083372c7f9c297bfc6b425521e49d39dbbe44de82cb99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b81cdefa1e1de06b2cbba95029e12e3bd4e48c276c438a7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82b6d170478e0db3d79f8a5f5af571a14ecaec279d5b8b508;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f04b771edf438f9c0279a7e72a3aa50a0f080481b652c83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98bf8f7cb054aa3834f46e9668954f72e33428b71cc43fef9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6da239540463866af00fc2317feeef6b2734dcc3229ccb3b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b9d17fc237f5f2c4030ac1761ff909868f257edf9dc02724;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80bd28c038f2e08e5093aea225a08ba41ba5d9e2cba1c513f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6aa2a509c33fbcc4369ed71e615bb431e7611a013cc40184;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h165fc035126353f7819ae62da8f4c58c5a70aa6e3300fcc55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbb1d1d94da8a8cc51f278934d6e4b3649e79cec842564b7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b9f145e4ba924e5acc0abc77ae96561e1581dc037027c1bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha26fe7578e922aadb3b25be0f843c237f5d85cbb80d28c705;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e3fb91d07d89435ebc3a34604008843704a4eec2ac2a212;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc46c2896143e384a80f4301ff2e84746c6f76ad9d30092839;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ce464297672e97e1c764469bb4aba0662a7b08a24f6d1f14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habea9f59a0c266b5cface2e9231dd6cefad75244dc58becfc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9d73a9c9c89cc6c1e50f023e9e9046a5a5d1da9a02d03079;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bd46294e2aeb394fdb71ea2c9bb386769f5b88125c1962b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb13bf31df4a8c8c20ecc4cd32e2e2ecccc203a6d4f28212ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65fe9ae723e9a5f13ed65893791a09c4e10db1a9ef70b9fe1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f68402f3442afd6fd86c0645984296253a1152aec9b82d87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc25d7c5bf36881f973172e096a12f1db70c1268fcdd3766e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h118c4e03567e161fc1923854590a091dc9622450f13709c7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43c54204223a6e5aa179e4aeb7fd636fda966eb88f310511f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d4c82b2960b8c97ea4804e2cd11fa15c2d461ba69271f5e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a34eabd2883c064e1538755b732466602dea12b293820b76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd4e62962cfc6ec869a614f0603d5f1e35e83208eaf5712e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c8fea7f6a0e77e922a6a60161761ff23590440d546065200;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he26fbdfc5c67cec23650d24064db66e66eb060ae1546fad54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haed14d27a3c0798b306737e6153f5efe697b6e32b59c672d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69c1ff367773793a94c3feb3bbb514ee8c979b5291a3e80ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36b817917da7bc79e80ff0b349202649483fe5cfa9c61ac1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa6608221123692565bf5e8f4b1e3908759ce57a08c5dad7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ed5364dd69486075507bd422a5d922e56dc9f1eed23514bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf051b9225536249a4bdc56db34e6f3d2117128ce371fee19d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc20e5bf01717612b323fe413c871eebf8b84cb1c298e0a17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8062d1f60b925ddf0114ec564180fd36d22d2cae0ad564b56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h396836ab14a1bdec4cedde08d3ab2414e01475ec230d94a15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd3bb5f520f2a43fe732d0a84768eb39669c46e424001cc2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h619bf58e79163760f143e71df4f4b712647b516842f99ee80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbbc7cb0a69cb0383bda7023f622f367f480723df0e04beba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd05b6c4a00cf2b68c1395a593d4d187c696a447846ec0780;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39008c2e8a691f1d38e2f0336c5332a6ed349a454dfcdf858;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4490f664ac46419c91491f7152981293a919bc37e406542c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc90f72792d27f81ecce93dca4a4e7c57c14a402d4fb0c7174;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0319bd61ed086f08e63956bf2e8e338ec3e0d59665f6cc71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e4bce5f5631b08484fc8e7d8a183c5d2fed24943b42772;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4cf3942954116808dc5408948cb65e6b68cc48958b226c86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h944001d49157f7fa26b494a7890a97508a7d65c950a852ace;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he54ee3217f783a0e4cca634cdbd8b00192aee980c63421670;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5be3d31f569e91542c9c08651a2ff7fd6914c7e64913e40c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ce811ae12d1466cc964dbeb9682fc36bcaf87667ec48fd88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habd1f6533d28efca2073090b8e5af73b41c20781262676b9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h708c874ee0fc5394eda7c237338257031033bc02fbca416ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1c091070a2a4c1e6c0084f8b67e9e98dc3e08c548116ae13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0db020127df640356c1b2d6df8c58016103b33ca1c53d9e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha24ece31a33e887cb6d39769b71d4887077fac5d5bc19d832;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had3c9b2c9f589c71ecdd4ab481f995ca1c40eac1b961d3470;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14255fb00a9651c1adcdc7a1b69a1d96cea3fe4f9c5c5b381;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bf251c146f14eb865aa2765576fc2a397a972e1109e26f07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d648416ccccc191ef4dbd3d9222302c247ecbd464352f5c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd059284281508f2d56c6f79232efc7d08ced8483629497251;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb65bea904e3137a14b7acbf71514a3ca35f29f2ca950281ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d4665f3b566572d03459aab3939e9c22cd96368791bd7f76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a4817cb8d155e4e9280bbafd357b3ba50156c69856ea3fda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e45a90fbdf2c5154be6f3997263020917bebb8ca2cf936bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74ed29af3e4eac9bdef9af24c8abb307903bac6114bca1845;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90e0dd96ddf86b32bcfa4801742cc2a1df621f4e5de72dc12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90706b722f4e4861c89bd1af287ab05b3a64fa2b8b260dcb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bd7808d4ef4651ead783545465fac00670c37afcca9e30b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73320abb0837365082ddd373f06fd186ae48ca9fb6f681dcc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadfdfe35700e331783d9713d738db1a102bddcc1df8093ace;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22992088823cdfcc2e4cb46314edb1b9ba585b1fb106d7086;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c9c21c6aaf4044c9d1a5531bd118e9ce29d1408148e70f45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22638ec4042947d82d645e8d63b9db9f6af591d0c75858433;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d382d3b25f1346eb523a5207e96d2b52621c7122e1428a93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb781e0c88cdf63b432ac3e35291bf71f427cd5e1defcbe883;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2fcf1aaafe63f3832fa82d655a250c4595ed6bd30756b806;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he731cac5df8eaed12868167976f08720b084a1fc17e38a77f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a85b6eddc084a3d0e9b453b43ba1eb201c405713d815157e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a963ec4d4b79b90158802d756b69d50edfaea3cadaef08c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe99cfcf49d514fa2ddd61ae842bca3e66bb0f1d0fcf1e134;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec7c6ac6207c65be5fceeeead9e7cb297170782913891c388;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28a32f304d1aeced3b9cb997638fa56f07b675868ad4b1fc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf37ee81bc45285af8b3156bdbb63a08b3c3c8c5471f82ea51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf382c6387f5b4d1c43f732f4f64e580fa86ab9fe30afe5c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had6f031373c4739b04f0c771c6b0984c88b0f5bf7ce28e6e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heabe8ad501e746e66375c6408055281393ada3c940e64e3f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a1788620b01b095d0651f0488369566d6c43f8033bfa4e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d587b414f451abf097413c57375c5b54852eb8a8a951e8ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7633130fe540da6f167bfe0ecc8fc201f55bc24906659d5f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7724c8980371019a7242b1f626313cb08563b96d3817ad279;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb9629139fda8d182e6635c3a3ec93d66f37b86e08390742e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29003370450affbf5bdd8934d8846105b45627450000214a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c9caa7d78730bd1179c01303c9bcd6eb82fbc3a9ac3a2088;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38f7e2af4a0148b0fea68c108394d27f328e52882c6ce510e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5df4c807fb7365ec9e9c867ab1c3572b18c4f5d3321c774d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1d8432d0391f378bc9a1c06b09f0b0d70d61175333ea0d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8dabab9595b5e55019feab9ad89808f2ad3d28e73a6d1b18d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4cf54c7ec7cda2b83da8a4403093bd2ff5aaf55b69d28417;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a02579cab11a60f7d08b2af65df00249f479789187aae0e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13434238d4ce5c1ecc5558baa846dbebf60f5c51754a5ba9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2c86ebd928bda7299bb2e121d41f8eb01908356a306949a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed2c35c53c0494ac2644da8e9628d6a3c3110d48c687fd582;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b613454d99d51b66e1633c374ab511e410bf6de36138ca1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5eed4a0379e44db5f56c4fe72dfe25430b1ddd77794df3e80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h810ca8c6439e9591a7527070d2b3308f265756917cd0672e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc08fe2b7a14de7aba7fb972465ceae3f28af78c5378b3348f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd333a259f49dc6d17c650a0e19ab58b6014e1374409ef1b28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ae81946a6817a27f12377a354e82f8fe0a48d1906f631d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7edb93fc016c04a6dff35381ece957e389e0b4a39b6a5caec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h351b4f4f6be1f2d2b1a24ce7c5064c1ba3f8fd07e3c2b4b8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3108f11565699c4d29d69bfe6b15df5d904c7b0aa6c13767;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc90aa1a2065e689bc34b4dc73841c4adc2d366e22a9b080e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e7a6db5784bedb401de67bb1f6561fea7b5f72d72050aac2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7109983bd4d04b257b009a574be9faa5cc1f880b88fea510;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39c9380a1dd581a51c097b4cda2029b890ff174c4096d5e61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b196b91bc47277a816bc0bb5761b24c7008a986bc469b3c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf71826efb3c3f047db59588df5e659339e7b980e01d862197;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fe941c4f4da0f175bb68697482ca6872b9e3b8c2d71134af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9444839aa65dc7ecd92aa3dff4abc322ff944a8101773879;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82df6cea98493f988119e3627251b36401748af4d968ab353;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fd27fb3d2086f84440593958ff3aa383743a3fe010ac370c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf72266e1e5550048b8f6b870ecd30dd3d8e966a83b14ce91e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55e9e64386a1908d154488a6f1c8938e7e464f5f9d2d701c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6d7b1fb5cc4ef9f5618a62ca376e266c9572c52cb40a2438;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a78dd40c56e744404cb91c4256e1843f87cf50e460d4d74c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b31b34d335150300bc1a7e1ae44c485547248b03e34684b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1eff9c11a36832e3a9ae848dbdfa100715c52e1000dd6422;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49b547a8b254e4e36d949484249b9d836c10b19c813b0b455;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab07266e98de5d12c232169e8bd18036580c0205d9c7e32a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50ef3de778c9617835376d85186bed0ac3490409ccfaf907c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h923682106c0e0f8414b11727f370f70ef8b328740c7680e12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55d4a5b930597a5f8c637359bb5e33515a53825ad7fd7c355;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15abda5df5af39217cc1108208874380aec747ea7beaeecdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52c169cb3865adf9642c3566dfbe7ee812067de07dfeb60d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99c25aabde7b21d4b33765cc88fd98d5dfc56dd8782411a7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea4eef42bfd7c60263cf3d4a839f785f6b719ba0fb2ce0738;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7e025b36f3ca844886a25971213425353290d23c5fe93476;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcf1364fa03d67d4b5d1d22b7e828305eaaac7447866f217b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9a231002360cfa88397a91eee86486a59c5065694a76f6c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1de0eea532402868a9ab13abf206d9cc79dc2cb7c7bbbbd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c63e76d49e66187b0634535d40f79474fea78bfe4d57c0ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heed796619feaa4c67fb0d5ba547057c9ceb55cca5dc08bb9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed93e3b5c406ea4795c0558dbe564148d7e93da231d41a01e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heef133f3e1bbacfcf48354ce2ebee6e0b2eb26360666d35dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45dd987df593a7fa683a04a55f174a469d00f0639540069d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72b38749aee70f1b128d8b25239935031b52ccab3920f96d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb411d62fef06cf1c03866b2a18fd06f45d0115ed5e614775;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6086587142a9e507a30928986c53d9c0fbdbd5e2439ad08c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf060197e40f4518dd82c54dd42feee704db242ea5cd72635;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc2e40f419c726191f1b8f745b8582aa6049426f29cdd6901;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h217926868a6e234ac2917ba38e80d3e23c302b4064ee4ceb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68b78960268a54aeb69ad62b6e260e259e07f1dc4221b3172;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb215efe77556d0e694ceafbe311251be66e611568307348ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24e1d8bd596aa98df057765e02bf661970becf9fa0dc3ee55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34cea7fe3d4082b5daa008aac6f69453dda2aec15aa02251a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53963f1c03312a0d5739ea85709aad9f582355f85eae6cadb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd02b5eb62858334adf7a02c4eb84f38130cdafb7a0345870;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bbb025e7a9698024668ad5849f78e147106d45bdeeba936d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2271f8588b8eebabb6cd527b529270b2df27a1d3eaecbd41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3416c6b05a6856670d2a044cb93af28bd9389fd3c0069a553;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dc054bfdc26519f96eadf389f39e77d7152464ba13270bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h662664885036a8ba59c8cd6a9d810b02c146111e8391f8c61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6032caca017ada0e7d2ea0679d48163bfdfbb3d5dafac20a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he643b44e8bc26acb04eed0b8f5d753b60ad45e6120b3fa3a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf40328b427734429273797fbfd82b88402ca2d33426bfecc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h429d09317c0be206bae6360a2161c29df6226d16a39be396f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h782805c20092e3c1cc484d5241dc175a362b5be02c6a47da3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h386f96bb7c109c128e8fd92c4cfca42f090f9e06660045f05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12e36bee2b50be7640cb894e4edbfea366fcc6f5293239aab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31eba8ecb9016ec1954dda8a0aa972dd2a4b1fae16a0cbe8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55898004e307fbbf05a2c9a8e23dbc452c716775daf58a50d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4dbdb67385184efa29f9c2b93f7390dbdeb9ba8fd4084f73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51685315edbd68c53723e3d8a8de5cef1c70b7225abeef260;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50df51764421f3c3c485355000297ce70e86a136d7c208f25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81cb45b0feec8cf3407ff57293b75b6dccd412817413a683e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedb8b3493739333a1e941f78730c6a36f815009c1638eb6ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e63865467c50630573e9dd05dcc74ddd989fd64617670a2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc819e7e97404c5172be236bb36a071840cfdb823f0ace3ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f645b1e6828f1056540e8e8464d92982d076dfd1b8e61caf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2647e6bd40c8f933c8437bce9fa1593c94a6a74baf4127cea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4953e7a57f1263dd114e29c1727d547fb4a0703a0636473c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7a6a5c4effdf3818fa0aff13265f9836b4c1f22359bd532d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa12e7b367ea99779994473b2d132bf50500ea4005f5a1bc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc06e85c5626420c8b6e4ce3cc6b3cbf26550edace617cd662;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1e7821360bf4c2fbea5c70ef2c8a58efb0da5584173f03e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5975fe568801601b86d01da5a25b3f7856d7bd4f6dac5d34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha418289c4efd1c00411ae5d2b59a90b679dc54474e2b82ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfad2fa5a03296bac7861b3050b7a3e07cba23892fe370ca8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1607455004398f2d7809a563fc1eeff057aea816478de77e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf81232cbc280407808e6e42e4e9de5219a48c1edd87f00660;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1339a2a5530bc4ef9c55eff9176d48b6135a3f1f7fde715fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbae8959a5fb3076ebf1311f6f0efc3e500b8a1dbffb259a19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88c27ed04245b5d68d6d8668c8f598fab520b0db3a8cf1fa2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb705619285b1ecfd5453ea6dcb1e9091ad61577c402060529;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8e86a30d0c056059de6d42520e236556d1abee8ae140257f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ea8ad660885df8908b0f9bdc69062921da22a66df7a0ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfda5a6c41b0ef01ee6b34e3e6facbbba07123d345eb78c98c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb35a6baeca7c919ca8ef01d8e9cacd4a8341c46c6f8b13bbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bd7d2fd4d830556539a0c6685194d1db7f46be6503d519fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa27d6fe36d9212d0a06d3b8b2d689f8ae9a1549a60b76792;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4474f9fff825b8759f31d68690bd19c144a518e642183bfce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c3dadec9dd7bf297fb8e08486b134319636feeae32b853ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdecb5c56fa809df1f466ed0b9e9aedbf9b71a74ac0ce02aa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92a71663f98ca2021147a035eee9daf59356bf2934c998a04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cbaa244f8eae7318a78d095c42e64b9d8bb9bcb0e90df3aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4e4e4c1504f209622e6b6123011324c0a00a64ee7c5df497;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde82e7c3c87cde216ef005ca7967cf37d840a1cfb37f066cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12a77fa7fc942b889fb693669605042aaad61b9ae4c10d29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d20b1bf1a79229dfec0306ccb80cf2f82195525ec49aa1b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8522f45722d7678ddc400cfff6befac29635a64425932e3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69898005bf89be8ecfb25b90f280ba0e8ce5d29264755e4ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69fd70b520f0d34928a182a4d3a77ef97601880a9e532bab9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73a10950a11fdddfcc21c21c1e40e508941ca55474dab8299;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaf9c0923e64d247575bab465e22daf8a87b410e856484bba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7490323b0b75d4c4ccbdbdb033f6a63e4472fcfa6831ebc9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52ec12c268fc7e65f187f4c3a810b0c5f00098c33c8072757;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd495493b6c23a6cd370160afe9376211380ef71c8d5bb2e65;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h582f611336076049c6a695fecbd230ee152f145994967279e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e4e7f4625e38c89718c6e9e94de60650ef59817c93a4c03;
        #1
        $finish();
    end
endmodule
