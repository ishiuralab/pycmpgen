module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h360cd1459aaae5fac0f7e3d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc166aab3f0559b869031d8a61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72b5f04fc2ba54f399ff335f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1ca799168e4b48d6eb329884;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4967a28384fd83f368aea5c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e7d4109593e63ee646a77d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha279db71788f49dc1e32ac50d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h879b57e8b54dab922cfbc71e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7387eb0a495ca4cd9d9319c82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab1aea50941daacde2309786;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84c9a6778ea9eb6bbec0885ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97cef3493c60c323933a3ef32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9c38b36e3eecaf9ae0806ce8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea8a92edae8bc5139b662ca28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha87ab4ace66b835ff822dc60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h407b5a624beeec0a4c0f2c73e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h677837fb6803d1776810e76c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h287115e7d9df966a4e50647fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6aef0f9bb57c6827609a9853e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71fc24d25f35caa5a7424b740;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd073d13ee2a0ee3899b01b58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1a5fd1df09513d136de6b3ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1f2dafb4fa3aaa889ca578b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1396a557327e0cc3886d607;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb1d9bb729537d0afe7732561;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b812f5d0d9c7da690abad1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5492dc500c074560e11b8ee48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bb1da4e226c89ac428dfbfc3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cdb6c44e3ad3e877c87d66cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf44e22d94945b6341c6b6ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha75dc5c50c00839fe83e3b51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h817735577d887c5329ef96f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3682325e6872bbe05d23d417e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24e1d7a96d3ab165d3e556401;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h161884f7f51cea11d6bf6d15e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0f516035c4cc6f70c49cc846;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20efd740485e47c95291cf77d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h884bac417b61ecec5141ffc28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dc1f34777548da37aa703068;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84e6a18a19f093d1d68476f9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ca8f37fa98e74f3a425cbca9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59e171f477edc13684f85cc97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93f8959072bc4a9567c67b842;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h718c273a5e1bd85aa4fbb78dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h948f9bc99f6b84bf8bd1a886d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8053ddf2053814b593e2ebfd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98f96b4faea3e1c1c24f016b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ebbb2208dee02ae177231b73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ffabaaaf678e766848adb449;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2405bc7c66fda222ece96f79c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f2c257a67fcf15ff53b2c402;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf0f1a46185772b4b3422a46f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52ad27275191ccb81b2ac3f3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h762a012f0212975615508bd58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6fe6efec85f9c6bd1566c572;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haac75d8f10d947a9b30ec5075;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf6778d817d8073da3e66dd24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0942dd990580e67ce6def89c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h995959829e8ad57dfdc98dc6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h974f01fc3ea0af6843beb6076;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdebb5412dd876b4c6fd0e8862;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85b3c27a3465cb679ff07b730;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c4731c37aeba55fb400785da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8c9986f098c0818916fe682e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f617c92eb92f87ad7cd82eaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dc400c80cd76beae6df1c312;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h816f8b84eecab6ef85f008bff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdccc1a2582f1fab9a84e6653e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c8845b39256911eb3fa3a650;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bb91c5dccdc73558eeb16691;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9de76cf75dcc33f0f21cc6d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc288a8c4ad45eb7623866dd77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f573b1899ea737802d48af04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc86fd4f58a1ff9e543e75722e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28a395b30cad7263731773e0e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9978080879e222dbdd7621fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab67e894e46900d3fc2b4af06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h816c4e09506e7757288a91b4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22b89e41b3a0539d0944e6b95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dbefa471f99719476cfde351;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f0512c61f4f07a2d7a50d1e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c15a83e510c9aca4190f406;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb30f126f1cb1cb84e5b13c75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9788015ab413eafa38813e087;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h368a87bdff46f7359226072ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb61328a49b085ed99f984dad4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c1fee0a8d24e4a1d54ac9035;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80fbabaf4ff2ddcc0e67e9b98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9640bd134b6f0f65b681ffe2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b72010bfadc721ff111ffa8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71fff5313c2e763e4b393162b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha206361273d084a2c1678ac43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ecdf23afd4f0acd16b0a8263;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbda60354ffc7b99c8f1b2218e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h985c6c626ab9a92d241715aa9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b7b91c3ed8dfaced28ce317d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7955390a9fcdccd4f7b93b89e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67a0af62baa80895b3b72d7bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2160718e6bb72ea83f3918d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b496da457546f40add4fdd05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1fc9c8f212d2aec2c914c645;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0e9a5eac19120f2998368162;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8c72d93b616bfe7ad9d9ad4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h421b70fad3f69d9a139a3138f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14f0993da57fb2ae8de55c506;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb794a7a360e44f0f1ed45c5d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a4a17afb0c0a8709c89d7f87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77305a54af4e24414ee2c2549;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26fc25c968a9b339184cdae5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h683023e9374864058b42a3bbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f065abb599007abba47c4b3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf73af31c0c2346e7b88e03c82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7582ed9a16807f465af817bd3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb29c4c61f2e18c5cd4661834;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63f0bc63e2c3545262e0be14d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bbe7e4c963a745e5e4d4bddf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a9c550f96dfbbcc6c95aacd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc54d9c488fa9fbc66e7a52b14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83b91e32446900ae6bab97101;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62ebdca4803250342cf8d047b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78ef03613f83602f3a2c5e910;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fcc30cfaf3e500383e1c6432;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29666652b7eb486f4d2e22d57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2a5ac8334f9da2027847759d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccd1eea1ed6dd44fac5649756;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa64629e0eab62a3e1fcb575;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1185ddab182dc208eaac453a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb23fc583f8b4eeef6864eba73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f4a977a33d81b5eea2fd17ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h749add7d7416840b2f9162996;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he03290dffd82c1b0ab576a036;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6aa3a5728e631503d0c49f9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a1f3c143c590642c8815a401;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7756fdc98ea9f5ad03aef1a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62e65e79e9ace65d0473ec5c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13d536e38257926a75381db46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fba961242d07df577e13d0ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff4167608bb14d97d97e5b8ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11daff69fe92b65332500c74c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9224d98c4aa34140658352e97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf492bd420837610ae9ed0e42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h270432c365745e7e3d79a5f63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h765731798e86f16446dce3195;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h908b28f676240960012faa743;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9eeda2ec794bdc1ac9b82bb96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb903f5996639d42abc560ed47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2affa5518744b0c9bfef5b850;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he47592ddd017c735bceb244dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf60f2217cfe3c7e7c9ea8d3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b0bdc69b884de0f8e5b73ea6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h214147f2a658f0d4c19fb30ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3515fb9423769b5c8785489cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e5d0ada91e168f9845b71ba6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae80735a4e9584769b0e2b4c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde84d68ceaf6c31aae0be284d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5237e2bbc01b31f2e7946d60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13d57293a3771b1800cfd27d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42896a4cfbac7d956a2101cd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4df842ca78eb3adb4f6acb3af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30b86449185f8501feddba586;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72c3cb5c80415eca9e1d8f91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h427b1d8d61b28f3b558bac691;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8299cac3c19e166ff7764d4ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb04d049bf23f8045a56fa4048;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h353a2367e95a72744892be3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24e4a3fcace3a59cef8177abc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74ef736390ac188387f177b22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h646507a855a711f45d9a23b7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf067828cb9b227142462b4ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed2964489e24479e349bf2220;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0fed4e40150846576602d3d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68f45261d4926da92d96c06b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfd41cd47e919780312b01ee5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6c8ceca3d5fef2b7b2697044;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heafdc334bc138005366a1119b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha506cf1e28a05ace4576dd0b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3390ebc1738dfaf650a79fdfe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95283b430f0bd9f50b16f299b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hced9df7714d011a8e8fadda87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he73c08c4267310c690727750b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dabbcbc00540091b71418fd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcced1d10621fa2cabfa4ed9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c3c6a9acc2e7a494dc6eb251;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h835da06f88a166f275f989621;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab96fc9af9f4f277b4812762;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6c9cf8637786d06113f868f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1f5a9cd9ecd78f71cb72406c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc81c0a3a2be8135cefc83b346;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde79d6f87c5433c31c2a7ebbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61186d806298f3a97dfc31867;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90e5cfad62e06ecd4358843ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a202d8f47e4783a3887e6511;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28eac68d2eba01f637311ba45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b74dde230276fae6d251fc85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22feecb87c82ae763f9f16b89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb1a2438a680c7ed45fae3178;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b52bfc7a364dfc4abee89187;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8208a914279ccb20b5db0fd08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e8f33509732a06bb46de22c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f1055857e42793b177b07558;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97c7ea0c72ca19a6b4f7f2f22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e7ae6932067b1d02cf4b3f91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48ace4d29bc18073b185fa70b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd8c09059c5b4a66d8fde7bcd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da3a445b36b5b0c0ac12fa21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe6c35ac3e863b795f58799b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b76d106c75e22ee101a5b14d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f35d9a590d153ee03ff8b534;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb933caa6127154ac65e24c583;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb37536aa2cee576d16fa94025;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf29a477c5ce40f4847798c51d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1f76820c36580b45cd50edc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79e8fcd1123ca43f8fcb32e1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d1eb6b72ba72dba7d39712ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6603d4d1d250a50f4f28c82e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e1676afe9c804cb32d56793f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57c7a6cb9bab70bdbc798c6ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc04f6a3d62845ed451ab37d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5c946b4e093eb5c807b82f1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7b066f5d3543e9f374c6f79d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69f72aa55ed264d649dbfb489;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf658311bacc227d3d0e40209f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h840e425b0dbcd2ae471c3ac28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e4fc11c30f8290891f504b3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3191a54ecf7c4239a90b10b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29f6878c46c71d1168abae443;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c75f64de693ea5c5a027e06b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h970ae7ca6e81ba7c51df343a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc42c84fb656b5ced13d54a67e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h471c7dd6b98d23df16acf59c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b5b35c3b9ae894e40c0028c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc45c67d07b0f69829b2d91f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71c1d246d16ca8423da2738d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85975aa2ec33f6843f1c13a10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fe9da3a81168650562736578;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae5ecb69625eb6a8598f434d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa27d136022cf36a6622c6349;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54627c295b4ce765dcf1a86fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23aa8405a58d234ce403aaaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fc2ca6dfc28166c0a80cc61b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e677eee004a2bf88063bd714;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15181fb2c588f4aa65af09af1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37f8dc69c0410ca4928c0a2e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1f09dd85d0ce25a9824af422;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9160fc33b48227014d529795;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ac678c216c01b5397792b396;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb13a5324f97392ee5d9eb45b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h209b80b13263fd120ee77a289;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h195498cd01bbb8c87ba7a344f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0343d11ef6de8803b82edd4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7e7e930cedf4f8158ec40907;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30467de5f37306d7faaaf51c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27be92b00e4388e4db2156289;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had3ad8de63c5dfc4e8a620e70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1876023f5dbdb7ef7b9b9e96f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14e7d33953135b6141f79ad7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56f44104450c17edff7e6fdf6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h484f20d600b466faf3a816441;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab7a9f765dd4cd110d9f9c9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf35119a492e37ceed788f9654;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e8d6bbbc92430baff6c47757;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33d5733be8941c9c0c622430c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68f3ff7146a1e2aab976d9581;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfc2fd397362aab2e9564a6ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6766b89b0c92a76aa07f7ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha09fb79dcf6586202fb96ee3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1818d21963d47db0ce7d1361b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9286121f6c0c612892ff2472f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67ad4035375be30007cf417a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4736b4ce0ea53ad8ec1f91df4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13e29fb5834800781bcfe7728;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haee9e3453988a09f9a5f7ff7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2520cc087f4622a249487e481;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89193d946db9ade6702b040b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58801bfe3bb6ce40a624d8a10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc40dc8a9a57d92434b9bcd868;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec5d5eca65d155ddb57702327;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2caa65ee284b97fa025c2b5b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a63ab6fdfdfda82f40aa218f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6beb6880291bb9e83347d2b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a56af2a55c375586571b6cb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c50511db0b84c5aa45b377a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fa9590d8633547256a80ff53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5aeaaaf7321d28f29701735dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5418f4bae526fce22568205ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h468e4887949e5f62317ac5b92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18ce35f7269f7b9a087d0b41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h876f9ae294a71571723a2762f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7abb6e7c5f4237804a180bc6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fb574f1fb6e9790025696546;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb53fbeb784691b5330302b20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41e179a7834904c4da546e950;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88b790aeeb0f81936ea5b0728;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78e851ed36e97aa4b5d60ca21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f02b441edc7779ff1d671784;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89c76e262ca19caad48136f70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ec983341b159857aa8f04618;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44c3559fb28cf4525a6f3a7ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9c9ab6e85050b47bc40a73c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7da626b5e661915b19c91c64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heea8289191cab16f83d3c8574;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17b4a2a991fbab5abd87ceab2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2882193480ac7227905f1ec37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h108442d2c2a4ca8406a3e44eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4f3343c5d0b875f413c1391a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd650d0f1043a010c7f372fb9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4908a4d16b1d6effeed0b7efa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c2fd8f417b9b32c0445ee19a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe109103e6a5892de096563ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9c2dbdf619c8983769124bb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27ba7b0fc6ed7decfee56c36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'head8f35e48a1472defd498893;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb6e2d1106a70128da6230125;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49da489edf0f09ac0fd2ef225;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h967a7a7555e590d071cd821ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc40d4a078faaafcb4e229145c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1786ff0f0cf9c71af70577889;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0c1417c828d4df67c618b465;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b8b1a025c8985fdaa95cf633;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda96b0f97724574f745423462;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79a1302cb8048d976773d9dfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5520af52eb4045af9dd296bad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heaeb4ff5dc4f65749d7c20b34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d6f0e48d6b56b50fb157201;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5deed849554565323fddd57bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81b2b25a7058d8029b6354a2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34fd9e83dd425773a2077c69f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc2fed0e442a881e142e641fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbab6837def2e9fb0fd04110d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f619800bd4ae7d7e25b22b44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e16cd8fbdb1d508073453f32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa6c9818bea36b70185900115;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26460c4a37e47b178109210b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd593ed212a3c5f9d8dc423f44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he942713b8ab48bdd0a8fb6386;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab6fb7751cc11198a4720c9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0e8f4e85fb1b66aa515e5b04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3ea38bc96dc63cc99c5e8c11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h937cf7f2bd1a092dcb16e78b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b71fc0fe43216663219d8969;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had5511e41f4aaaf68717b77f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5678d0d753d5994884ae715b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heed414a60ac6cda58ba2eee39;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1e4c9f279aa104b3201bcbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83544a05a66d35696566e8ca8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9913520eb65dfc3b343f42b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h211b360f15c8312e1afe5aa5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b2d5c3d7187243d7437d2f97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53cbc57e80188ef7146a3e6b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha09ee9c18a9f5e1b139edfe6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20e2f23ce85b7ae816905294d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6465964753724269d0bc288f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cfd59ad7a8e7bd1eea79afe3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30f31b2271403fe40e5319eac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc773192539f2639584d1fc18c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4c44d3ac1a8ae0d206ce2d82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heab7ab05a1bf80e2f688263de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2268d07b3e950cb45b0562d17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8af9f7f4cc16f3f85819fc92d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he07f3f0b43c962943f1cf711c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3aa19c71223527e6184c7ce6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h712d067a0872fef6e96167e71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9a532ce012540871871712aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ffe4f3155400345e669fd342;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17af70c32abb1f20ac38c35e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93d3e73afe530aa5d10c357b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafba28427b6d8e0c2f0381a5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30a638d8e9a61e771a5249532;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc487d28d4596a6398b791b944;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22f0a9e3fad50a4ab04a57cf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde48f5440429c7e5981b38daf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha74d35dcdff2bc320f3864d29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8084dfcd2041082003695e9d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98adca925dcca1a74c7ea7d57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d5ee9c411ba8a2fb8bb484b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h777a643983488ba0392d57e21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9388a7026c9988f1961e6bedc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb02328c3d5ee8972c2b038e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3de7e187f56a53bb8f2daba69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha47f5c172c953b9d88feb0544;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1921db9956a883369ec8aeefe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c5801f95809072d243ad8623;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44ba1a1562254a63a8e887b91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd122322530ff97487d5b3082;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35eb5936acbb7d4f38d088af9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ee51d49ed6b8870d33cec292;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57120b32c744c6541d03dab60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97b2f126ed8dad15464e6076c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd81646cd6fc61c610bab0132d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c5fdfe2b371f220b3069482a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he52426e345024af7715d1a8f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87e779f4827031ce15d5e2f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6595f7308037ec628a1842cc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7dd64297ef7c0b779dcfadcd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc798db9ff884ab237a34c9e38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h617edcf003d84240e991d5aa4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h239917e362b339cff4c2addb6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha557944730dfbcffa464209b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3ad6fa0a99ba0c5debd230f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7696193131c0256831457617;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5a8a5bc2e5e5bfded2a27552;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30f9d8d41000195637431e775;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha32e66fb61849f5a0e892b8b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae879de2f664064d6d385582e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47bb617fa2e2dd31e9afb5256;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e8b823f4ed661a79bd08bdf7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadf885a2f6111b13e973eb33d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbffcd2ec44f707be3d80e8ce9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6568c9f92ebab402d2632b3c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf982db4e92c7c18b675d2c7c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2db04068a1e100a79ee0cdaa6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3bf4cc3098b03919df4a9ecd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h311a52d52c602bb55e39adbc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h678f59d621c213b3f6d76e055;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2bdccaa489db609925ddec7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5954560bb55903d05254a27a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a20c11c0386b2c12fa1eedc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h822162ec7ecc187a078552f12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he94c9364aac5d98f63296d518;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf114a49f6c13cce84044863ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa05e4af4e6626d236455363f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f898d740426c780e08366645;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1307175f40aa22b5fa93fee31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h984431a5cead6b7c9f88b77dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf69d4abd3adc078e95f722767;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d2c7bb61b607f032273f2a60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7392c4ddf643d5a00bb4b048;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eb11f361bb8f59db3646736f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69c7973c2cd6eba792d09ab3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbc87d8889aba282903ed81b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae510f8076c194604cd68a27b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66a820039f2f60a45226dc9dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h698d98b4fd5749d61cfa24bff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h270f23fecfb5be2a6f72f5bc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef29fa2f338e011b945b61c77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38bcc86ef6274db2ca2777e05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd101ae40a5c5a8982bedc042c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b84e611be0453ffd59316403;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae76d6320bad3f10aede412fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dd2b0ff13801e22e16bed2ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h844c21367d71e5c6c707884ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2dbf257a5151c5f0284e4660;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2111843a9e1301425729f8f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h662c1ac6793494ce6aa3e8096;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78befec9233e5a4fa5f11d633;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64787510100edec85e435ea2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h496062f486d1f8506ef90104a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b6e58648d1f578559f9f3be5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9aa2ad808507fc07348ff9fc1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e016880f212bda4128218585;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h516a4ae791604c5d539910b1d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2966a0d8831e04c220690adcd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbae01b0321925e8ca6d1be3fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf76cb1ec202886222970f7ebb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfd16379efd75d5b8b3391283;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he100575659c99ee1c8dd0e303;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcf5fd90e2f337839cfb2a29d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6edce3a0df73503d515d0f456;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11746aec1d9523751450d2206;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd7ca2cfd253d0fce953b4fab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf98336d0cea554dc9876f8dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce535be7919293f36e84784fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h452f75b4cf2d4aa16cf59b438;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h601d97e19cb4c4909ee4961da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd1bd59e1993ba8b059df31cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67ac67187a71fd03458221b59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heec657a0839d3d83fd944db4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97ed9abfad5bddc9ec829d58e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c2bb2bdc45b63a55e9195b5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aecfb02675299ee9b1e770;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9dd410fe400b3ef23db5143;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf15eb8c20a8bbfca9c2678eda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72e2b6db49dad3da3981ce837;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc90cc119258d7bb22e9a5933a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc59d1897409b774b82e60c2af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d19a01486301faf106cb5701;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34fecd9395c16822e2f7f2c15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6890e3a9daf2a042d478c73d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h262690850e354e025f5d4edf1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha02985270f2838604f569c1d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf04d1bc8ca8f6a2b8e86739f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14498e7616eb2557c642d8a9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e632a2f25f9cfe9f2eda5742;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h333318d07243908857c8c75c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4bf15f6e86e15a2336b17b95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f2171df7ba50c6172086522e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a6460b03a60119d9d0f3d3fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc0cea480a06bf2aa55260c7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81ba824399df3db18044e810d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb19aa3a84e8ffd4880cab050;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1913e18efd69d4ae96020107e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a3608819f32c2ef43aa4d9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5974f5b7a099666248f3f367;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c1233db82a534747f751fa10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15b5e4532ceb7bf32de33f543;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2c24d5a8bc41877aff16d2ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8831f29b2950f02f37a91bfbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h147b24ad5b0e7bc84152ba7dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeeb8b407e25bb77b3b13cf7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d8236f74a2bf5e5fb53cbf4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75b2876107a756092c65cc25e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf814b183e62faf8488ea1b226;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42faf42e73afdd284a748743a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93cd57acddd2740fc69f334d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0027e53c5bbd2383f7623d0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12c991c2e7ee5e17e308445e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c8e218ddcdd86f8669f7131;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f512357c8fd52ce29d73f398;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5890679291ce53d74d85b9ba7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haad4878fac3a6db474dc7716a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h531ceb3e2afde8f5dc1bdfe6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h642c74b2236624127b926e381;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd82c472dfac82d58b309a3ad1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b36fbf4932bd26c4237a1b51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h331a1e5630465d968b85956dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c2bf9a6a05b2d657f74ee054;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e4a89b96c2479a4fb85ee708;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccbb157ce11aa10d0ff3a4b70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8903ab54eff84290ba3513af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h506475d38e2acf374ef4471b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52905bbbc2bebf0e99a1db3ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f0cf568021670d61696a8eec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e059f4aaa38f2e5497651252;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdabaf5b23d7094fc7e12f02c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ee9d8da4e3c8555295022d01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h284dbcbccf5c9b2da1fe70c52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3557658c49ab1db24ca5b3e52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62fc44d15ef52536d7053fb2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c55340c61bb7f18c99098b2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefd35dd32c01729b593ed4a2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90b4a74607b7a88f63538effc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1f7cc31b31f3be97c88f32b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf150e454f95888e06afb12151;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haae2a90f5fd994b719e7b78d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d5517f4cabb0d9275ea240a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8adb87d04957bf9aafa8ed4ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55ad43199e31cc16de5ed2958;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f54632aaf038542b2bb6b32b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h821fa2ec62aa7080b40891b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he45f5939ecd9989d32c3a4f5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5382e56788049064c3e0debd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hace6c9e47b945ace38ca89861;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h510e4f7ed7653b13b4291a98a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26e667ee7dc357ad1fcf99db5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff182d3db3ad981979ecd885a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e62bd1a2982838cab5061c77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1ee8b3dae849fa11294657a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84171c9fbffe4562c7c3fb918;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h611b6113f04fbe0c51fc993cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he49de916793806b798e8c3a05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45c88520768a338f784325318;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc44f3583ee9b60cc613ac9e57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b054eb4731baa938b81da570;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20c53da1e9c6015f0b190e576;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h850fbafb197b233eb4f4fa1b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd257cc5a01aee648061c3f8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55b3d52f76e698b60f9d4ea63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h788b52ba2f7286abfb6297d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbddb8b41167588ce1b63d8ee4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18d2d1df8bee553d0a06aba99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf10ba357871c1e33f7b164f31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h493f1bf45d07ed17d0456832c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc0e041b8dfc54f3326f1a052;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf16ab500e505725b5842149c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d978b6daabf65e13bfd88785;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h895f1c9d1c8ba80f5d84e04ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8187e9a935d62c0939aba65bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f8e84acfefcc10ca99d4f1cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2fef624e71541f543ce0f5e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3573b2975b2f50686ac378dd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc100a3062fbc33b925c5217d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65ff861683f0b5bbe4607b522;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13d3fa6f203b1f7a23bfb9f74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac269341ab85dac7af64c32b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c394eada735f515eb37dde5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8722db57eb7b894609f5f2af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf67c19306f2a64e3529673cc0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62b13b423c37e6420ba22b2c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ebb8ea4b5d90abe3b8081024;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h365ebfc50025893a27433b76f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8562b3a1290e3505a6d734f3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h321979e99a70e87b607299e21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h390e5f06f4c6b43be34732871;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a3baef903723ea56c15165fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbff6ec4c5837cfa29c782dc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8838d71b75a4543d4740d995;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12bc3bab4c0986b4126830bca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c67d618277525c209fea5969;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21245eee5a3d306c2bb5c1615;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bf11f76ba99f8091086e7b43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7eaaf7f7802f12a58c15f3c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a3303413ce8ab6364407f757;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h746a7ade6d50783c5832cda1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h145af72af86ea0be8f28effde;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42f986a51ade7d15f47bec462;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf51a58f3b9f9b85087f99c5b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1718e51a4cc3451e66788e5d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b8360dcc0afe32cc166d00e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he59aed380fef9268cfdeee430;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h404901b8f586f15abb1f03eec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h376ed363c9892f9b4fdce7472;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98a6b4ea5f5aab84868552bfb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h444c6d54e8ef8304ebe7ab8f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87f609a63d2a734bc81c48cbb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9d1deccbdfee690218af7574;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ce2ccbaac5efa6e2f67beaa6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73795a1815e804b8463fbb654;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hedc381032b1c5daa178b54eb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc814b7b2c473de578c50ef753;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e5e703a8ad16cd6ecb1afbc3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc19563657003da6fa4e8f421;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24bbb069550d30a697436e07d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ab9da7af31fd00935b74fce3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5843f5ce76d75c9be2c51afeb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d43f8a05ec90d2237597b1a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h823e785b05e0a1f684c3ac9f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a15bb5c197c0f4fc0ac81148;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57932448dfd5ac103b3b7136c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ffbbd9f58af12bf66d35878;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he31eac79f8debf12f78c05cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eec4cd4e045a86226fcd5fab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71d51fe4d42f23650bd64ac26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9e9e7c67e8b35730506a8167;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a5e5676f3c86e45821874e54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae4fc308a67fa0b3c8bf0ba7d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6dcd4b2be525ff8130cbcbd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcb13edf3aa010cd901b3277c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bf0dd210dbee1c706053e3e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6321041efdb8edc9b977c4d92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13503509bd10ad0d90bd7b5b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haabbfd19a9b0685521ef51fcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc7f76040192aaba7104ee938;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5593ec7e75abddb86e78992a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h943daa263b2337c3f737465fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ea702d4d94e406eba2c208d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57ab1df8f31fe51b729f2e548;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25e747f2a9f4486c8e1f58376;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb9f4baad8c530ce039af726d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2e69737efff1c025d440cc48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c79d663bcd36b705e89f76ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9326db410650041f2eff1e1ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5568a6a7fe2e6366a910296f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ad0d590fa1e3a0cf6dabbd82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h871335d1fb51cb45f099ce93b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3edf6c82db4771af4d0727ad6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h192e532bf5a8719ccda62ec44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99b516091060cb2743e8bd6ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e31c77c26b94f254b84879bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0347db57913ae64b81d1b617;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8908fecc0ce0161a0b8e7cbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73acb0bb41e7014d6b8b391fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h230333edc8a3acd0cc369e6e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e88a6a8eb50e9c43cb179411;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf44a8aa04ab794e745d9c695d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cdce9232848588e3a8978d2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd29c105a00e94e0bd99febbca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87f86845f8a54760950cb71a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0e42e043d0637724f4a866a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c20a1a960c73b57ed85257de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33df6268a118dcb0513dc90fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28e4ea57b03958506ba5382ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h719c5a7beef0da95aba26b5f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h554dca847269df1837a1b3a1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h682f6a4e7b9f1b3d6da78064f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38988700b347c28783cf9fbed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b06eac5ec8401126e37a3c86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655efc40708fdd5d187c18c5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b064568873a71692aa7f21c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h720438428915dc11cf4fdc3af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dcfcd14b67ed4d8fe43be2d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14d5661e644d5b6b0db79ea35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb55e456335c5f229d6cfc41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55840482b380d733dfda23a72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h783dc7724b216681f1f9a9fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h917cd3a5b9021cb336b787944;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf55c5d0eb3deb7bfd98364f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc83d92a9df77a0ad679d88f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f1076d12d2449aee4a2a3be6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6d491db0a6745d5920db776d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47a7f9e0c62fa855eec994b9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dd328f2e561da2ee1e26a83e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h225f00e0da3c888f33fdd06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9a31d2d5493c813c1bff0e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3741e664163be5bd2306f8494;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b037bd2437de932263ebd60b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde05e4c92964c91caac6627c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8bf9ca398e7057fabbebed97c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aa8e60995b72751819f575de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb425e4a087e50cbf086c525e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90bba28e05fd7514ab4f62d45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9589a92b1f77e8a5c6a8f035a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa8b1d7f6ef96a8f844c82345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9abe096f749184a8f0ff56a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda352d742ac01a275ea48d9c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31411208c8ac925789b8f62dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84e8a09d75dab5bd543e236f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c1f5ede031dadca6cdfd7d21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fca30a92ef90130319f91a7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha522a3453070655317be2e962;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb87b701a278c1200927e461f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf4aa050ceca8203d9bc020db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf63a84e487015dfad231a41cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb449310d806c617399524534;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f5c11106705a0b9e9988d574;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha08295bf2fe940d7f6d47cb9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e450051d2220bd57d209a1dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7367df9a59424f94424982f51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73d1d9481749071313e8a7585;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h129f649e547e8fc37761abb6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f1b00969abe15c8e8de23a7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcccb9c466706bd5f5dfa8976;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c4a81191ae7566b36886495d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33a45f0b143608dfb7fc4f936;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdef7d5539ca664d13c5c093de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81ced0dba7a5f9ef8d5bcc016;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf3bfbec5a75d19f7000beec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h880e6c3aa256fa7a98d4554c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfc455df49ce5b4b3c04c3be7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9066b2f87cd7a178128fecfb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40579e0de012ef434e40b9852;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9778cd47d44589b9e18ca4f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd88824c925049c49a44052043;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655c82a5a8ebbeb88736f016;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90b061b29a1d5f80b1356b5d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9478dbde91f22bed6588137ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9849eee743435d1947c4b4a88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ec9ce98a21b9848c46bc3b84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h716ee5827adf33d27c10f9d03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbac667d5c19c2ba3fd1e0120;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf44c4bbd45e94b8b20dd60b9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca8147cb5155951e3b8ede35e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha03909df7833d029d1c4a20f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc69ce0b5b422b750be47eba54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73fa436ae0a177ff4ec9bba2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha86517fe72f0a45f1def9e0a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc94cc9640cf37003b9ec957d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d25e493e6845102f5cbfb07e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e555a93944e13be0c0dd0d66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef20392ef735e98872164d64a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81ead6117b496456acc7189ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b6e270d5d55f992d34451c72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec70f413325f1a7175063a5fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbf6d3fa9f1f88e86d76f44c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55d23fab50ce6ae762a543673;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5170e83c63dd2db753837f540;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd55eb6429e4021c8e2079ad5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c06904e4343cb12825585e52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcaa7065139ec823e4e93c445e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e7a041dd246c01b6474dfe7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac20ad5d33e676448017a9c09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5a5808448653ebf6cd767143;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36d3229a982cb8b7359021027;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbfc60462ee509c3234ab8858;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h826072295bbabe5450f9cf42c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd659d79353b65a662cf04acc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19c6c2795073d14096acb500b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6db2014c78eade30fd9a9c9ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h359469573aecd04f6acb290ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8df5acde2fb1ca78d5f01a319;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h957bd6722e5fed3bbf6cb36a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h168fc5de71041b64a5f8e0976;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23f7f406ebaca5edef1919e5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4f8faa85d6a8bd4df4cc5556;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7b15f42b55f537f047387d15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2b6144529093834484d2b6ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h120fa20d6b28523f1ebd7a64b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbee92ead70010b24f879347aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h521b5dcaf6245ed1786164eee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf42164477a3ff7ef3c8fd9412;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5be739a350407e1aa13ab57d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7504fef2a3b74eb95bd592501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ae78de683022819c09f927ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8356de0e93eb967998706ac10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9bc4909dac4411038fa07d94;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffcaad41e4805c5ca297c96e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57aa8faa0952171e1ddde3858;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61e273296f3c964dccbb9542f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1303e88bcadf740fa1455ce6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4b91d597024282a214681dfb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h788535752014712c313e2c1c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a3b84888dd2c8fc3ef2a698c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34968ca4c042b4d79620312e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb81d986330964638fba150854;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h949c740b18acdab3248cc8eff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42985689196ebf7ff8147f59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde30c3ea49d3335d3a5819ed5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae0abf647e8c75fe87e7998a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7adbd9cd8129d4de04c4688b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43fd5e7ecb78e49624b68ffe3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61bb4deac766609f6d314a37f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd076b374f7e25b365f9e024bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3462cf72948b69d138575585b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2241b1de165f699bbacfe5771;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc45697c223bf207e91d76e7cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4d15cb1bbc785698673ffad6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f7381316f94241e15e848be1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha666710e0b1308e1e254ca485;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d75368cef5036862123b4ce7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h864028f15c1018c9542c1e358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3064453c66e98973129bc5d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7d7941fd6f0880fa15a2f1be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97267f7e31d9906498f22f938;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf215923aa3d1f9375ca98b6df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a42bae0d7f3aceb55acf9107;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6852797cf65e7d46c74357cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ef017d6a37416c4c6c0383f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82a294ac55bdaeee8cedf452f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4a72adc39dc2c845990926ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4536fed59d13dffa923af25bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb21a7ff35773ea00059cf5971;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h956b5978cd82d23f95e8d3c22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha877ce1ea10826e3068e168d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46c3c54daafe78316610027d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h548d206522f35b7d29cbf7d8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf722f1a43571d9086584c6758;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37557a4668589d8c4bda4d369;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff8040b8575985e9e5cec4a5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24a5ba3eee9addc5c3acb4c3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72e898f40430d1be1aa890841;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h171185e10a14e47d6db225723;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1fd7beea18bac4840598e08b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h792907f552d1d6ddbaa64d169;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5325e846b0471861bea525538;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h467e30d5b6a407a5a6cb373b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd6e9ed9d38c0a04663795195;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5a37093dfbf5fd0cf89145c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a03f2cb5ba28e43759e1397d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45ccadec187437a3657644087;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h839b020e78d8f37da570d5df7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5f8b1f60934cbfe88a574f1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd570ba7b92d1f05f1d8402367;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha13094e390576b38cb0343499;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24e92f2414197a6e0a48311aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf9c0c484ec733ceb3d38e136;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54e429b800097fc5478e1965d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha22c85e36e1fd8c84845a4747;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2998ceebcebc4b0cf2700a58f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0f0dd065b9bbcf2269e461e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94605a75ee4a078be9875105f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7a4e9a65e5877a7021c2a12e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ca9b4ab28291ce32cf8549e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23070a30958efbcf13d336a28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0c181f6e6838f33491444355;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf07ad6d015b752422de1e57b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd37bdc3aa74b6b76ab5ab36d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41154db83dba738246dd30d04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf49ca91511e7d963f9cd9a057;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e57d76e12b446cd1300f38a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8387d8e578a6a7ff46ebe467;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31b6d84c42a39bc18c5261b87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6785545d666e248b19c41aff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h168f3a1f4cc33545458ba94fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf01df9c4c1302ed05c547be06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19c6eed1a72dda8fd92cd4fe8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h245ca4e5ea506e657b5de2677;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda19152fbce4473aa34d61ba1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfb4be54550dd1f2852eea2b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46b43f5dce9978db1ab2eeab3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he60a35707068fb44bbcbc6dd7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habd2e0f3d9ceec302b2042eb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62477a09dcf8373140c8ead24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h450e30ef8b645f761cb97d5c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2071a2acb343e56324a876799;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6ce280a96e60340b60ecc6d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e50329eaf9353a71904fe1d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf535dc6ec8480c7d8be717de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22a6e1c3ea4ace602ce4ccb8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1aa2b6b9bc08ccdb650dfe732;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe4f2a965e57a594da1bc06b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1560ce1b9371ee3d427a76d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c5d4634f9875cd4caee36794;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h944d7607b8572cbb7ba8212b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc82b2decb05c6bfe5fa83b8d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h348a1062c0d1df9232895da0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha683d0767022165d3107f127a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h819894b0d15d5940841d2731a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50a7dd9b1e3adbfc0c8824641;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h724a89a913c20f3e02e1ccbd7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37e1e04cbdeeb2690eec5c8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa10376317416f3698f5596fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c08fc07fe966eb92b7442a53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c7d869ae1d833c8952e0b56b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h754e94818d53f8226e47d177;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he742ca979908ad141437f535e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa615bc89782d79756913e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da1414188c4a92a6c6cc2308;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5b1ea5be4bd733e67f273f89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h799e6d0630ce7f88fc2ef079c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66f3819c24f527cc718648b1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36028ec57c415d9c9d2bf4cf0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70fac820fd1f4b245b4d07598;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3270e92b135d7e895bf18a14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d778df74a1f59ac5d928df3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cbaa62770f9944ed4334d76c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61bad81c3f6b8fac28bf501b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ef739f0bcac51a2aad088952;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf32568548dd3c068766b6d53c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6542829393284da691b767aa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3372dd9bac6acd6084d88d22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cc9436352a02b6af55116aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae44172345999fbd80c9326b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84654b77022b731d968db0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaffc774a494d0f34f174187;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a60e71e17151575f91b111b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73cb8df85ed221a2d531eee7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb627d4f55f48f5381e0ac3166;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e59fadd88c4039ec17529617;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2695d2ea7f75725854b66eb48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfca342760a402fa4add6b89c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe9ce698d2435b3ca1c11444e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c1157e41d135d60c97852f85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb719dce8c502f6a61282f7af1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha853ae6ef0ddfe54eae023e84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa8ab29efe7683ad37ba1e7c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd02decf7c13af72a25ed0abd3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f3acb06499a3bc3182e809c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeb85a45e89837e46fb608eb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94951d1ef64dc1f9111fd2bee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he72ed6f5e16b1328c30e009a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha117b87582c19b8ce3c2e5158;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h773da4493b867e639440fb8b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haee11d828eb5d76f5c1143739;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bf478fad63c1a34c9a21e19b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h267cd46ad7a51d40afa4b416;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h338c098d3aef160e126f771d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5cc6aed05525053d6ac83870;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93835c94d25c36872d4f18ab2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b27a7fd80254c5742b4be1c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h428a817da8e9656ae8e88a2e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80dd7e80ce3316fa244e291b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h749abeda5984530c5c1308558;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h867644fe3b908570e8fccf08f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h610e31e7fc2b29c2a6e224183;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8403ea7e86a6a2041765513e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97f6cb5624caffbac91c2777c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb99b7406e1fd0b2d30e780ecd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a63a7418190fe27cbd6a675d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c05e541859485f7f53616a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa6eca6075f8ab0002c14797d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb5ef416ed1ab0029a776d727;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heac1fbafb79b9b57d13f94a78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e6eac5eb254347c1edc7726d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h727972320ea1ef499a0f1684a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39e370213061835714c2950fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha71e908142049b9ef970f70bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c3015eeb855a2da3ba923e97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcaa8206032a825d906b1f391;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0b619c9c6ef788ec1ae74be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha753efcc923ce495b63daecbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65f4e5de087a4d355f8a158f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h709855b9457b45e2f7b6ccdc1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e52b0b1acc116bb43b31e1d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96fa2c6686b92558a48003b72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd952dd79369757d9166202ff2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he16d9a6db29e8e9c62e702b2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h385c4b2968d16185a62c3269e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h909743d6629bfcbebd5f8f626;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h885fe124eaf99771802887b1c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2a133be85ef0dc7b2abc64a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1aa45f6ab55ef7f219293468;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefb801ae10f19b6d85608934c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heba91fbc61291967aa7c3907b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h890b2e592eddd2a2201f71c87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08b8094037eba0f9a27d5831;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ef5fd3c0ca1f591c5e1d29c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e028952141bcd2c019af3dd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he00a16749764f15fc84a9a157;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ea72ce1ab5f3e1a0d1515d93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc95dfab32fd9e9ab90894b08b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5641f54a62cedb6629b6db682;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65267acd223306edf2c8879f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23355f0225465a75745948912;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56da03105621a24cc62d6ec2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a3925bc0ac1678556cf25374;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ac1000977410c3c6ce92f04b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88f6ef2ceec7983ebdbdd83bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h374f0e19b8f8514ef159a90f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47c2c0c70ff80691ddb70587b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c1a2ffe38e4054add5eae8ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8575b3b2fb303fbf910a2c784;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a59021acf8e6a77a4a924b08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he79feb47443873dc45b88d579;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65d42afc31c58379132c39c99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb7f3ec19a0156a229dddf899;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21375fd122c3aa378300ca45a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb2984fde4c77c5dee5d2decd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57918ac2ea9d416caa69aefc5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h304303e5d574c1fe8bb5f637;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22016d1ddf76364f20c7fe27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h531b82346c31f6d88db5fe951;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf539f548ae936c08d2fe5f0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd296cc5acca0e540c650521b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fad250d0a3db5bcc44fc96ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h359ecd555bc3f6085256bd02a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdb84c8e46f9ca6ba539c03d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd7d69cc2d1b98132a4dc8e0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbd373709792317ed464432ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc2520d7551fec8565721719b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2df6eb4eade3f278719fe09d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d21628aeb8067e1c215c61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37a66c8057e1a333e56f5813;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bdb411065d8a9243fa0145eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90b379010181dd742c6b842da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb676a6f372ceb8acafa16d53a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f946bfd8452d5372489abb27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b2a42424d3976320038adca5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f404bb09c8434c65a6cbfcb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heacc2960ebd41e4854f7fb474;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74df480cb48a912be5a8167c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he34f0ea806017eb4aa78f7e2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdccede75bb13eaeacd73b7801;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h952c8b01c74a7fddb5c3e060c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb3ec94bd955802682f90da5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca748a854b0298af3c1c3cccb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7dd6afc075fc8de74202547c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5a8ea6c134e596f6704e410;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9be5ff122aec3f27f67d6abc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60311ae11e52e3cbd506880d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6a7ffcfb17a059e7b920c2ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f92347cab4fd75a163eaa74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6d0d89555ad732216e8c7af7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb31e97f37987298164f38415;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7656c13c70d6e8a988a74663;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8935835e470ea9e10d01e0970;
        #1
        $finish();
    end
endmodule
