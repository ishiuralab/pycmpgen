module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    compressor2_1_32_16 compressor2_1_32_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_32_16(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    rowadder2_1_21 rowadder2_1inst(
        .src0({comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [14:0] stage1_0;
   wire [9:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [14:0] stage1_4;
   wire [16:0] stage1_5;
   wire [18:0] stage1_6;
   wire [11:0] stage1_7;
   wire [13:0] stage1_8;
   wire [14:0] stage1_9;
   wire [12:0] stage1_10;
   wire [10:0] stage1_11;
   wire [15:0] stage1_12;
   wire [17:0] stage1_13;
   wire [16:0] stage1_14;
   wire [10:0] stage1_15;
   wire [8:0] stage1_16;
   wire [4:0] stage1_17;
   wire [4:0] stage2_0;
   wire [11:0] stage2_1;
   wire [1:0] stage2_2;
   wire [9:0] stage2_3;
   wire [6:0] stage2_4;
   wire [8:0] stage2_5;
   wire [5:0] stage2_6;
   wire [6:0] stage2_7;
   wire [6:0] stage2_8;
   wire [7:0] stage2_9;
   wire [5:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [15:0] stage2_14;
   wire [3:0] stage2_15;
   wire [11:0] stage2_16;
   wire [6:0] stage2_17;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [4:0] stage3_5;
   wire [1:0] stage3_6;
   wire [4:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [1:0] stage3_10;
   wire [2:0] stage3_11;
   wire [4:0] stage3_12;
   wire [1:0] stage3_13;
   wire [6:0] stage3_14;
   wire [4:0] stage3_15;
   wire [2:0] stage3_16;
   wire [7:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[4],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_3[25]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[5],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[6],stage1_4[10],stage1_3[10]}
   );
   gpc606_5 gpc11 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[7],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[8],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[9],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[10]}
   );
   gpc606_5 gpc15 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[11]}
   );
   gpc606_5 gpc16 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[12]}
   );
   gpc615_5 gpc17 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28]},
      {stage0_6[18]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[13]}
   );
   gpc615_5 gpc18 (
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_7[24]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[7],stage1_7[8],stage1_6[10]}
   );
   gpc615_5 gpc19 (
      {stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage0_8[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[8],stage1_7[9]}
   );
   gpc1406_5 gpc20 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[9]}
   );
   gpc606_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[10]}
   );
   gpc606_5 gpc22 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[11]}
   );
   gpc606_5 gpc23 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[3],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[12]}
   );
   gpc606_5 gpc24 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[4],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc615_5 gpc25 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16]},
      {stage0_10[22]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[5],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc615_5 gpc26 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_10[23]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[6],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc27 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_10[24]},
      {stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage1_13[3],stage1_12[7],stage1_11[8],stage1_10[9],stage1_9[13]}
   );
   gpc615_5 gpc28 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_10[25]},
      {stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30]},
      {stage1_13[4],stage1_12[8],stage1_11[9],stage1_10[10],stage1_9[14]}
   );
   gpc615_5 gpc29 (
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_11[31]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[9],stage1_11[10],stage1_10[11]}
   );
   gpc606_5 gpc30 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[1],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc31 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[2],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[3],stage1_13[8],stage1_12[12]}
   );
   gpc606_5 gpc33 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[4],stage1_13[9],stage1_12[13]}
   );
   gpc606_5 gpc34 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[4],stage1_14[5],stage1_13[10]}
   );
   gpc606_5 gpc35 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[5],stage1_14[6],stage1_13[11]}
   );
   gpc606_5 gpc36 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[6],stage1_14[7],stage1_13[12]}
   );
   gpc606_5 gpc37 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[7],stage1_14[8],stage1_13[13]}
   );
   gpc615_5 gpc38 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_14[24]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[8],stage1_15[8],stage1_14[9],stage1_13[14]}
   );
   gpc1_1 gpc39 (
      {stage0_0[21]},
      {stage1_0[4]}
   );
   gpc1_1 gpc40 (
      {stage0_0[22]},
      {stage1_0[5]}
   );
   gpc1_1 gpc41 (
      {stage0_0[23]},
      {stage1_0[6]}
   );
   gpc1_1 gpc42 (
      {stage0_0[24]},
      {stage1_0[7]}
   );
   gpc1_1 gpc43 (
      {stage0_0[25]},
      {stage1_0[8]}
   );
   gpc1_1 gpc44 (
      {stage0_0[26]},
      {stage1_0[9]}
   );
   gpc1_1 gpc45 (
      {stage0_0[27]},
      {stage1_0[10]}
   );
   gpc1_1 gpc46 (
      {stage0_0[28]},
      {stage1_0[11]}
   );
   gpc1_1 gpc47 (
      {stage0_0[29]},
      {stage1_0[12]}
   );
   gpc1_1 gpc48 (
      {stage0_0[30]},
      {stage1_0[13]}
   );
   gpc1_1 gpc49 (
      {stage0_0[31]},
      {stage1_0[14]}
   );
   gpc1_1 gpc50 (
      {stage0_1[30]},
      {stage1_1[8]}
   );
   gpc1_1 gpc51 (
      {stage0_1[31]},
      {stage1_1[9]}
   );
   gpc1_1 gpc52 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc53 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc54 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc55 (
      {stage0_4[31]},
      {stage1_4[14]}
   );
   gpc1_1 gpc56 (
      {stage0_5[29]},
      {stage1_5[14]}
   );
   gpc1_1 gpc57 (
      {stage0_5[30]},
      {stage1_5[15]}
   );
   gpc1_1 gpc58 (
      {stage0_5[31]},
      {stage1_5[16]}
   );
   gpc1_1 gpc59 (
      {stage0_6[24]},
      {stage1_6[11]}
   );
   gpc1_1 gpc60 (
      {stage0_6[25]},
      {stage1_6[12]}
   );
   gpc1_1 gpc61 (
      {stage0_6[26]},
      {stage1_6[13]}
   );
   gpc1_1 gpc62 (
      {stage0_6[27]},
      {stage1_6[14]}
   );
   gpc1_1 gpc63 (
      {stage0_6[28]},
      {stage1_6[15]}
   );
   gpc1_1 gpc64 (
      {stage0_6[29]},
      {stage1_6[16]}
   );
   gpc1_1 gpc65 (
      {stage0_6[30]},
      {stage1_6[17]}
   );
   gpc1_1 gpc66 (
      {stage0_6[31]},
      {stage1_6[18]}
   );
   gpc1_1 gpc67 (
      {stage0_7[30]},
      {stage1_7[10]}
   );
   gpc1_1 gpc68 (
      {stage0_7[31]},
      {stage1_7[11]}
   );
   gpc1_1 gpc69 (
      {stage0_8[31]},
      {stage1_8[13]}
   );
   gpc1_1 gpc70 (
      {stage0_10[31]},
      {stage1_10[12]}
   );
   gpc1_1 gpc71 (
      {stage0_12[30]},
      {stage1_12[14]}
   );
   gpc1_1 gpc72 (
      {stage0_12[31]},
      {stage1_12[15]}
   );
   gpc1_1 gpc73 (
      {stage0_13[29]},
      {stage1_13[15]}
   );
   gpc1_1 gpc74 (
      {stage0_13[30]},
      {stage1_13[16]}
   );
   gpc1_1 gpc75 (
      {stage0_13[31]},
      {stage1_13[17]}
   );
   gpc1_1 gpc76 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc77 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc78 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc79 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc80 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc81 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc82 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc83 (
      {stage0_15[30]},
      {stage1_15[9]}
   );
   gpc1_1 gpc84 (
      {stage0_15[31]},
      {stage1_15[10]}
   );
   gpc606_5 gpc85 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc86 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc87 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc606_5 gpc88 (
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc89 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc90 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[3],stage2_6[3],stage2_5[3]}
   );
   gpc606_5 gpc91 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[3],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc92 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[6]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[1],stage2_9[2],stage2_8[4],stage2_7[5]}
   );
   gpc606_5 gpc93 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[2],stage2_9[3],stage2_8[5]}
   );
   gpc606_5 gpc94 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[2],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc95 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[3],stage2_10[4]}
   );
   gpc615_5 gpc96 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[4]}
   );
   gpc606_5 gpc97 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4]}
   );
   gpc606_5 gpc98 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[4]}
   );
   gpc606_5 gpc99 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], 1'b0},
      {stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[5]}
   );
   gpc1_1 gpc100 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc104 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc105 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc106 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc107 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc108 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc109 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc110 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc111 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc112 (
      {stage1_1[9]},
      {stage2_1[11]}
   );
   gpc1_1 gpc113 (
      {stage1_3[5]},
      {stage2_3[3]}
   );
   gpc1_1 gpc114 (
      {stage1_3[6]},
      {stage2_3[4]}
   );
   gpc1_1 gpc115 (
      {stage1_3[7]},
      {stage2_3[5]}
   );
   gpc1_1 gpc116 (
      {stage1_3[8]},
      {stage2_3[6]}
   );
   gpc1_1 gpc117 (
      {stage1_3[9]},
      {stage2_3[7]}
   );
   gpc1_1 gpc118 (
      {stage1_3[10]},
      {stage2_3[8]}
   );
   gpc1_1 gpc119 (
      {stage1_3[11]},
      {stage2_3[9]}
   );
   gpc1_1 gpc120 (
      {stage1_4[13]},
      {stage2_4[5]}
   );
   gpc1_1 gpc121 (
      {stage1_4[14]},
      {stage2_4[6]}
   );
   gpc1_1 gpc122 (
      {stage1_5[12]},
      {stage2_5[4]}
   );
   gpc1_1 gpc123 (
      {stage1_5[13]},
      {stage2_5[5]}
   );
   gpc1_1 gpc124 (
      {stage1_5[14]},
      {stage2_5[6]}
   );
   gpc1_1 gpc125 (
      {stage1_5[15]},
      {stage2_5[7]}
   );
   gpc1_1 gpc126 (
      {stage1_5[16]},
      {stage2_5[8]}
   );
   gpc1_1 gpc127 (
      {stage1_6[18]},
      {stage2_6[5]}
   );
   gpc1_1 gpc128 (
      {stage1_7[11]},
      {stage2_7[6]}
   );
   gpc1_1 gpc129 (
      {stage1_8[13]},
      {stage2_8[6]}
   );
   gpc1_1 gpc130 (
      {stage1_9[12]},
      {stage2_9[5]}
   );
   gpc1_1 gpc131 (
      {stage1_9[13]},
      {stage2_9[6]}
   );
   gpc1_1 gpc132 (
      {stage1_9[14]},
      {stage2_9[7]}
   );
   gpc1_1 gpc133 (
      {stage1_10[12]},
      {stage2_10[5]}
   );
   gpc1_1 gpc134 (
      {stage1_12[13]},
      {stage2_12[5]}
   );
   gpc1_1 gpc135 (
      {stage1_12[14]},
      {stage2_12[6]}
   );
   gpc1_1 gpc136 (
      {stage1_12[15]},
      {stage2_12[7]}
   );
   gpc1_1 gpc137 (
      {stage1_14[6]},
      {stage2_14[5]}
   );
   gpc1_1 gpc138 (
      {stage1_14[7]},
      {stage2_14[6]}
   );
   gpc1_1 gpc139 (
      {stage1_14[8]},
      {stage2_14[7]}
   );
   gpc1_1 gpc140 (
      {stage1_14[9]},
      {stage2_14[8]}
   );
   gpc1_1 gpc141 (
      {stage1_14[10]},
      {stage2_14[9]}
   );
   gpc1_1 gpc142 (
      {stage1_14[11]},
      {stage2_14[10]}
   );
   gpc1_1 gpc143 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc144 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc145 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc146 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc147 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc148 (
      {stage1_16[0]},
      {stage2_16[3]}
   );
   gpc1_1 gpc149 (
      {stage1_16[1]},
      {stage2_16[4]}
   );
   gpc1_1 gpc150 (
      {stage1_16[2]},
      {stage2_16[5]}
   );
   gpc1_1 gpc151 (
      {stage1_16[3]},
      {stage2_16[6]}
   );
   gpc1_1 gpc152 (
      {stage1_16[4]},
      {stage2_16[7]}
   );
   gpc1_1 gpc153 (
      {stage1_16[5]},
      {stage2_16[8]}
   );
   gpc1_1 gpc154 (
      {stage1_16[6]},
      {stage2_16[9]}
   );
   gpc1_1 gpc155 (
      {stage1_16[7]},
      {stage2_16[10]}
   );
   gpc1_1 gpc156 (
      {stage1_16[8]},
      {stage2_16[11]}
   );
   gpc1_1 gpc157 (
      {stage1_17[0]},
      {stage2_17[2]}
   );
   gpc1_1 gpc158 (
      {stage1_17[1]},
      {stage2_17[3]}
   );
   gpc1_1 gpc159 (
      {stage1_17[2]},
      {stage2_17[4]}
   );
   gpc1_1 gpc160 (
      {stage1_17[3]},
      {stage2_17[5]}
   );
   gpc1_1 gpc161 (
      {stage1_17[4]},
      {stage2_17[6]}
   );
   gpc1163_5 gpc162 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc163 (
      {stage2_0[3], stage2_0[4], 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc164 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2]}
   );
   gpc606_5 gpc165 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc615_5 gpc166 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[2]}
   );
   gpc615_5 gpc167 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc168 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], 1'b0},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[2]}
   );
   gpc606_5 gpc169 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[2]}
   );
   gpc606_5 gpc170 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[2],stage3_14[2]}
   );
   gpc1163_5 gpc171 (
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage2_17[0]},
      {1'b0},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[3]}
   );
   gpc1_1 gpc172 (
      {stage2_3[7]},
      {stage3_3[3]}
   );
   gpc1_1 gpc173 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc174 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc175 (
      {stage2_5[6]},
      {stage3_5[2]}
   );
   gpc1_1 gpc176 (
      {stage2_5[7]},
      {stage3_5[3]}
   );
   gpc1_1 gpc177 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc178 (
      {stage2_7[5]},
      {stage3_7[3]}
   );
   gpc1_1 gpc179 (
      {stage2_7[6]},
      {stage3_7[4]}
   );
   gpc1_1 gpc180 (
      {stage2_8[6]},
      {stage3_8[3]}
   );
   gpc1_1 gpc181 (
      {stage2_9[7]},
      {stage3_9[2]}
   );
   gpc1_1 gpc182 (
      {stage2_12[6]},
      {stage3_12[3]}
   );
   gpc1_1 gpc183 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc184 (
      {stage2_14[12]},
      {stage3_14[3]}
   );
   gpc1_1 gpc185 (
      {stage2_14[13]},
      {stage3_14[4]}
   );
   gpc1_1 gpc186 (
      {stage2_14[14]},
      {stage3_14[5]}
   );
   gpc1_1 gpc187 (
      {stage2_14[15]},
      {stage3_14[6]}
   );
   gpc1_1 gpc188 (
      {stage2_15[3]},
      {stage3_15[4]}
   );
   gpc1_1 gpc189 (
      {stage2_17[1]},
      {stage3_17[2]}
   );
   gpc1_1 gpc190 (
      {stage2_17[2]},
      {stage3_17[3]}
   );
   gpc1_1 gpc191 (
      {stage2_17[3]},
      {stage3_17[4]}
   );
   gpc1_1 gpc192 (
      {stage2_17[4]},
      {stage3_17[5]}
   );
   gpc1_1 gpc193 (
      {stage2_17[5]},
      {stage3_17[6]}
   );
   gpc1_1 gpc194 (
      {stage2_17[6]},
      {stage3_17[7]}
   );
   gpc2135_5 gpc195 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc606_5 gpc196 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], 1'b0, 1'b0},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], 1'b0},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc2135_5 gpc197 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], 1'b0},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc615_5 gpc198 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc2135_5 gpc199 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc117_4 gpc200 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc201 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc202 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc203 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc204 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc205 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc206 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc207 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc208 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc209 (
      {stage3_10[1]},
      {stage4_10[1]}
   );
   gpc1_1 gpc210 (
      {stage3_11[2]},
      {stage4_11[1]}
   );
   gpc1_1 gpc211 (
      {stage3_13[1]},
      {stage4_13[1]}
   );
   gpc1_1 gpc212 (
      {stage3_14[6]},
      {stage4_14[1]}
   );
endmodule
module rowadder2_1_21(input [20:0] src0, input [20:0] src1, output [21:0] dst0);
    wire [20:0] gene;
    wire [20:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[20:20]}),
        .S({3'h0, prop[20:20]})
    );
    assign dst0 = {carryout[20], out[20:0]};
endmodule


module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor2_1_32_16 compressor2_1_32_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdea912ea642788207f350ec3bd02d96272e50340abb5d6794b714693653becd68dbc56a0c1f35818be56fb05d97a218844060100f19a71415870e31ddc2b565a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7f44f3bd43ace53c14124c5d105a343c01df3728b796b72e913ced0973008294239085b1e63a5fbe01e433d5dc53089270d2dd7155e1f2d1daa22fdb5f9867eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7e4b0472e3bb0a8c829a592d5c1caff8e475a3aefef5ce27a460b3f7a0f8babd35049bca5b82eb7951e8b1d04050a5eb09408171aa16d273f48688ac8475c64b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haa90d1d44d6fe4fac7a008b2b048f330c95818040f6d0bebb9973dbcee90bdb09f10a18e5fe2ff3d1ce51b62fa7d3afab55b08d7666dcc2be98b8deaafe6c55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h41d5c19ae8719a00db78952c74ce4e97b53b00324ae16cd80950dafcf5d2f475fc8814135f640a47899060e67599a291bd43080bc1c42910e37e930da85824b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8bb8973f31e90c863fa9ab158fe83ee555f8951beb4901a94a89f0cb7233091a2a5dca3732b703522f7549e96c06dafe234e8a851d002199d6120a038d9ddd65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7f0b1ca2474df6ce6fa7030fd9b6a406d0009a4f51c53463d8bb07074b24d791dddf3e2f661ec50ed16dd971d00127daa5034e3564b25fc8f621b0cbe906a2aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9136c3a32a440b4ee0cda127fc9cb541fd7e39d8d883f885fdfbc4cf518716d4c5336c704f8818c3f64f8d6095ae41b789f715c2124215d2a1d7e7dbb4ea881f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2f854d32ca31cd08bc52326d01c61983d61d903f12b8f51677ec71fbac25626e3199a804e7c1826418f83caf96bb2534971c738926cea0041776a6327ebb1a82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd7c8ea1b20c9ebe54e104db97e7c14499c7e897480ef4e674eb553e1eb8a41d101f61e7dee7ab3353ff0bb5496e91cf8fbdf8c83a2f5c1863de4e8afd54d315b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7bb7015ed48d61e2532aeaa6752c943a99ad8c73e3ac9e365bd1ee5e1221de6a53be01e2a9a911cef52f540ccafee56bfc700cee4bbb5d04c523d0aee56eafe7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h82ec1a8083534183991904c148a8757454992266c858601b3eebad25c39b796e073f6181a0c11876fd7f10b7e6e59abaf3ae48251f98fa97436b78b5e0641ab8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd13544e681432020eefaa93be93aaa26993df662878f91faefac98f32a5b3a42a7b898dc27c8c6b6091a20dad4e9edcdde462e81ccec76f8c35e1e25a148683d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf5784bee62ba909274ad7c624eb641a400d78d660262ae42322f1b20c7bba69c957990681cf09e8c1999f93233a4e283749578c6d2db0c1abd9041dfcb2467fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h73388ce879b577604e6b608b91a38a231c721d13afac6ca45340b3141dff39dd75101f9e8cc8106caf40d731e441d93ec097451a2a5cd7235a79fa2363c97b10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd7bd49eb7a985611ac393549b542f7840bf8a27e5fa8558703a4aeeba89346c35546a1d25b092e0b329f6865598947a9ed7dfd9eff67ded34faaed4ab498d1c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8290450170f179819ff4cf4a7484e10f2f2a1d76472f2c446a094b0ae10b39981181c68616046bee15700460dd79b04b3be7c7cb06bfd9be1c0c8d7829aa3668;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h14b65e5654628e890ef77334e70c0cf52502b296c174900f8d3127df0594daf9da7a1dbd51e3cd301a1088dccfcefd0e559c25683fb4d6dd42c5b6f64beedf42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6cf43cbe193b8c6055e2b5b14f39cdda654c1a53c40886bf78700f8b0e31459e6b786571e82f6b8f67a3ce12873fd4da0d34173f4c0a2530bdefef5f3e952c90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h37b5bc4dcaffe5ccb4a11e1d5a1cc8630cdd3b536d1675b1969ab3d56bb8a66bc1078030687743423dff3637e5af603aecca3085ec475ecea61502caf7e33e38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h91d6ad3c969a4742efe38276c64bf5cf6c5f37ab90be60a94022025db25076fdcbd5d22ffeb7050b138429522be75dcbde00bb97a65cea66c7e88f08043494c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6c0d97cd493f3d0f5a677a9e8e4f60b46712292a3edd7bb0668e8a5d9618a0639ea04aed9cd951e46a90d3eaee72928d897fa7903f6b37f365fe0d8df61ace7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h536a0e55303c6f044c7204cdf8ff21991cb11238833db7070b118f4e5cda283640ae74579124542ea082f148a89d2ebd0dc3e516c89d2d9a0b82385a1be23051;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h62a6340178e4d9c9f6d44536065adb580388fdd08c1b4b036f186bca1d883117760ff0de73537f33f4675081827e8ea23665fb8e603e3ec77d05d7aec9c7b1c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hddb0bcaa1e7e7fa4d34d34a7ce78b687468e7fc18b1204109c5ff5fbede8db9043900c13f9ec98fdbe34d01e5399075153c882e1a299b26d8b1f3483ff6733af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hff88657a35ea22f855f827ff4a3e6082046de41f7fc609fbb856e678d9537767183431d370aeb4acb11592748a81bb3316649c42293bc180f8938651ee07661b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1f49fa5e6a13ec6e79c3a979a762d21a45530e414f2d26899ba7c9fbebb97e1e7bfa497faa044a9bd81c9356b01f0e6ea107575ac08fe173ef95645a0bf34b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf5d2e507aa3bde08028db7f48a07c6c6d1f7fb20ee9e66b6bfd3360ed9bcd65010418d03e3cc1a1218540d09e33da33bb10dae2d705f5657ec932a67e5e8bf78;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9c33a6bb46256f7411964e506e9d86f029827e0f7b615eeb10d216b7c35ad375afe87396dcced2ac6403f3ca5727007fd92342ce96dd0255295eb414c7f11bc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6401b07ead7da0b0d50bfded87e1bc29f4e4687a8c7d5f8d33222a4e802bf3b0867caa9040524c564c18c9f7914221fda71efbbb254cdcbafde2f1afbf57e445;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb809d0db43d5e1f216834d8f5a7c4afd237ffbac006dd78fbb0451a332d5ef9b0a818a1d8f447f37e193f7f1c6f8dd829a1dca109ec9820ac27800c1d3942470;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8c94d5ee8c7cf7daeefec749ac23621e331d8b100a168ac710789382c5fb8b17d8734410164517ca05d5595dc1d53831ec06e38d6aed49f842e094efdb68cdf7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8733ddf7c3b620bbf24e69a3ffd83c0a5e093a1fb078f8afde0bb30926d925b6e930df7db850a73591ede305d20931bf053bbde5cd74ac92dabc30e2c0505979;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h83ab432ec1b43cdc073a7d0c17dfc5f58a35030df2ddc23f1e7cfe638f854376bf364715384e2acfc561ee57e117add3c81a28e5d07a164aa2602e9e381c1901;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfb7759b14f2c06538db970854e8b00c6bddad7146278e10c67cb2ccca9589a7de1be3d5ab14d820240031fb356961572bbad2a5df23d693fb5ca493c34625365;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf24fb5091a01a41ef7a92c1f0874cd4397b1b293dcc2ae80b9ea4db9854ff34cb5b464a004707411a6ceb88378c43290eacaac1e0939f4637e924bfb6fb01fd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfb73c0b291a9bfcbbc359664760ba5a71b512dc5e7a6de3f9855c9bca3d8920c7dc575450ee003f6724ee1c26d2139af33b9e64dbd3ed322ca9c3dadb70ef7d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h83268afee645098c74a66751e3a20c288643fef72138738e19fb19df100921251a1d3dcad3f082a7fd03c1d1922d878fd05b1d49874b6336da419a70178f5c86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6eddffafff7cba4c3385693a4d7a30d87f1381b150dfdbae3f56e678c82baf404489d24b52dbbe48d5a477df04ece3a74894aefc19ed4f5448a5cad15ef85c0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb921d34093081c50075ceef09432c78c93252e73e5358eff2e36ad116dee78e3f1779e953f58af2d01d56359bdbc80b3c10e0dcef0d7f922984d162fc7127d0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb37b125d6333d2fecfe2ee523b8e9a94302b5777c2395d6ee668a01a4877308955820f15cdea526a35340fb2911b301f172797aa4174d3dc649cb86b1c907526;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8708ecc0144f5360ff3c143ffcd4d03af1afb4a2db1a98176c4bd4f161aab2f4d3224d1d043a395692ff13ee3b6b6577442488312d6e782625eaaf4ec866b2dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h520a9f071cbf6a341840ac26ec7bfe39573fa3e22d437c4661a3e6fc399787cf38ed4803e964fb54cfcdd4b1554f64531dc046416e971fe2d4a918c01918f1ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he86b92553584906b673ddaa86bb75d9115a33d7439132abc070438a8fea6780c5001b7daf485603aebc90723ca227ed9aa55cdbda694555140754450aabd07e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h463520f8f2afe73efbae3103ba6a80772e82c51f7b6a117261c982e75ac01e3f046e7ecef38dd58828908dc9a8819f2ad72c9c3660a095c5c75c3d16413856fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1a305c145b3a3863533f37782c3092e16963fc952507f3c37ce5e53e868d93e64ddfc57ec931fc83028b9093b613167e797633fd5b3b06cac1a3688067909b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h516419886e709482a251873a841b8c78911c31da0ae17b0dbeacc1a6af1419fbabeb7802768c9ebe9e19ffa1bfbdc077108b3c5e4cd33f2aba45a841e8a4d5f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2f2460914851ff0031a5d8c13ca99cfe81c452d463bc9cbe201cae80a6e63225e3daf07d457cc0afb2ba3282c93e9948f798215a3f1d0d8d7799641e2f208c85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3919bf0c3599fff4f9ebcda7e43f857a1beddd60fc95de7b777a844615f88257de72dad4a08338293e91421718a5b88c293f32278d617e953791c8994c84b988;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2710913549606aff32af7134866e1b6b80fc50f80687ef0a538d560300924889af9d7176e6a26cbd1b258835ec065e97641c9754400389c646e6f41efe7af63d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7ab63de56d742501703370e984b7a11a16a775e500bec1592f2266cf0e7c3e7dde0ce02f04ac477cdb46c9ff6602409fdd98d2309d9763f34c36059c685c7d49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hda8c795b6d1cbfd866129a07d123fb0ff6c82151ae36ede69640b8272371346f271f4e2a3864ef925375f720337ed2b0d077a9e074e83a9738e13669390183bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3450c27f3e90d976ab7e604a7c70c9d87b0d8b6f4a109feb59b581ae1dc327c575cc39db157b6e285ad2eec1584488d818cb5f4e35ef151c31d73f4eacfd025c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h15450c4bb39d9fe801767567342e263bcbd5aab42548e26c507dcac00c200e1c08b963a7f83a61f5b161f288ee524c8b4f41923229d601f342c80dd0460b071a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2c8dff51372d2cdecd9b0c96b3375197e56f1596ce6269e89e958609d925087857b84c5fd5356c4ab11a456f2788c9aa6d9ad52d954e68327df41ea3d909068a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9d365e0b8859d762901469e5d7a180a7c454daca5f3d8f1fc024e268c60516f5e5143714f7a328a20fe3863d6933fccacbf6d8a87499dfb12aa9fd0990fd108a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4806bb24ec2ee5f77183686c239d3e6f0b803bcf83e99a3a8ed2ddd6a22ea996bcb6a590fa28f9de1cf605a1eb0fd06dc0cbffa9ddba4cfc9cdefb52eb1c76ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he2b47856322981c01fd90f2184e3c4203b8d6cf42b1579320c576acb4f5fe39a17c82c0076412f99a2d050b9c67ef8b460a04092ac0f4986d0c3e592677ecc82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h22d7cef797547f81f336d6fbc634a7202d2339b60f8fab74494b04b925a6840c130a4a468e0b08cc4a85b9f5710f4df0c136a0a95476684fdaed0ce7850d309;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he468d4f51bdceb5abcaa2d579013a7132457257689ba220bbd1f5fba2c26792600f0159bf4eb45b87b43d14962576b10f8927ba266594ca44adc8953bcbf0027;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7d0aa3e3c475d9f165b2ef5b222d45c14baaac05f04a7ae6cc94f5d8eb1f1e701c73e73b46509a45df7ab2a0926a52fdfcabbf69297e7181fc391422ce5e76ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4ed7d32e5427e92cfdd151a4e037760bf2e0e39b8d9bdc920dcc3c3b96fb1966fc77c69b6198ef545ea91fd859c2b60852f3bf10ceaa6f4d7cfb589b5944b8fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4583d09df78f2999ee99953443194381b0fb0e90c978c9596c43f1f0be4b1f06eea4759d339439236760b0a77165566d2bfef52b400ee0a0cdfc66a190e299d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hbeee6bc740b4bd2753703b2cf9c87a124d11c491f0d283f9cba08632a1171b2ebd313dafaada2206467529243cb1c4dbfa40b6fcf316c791b81906219e047b57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf2fc7d1234587e1559b28bb2a59dcb45dcf7b1951a8dd9abb88f0ee27d0fe9686ede3fc9c1fc20cccce6d998c6e30827cd75e1ae0f91f74f4ab4a615dd2bdb86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc0b6fa0c4dd5b1366d70004461c21fd858c8f30188d4fcea46578ca658e56fa49d3a9035b5613f4269f13de8a371a000082ca139cddb6a099bf806cd65b80336;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdd98d231ca203206cec97291f113cc926938e843863a8328c17efdfccc466ea3fb23dccb0e17cff7c11237adca12ebcf9ec98392a0ff694877e85e346f9455c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hefed7f041167530743a94daea46d4c90d5959c0a6d8afe733e93a8ee156db8d3c5bcec97cfb7981db39cef716ea9ef95ece9ba6678b8ab03d147adf68b2c4e40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7cb9e99136ade62d078135602055ffbaa467a83d37220364411418cd00fc1b0ebb6f331fa7519ae4c17b1c51cf53a69c73c5a85f904db29a634a8cc59e9e8f7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haa3f2e7ddcf33023801564d4a2f7bb7ae1f14bd70a4f4b93a916c692f3c277ee780310c0a4ee1fa1bfe4e15f54c438994e088468831a168212e16f2f146533d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8488487c79f7bd574366d132846569fe3d39e945b27bf6733cf8debeb5693f8131db454a5cb6ea5b8b40b8bd89f78a66fd76b968480216afee46442d15f1b00a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h51b658b8210b5e7e84e12ef8ae5dc6abb6bd7068e7c493dbcb8de3d57b7f1e66c50f378a28c38f7d7a349bc811581f35cb8e12f159aa9d2fdf49c366a8371c53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdd9b841d87e201490c3da50a9f976e4683ad99bba7a7692de60cec77d13bb1a02c4e8e9d224efd6fee2bd9810f45caf129f6dbdb0dc319a2991722fe87695cb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h253938fc1911309083cac53be5d2aaa301be2c4fa10f7dc05936542151c33a9b1a31d47fe03b2306d5db0eda874a54159aab1d6be52dd757d018e45c4944767d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3175afec8c09517fda783cba5fbb0f30a5a485d0693e1107b5dc8f6eec20d60d20ad22aa4d93d41168953e3abbaaa5baec801a874b34d5af97cee9c560b517d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6a0a96afeb87fca66eb0bf97df6f1322e52ea5000e111b51503ee74fd77d809f7f3528d96f9fb443d3e753fef96ec9bb64ea42085b337a3526d8f9f818eea7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdb2379033b932908102d2e049dec90ff5130aa528d14f67250b156559c9f852f7a33a38ddb3fc8af90b80ce7c445d989e52866416eb4d2cfed427151b54ddd87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hadf8fc79df019786f58925ca0eceff9067c0a586c22279362f99f577bd360a093248e11e170a09a2476546cf3f27d45140eef5d34f7b8ae976c566a1c0b5bb7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h66c5c517a19ee9432b1d731e3a3a8b64af179cce4d5d1d6c72f2c16322f6483334563ad31ff8ec48f83318c23f13a2c5edbd65e0265f30099f47b7a10f8bab1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h88b4febd7110f9ef3ed63044667d4bb13a6837d4bdba3fae4799c726908b0efd48a7548fb3541b8309ada3680a6d487e822c1630dee6852a442b4c9087fa004e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1a0821e75d6ec4e780b3902c79a96119e3639b03c8f08dd63464565c9f85d9685d742d3df232aaa10433c39b1bd7a60f7b5e6cbb529ff092936bc1ee0bebdea5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha9c24437f3579c98231072375b82574241e8fdb3e01aed35be2ba7945f0d7be260d2ae92c9fdc311c147274cc0d8401daf036e5c80128dbaf0d737b71915e60d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf393d890fbbf72554e4a4305387dc2988429a8ab8d4da3114e4e87b61f120ab9bf565aecc19be19d56ccc12cb0128cb9f2a6db7409400dbef9c78f93ecdfea77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9f543d78da1de446d4819db4204b23060c745bfad2fdb7926c069cc5a4c6bb43816caf4b73a99edea997ed81cac1ab9da3ad820dddd4435e3d3fd662c2889b3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h81e28ec9188b46e1d1c10282102070e842ba716b7b45ebe04d9d9aac7bc1ce7d779081d8eb4181a57cbdffd5dd814098ce90f56225ade090b71ba0bf6c2133de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7f3fe3c8ccf0569f9fba2cfd5f629eabf316881f53b8bd22a4d01efe858d4cdaf1e98f3b066692697e8e15f4fe78ddcf2bf60300ba779382020ab38e745a8cf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1bb693b499da809ad1286418739a76752431a60ff35aca02077bf8ef1725e663dd6b7e420d800704f6b65af5dc0c73e47140df5a15b6950e5422fcd36dc885f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb55c7d109832da95eb91d8f67f0f663f785c95be436d7d8db7f18f359b65d9c7fe1a2521930ab6e076ecd681392114297af90fcbf0bca75665d932f10d8e5ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2bd4bb54b0144f220cb67d8373884a8ed0c6b2dcdf3c35ee951d8945af3410777dfebf8897fc280c35cafb64451ef08ffded34a2369f843211e5bb4cb8e3929f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h65689c37f32add481a0ae21e67a7c62c89cb2bae75f9f92bef212548e150002398c312615ec901987f84ce8f30351c4fd5c3710ae10d203046073498e21a4755;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8a9c494f1490158362b95ecb99771186116841fc764052eb0b5ce137171193430043431149cd96ec2e5cf2f1b1583ed07c9615657925747006e077bfdb540628;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1b1cea71eb864da85ead9bde015363250e6eaf4d83ada5bd7ff2a22edd6b70e3df50c0ddbcc4a481a46125ca10fc2d93c178d75fe126748a4d67e9267107fff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7c5d3712e3078df097cbb45ec1b8952b935a3c4ad10072f0b144f5979086ccc39d92bd556e663383894bc29c2f36b9534440f25e7b6b0195fffd107cb3aa8342;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h736a96c9bece25a2682187d42e22f89150f5dda7575c59ba88f566206827f0136c8a3bd401d5aa3db930b024286d8267517dd300d6e2988980a14e9354afd739;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'heda43551e52c33b81736cf26854b8fb1784e4d0e12e1ded23ac4add3c54df96d44ad8d4a6cd0a3c8f233a7f1589ae2648ce1c498add1229548e17a5d64048b0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h119beeabd19f2685650b9fd91420c3b1ca0205cfbef7c80a0481b7aefe1b00e06681ec36431d583a8db34b14ab0c67b3df09f3719f0a557ca4b247c156fc3040;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h64c74f91963911753d02757fd69da553f44427e5615218ef72c45fb95f09cf602dd2b8534dc9163a72b0dc762adf4f5e0f5959535182098397138a12d7768ad4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he188f1304151e6b09d782d68ab825d9bdeef1d23ff04403688055a286d2cf5b4ad8fc403daffee183cf0061fdb0e1d34f2ecabcd3877acee97ed511977a885e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd899614ddeadb22d919f5a3498536d8ab846696aa9fc94628fa4114439ebafa77e82675b96cd3f2b2ec247540ad6b2ea1f165f9e4078e91e19c76225dec2046f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8e13d14b392ff78ce0161d6cab754d3155341877feca46ecab1da44687308f783954138a9e03f8597be9aefbfc83077baf648d29fe8ab6ca8f1d72a9b3660b60;
        #1
        $finish();
    end
endmodule
