module testbench();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha05d2452668466ffd1d49dd55ca08f325a1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h305a7834f01e84ecc02f02957d8e64e8900f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1a0338c399606b96885cb8f618e8fa869ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4998e63b63037583703556ee22b0433c4355;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4786d1bb07fbf712ebe382767ce408791fa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha208c7c4678758ff55c5a520eb2ccde4d65a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6d0bcb4248d0fc25366c9692c740e17cbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc521b0bfaeb63f923d73c9206a12ebeec97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcd7adfeae4975670971bf9900e4cbdc2f01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9722cc3ad393e91a46a9d8a37f3b9b63da16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc00fc51bacf32a952df1b38f6ec1c0bcb98f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a64c7922f6c887e320bd582a5d5508eb527;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fdf3a8d51f10c33af895f093b8731c393c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58e3523578ba4579133fcd767cd4b15a972b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he09cb6eba10a060d608c8354d8614eddc95b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd66fa0c9145b637a2090bd0a518626987443;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b518f61b965da1616a08baec047151f45be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b142965bf8479eb45de693b266145ea359f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6df21856431106828cd63326e60b03501ba0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h427024779c1c33e6bb061face31e81ff20be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b06a922e76f6c72471196e5da45ecd216e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16d77ce4587acf0c145b18048688a9e65fec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85961fc87f10380720aee3de4dc359960986;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3822ab36ac1137516530566a566bb24d2e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb617fa5b210be9d61bdf07f67494e7ca7a14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0385cd3787f286f6b894a915a41d144e5ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e4743980ac6fef785209ac946e9107d02a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f77d1df74c459410e97f0a49400b58246dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63072a714aaafb32f0ee1ae3f9c3b76e510e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6af78fc2533c6f67cfc30bca49141a907507;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ffcdf5a3ff4a5bb9677a11fdc4e9c70fd07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf34ef0dc1bac53c8d60043b48525fb21e12f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb31eb35cfbe5905f14ffa68f525f667cb935;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31b38adadf09dfe3744d57973b1486bdbf39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94f52f7fe3df39a1b84847f653f6453af05b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf4aadc727a5bebb88c8c920cdac7355623e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a0bb948f58e0653b1b4f5ec05d41ea2489;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heaaae91e9b03434ef44eb1ee6958cbd9ae34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7f607cfec59e1337a9e5f003cc1df11b0ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81987df78888f6b8b7f86f19e8ddc4de03ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44794b6b1d9ca062a66bc0c6e875b6efc915;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h976109ef7d0e3ed1e572cf8d2484987a9439;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0134b43cdb84bc8c590175e626b5db854;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c6e5a0aee7272943f98ded22ed95ddb0647;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8a4e3d49bc46530e82e98ba52be06364d3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h683ab341f6323d8eb49369e637665cea27cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63d9096f78906891bbabe8965e8a66c6fc2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8a41c465ae0f5401a58afa7d01e17250a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ff1ebcbd123e7abcd16930eb77f1e77d909;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac7b7bec7794ae213495e93f64d8e5c53d16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0f51120308cfdc57def39d19c6409e7f7c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h623e700141ba362bdbe25443a626c0f4b345;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb34ce7c4afcdf532c7153fc10eb8e66ba4ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d44bf02e0cd631972b4989b50bb89b01280;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38580c22d268d2040067155193851400712a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63732d3bd09752b3f1e2188a149092867505;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0c50e7cd9132b453a671902c6900ef416c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1507c05a5fb193fc1fd1962fc6bea8aa75c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f9f2167858d85f1dcd16abc9bb52511d948;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae23131225fdae0023aa4f2cba044a2797b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf42cd5d1a3ab3869830e87e349fb4ae10d01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h942f5ef85dd6ccdad5a6af8fecbcd4b2b4e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d4de10d2308dbad4fdfb7f4e106a97ba39d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3bc76e32ec63423b33e96d3330f3100e1b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdbec2c9c62d99be6f7433790924ebf61e68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb57e9837422bd7b97e51fbb31652305c9b9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a2f459d6e2d86a3110f52c29548f692520;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae8a3482e506c3e02b3c5c733dd396de9368;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b484cb5fd29138b272a7d635c942a9a6a7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h859ac5c782aba85bb920b3837e0c740897c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h556b8fdf0ef74a8f3e038d2a78572c2ab01e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ecc5a17edee5f626a6e8a189c6934047ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b10735c4bdc385a32479c8a53d18ac7e241;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1853063039f9c5a1519aab2c7bc3a3d3b9f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19ba78f74f9975a214b6ddd2bf8c89b4c213;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a3434f9c8cce2f2aba9b42b4af41737701;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd8d42f33c91ddca7b1eaa7e624647d35d53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h969fe4cf2d1aa692ca2e202c1dd05e709ca6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a751b7cc2acb0e53d0b5a0fc79d09b3f694;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbedb90719934af2b61a57e4412b4e0ce6691;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33a2cc5e759f70d69b9fbcd1b2eae53f7b31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha57d88768925d9598d25553f86470f3dcbef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haff6965c235a9b3c1aadad2342cc06a41056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he18917a1e2bca32ecf743c4b123fe402ff64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73453cdb1e26dba31b4bbde2eb04e1070db7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h883ce6cd7df83e9b77cc79ba0e8a600a19e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f1ee8c06f24a4a8b3bc998b9903e7e2d8c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h604cc7e77ee4ec2256de9c4fd39c6daa8b82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7df8b89ca1f4b295605f7f6a6c6f1008ae5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h461b68a406679649bf9074bec2adee1d24e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1de10a07a15e2efa9ebfa7aa9f15a47b3721;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ae3329e9c0bc84d3d22928d04c0c81fba19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2ee921d13a3b6f147faa17e49473753205c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94a5438f6e5a80ef8ff7a76939630153e3de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32ba0be8944748973a94b3aa78ff3876ec8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b9c5820dd648208c289fcf0e77f197914b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d2dde30c7490143b465045163ac9fc7bc17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5da5f7cc912c35bb8fc6aaa34bccf362b702;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f0fe6c0dfb89e4c637da82e6085e5d2fb82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd957a45e22efe007e6dfbd8ea174fbaf8271;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h220659873af4f56d6eef73ee97cb3fb91b51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h814013b916124f6bd4472996d838800141e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7d7480f002dd67e8831bcb63235ec4f585a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7773f4c1ede026f7f829ea09e1fe91dbce60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8014f9591ec54a6f79f374bf032fdf6ec2b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17b112d9324bb5e6d3a046f97bb236146490;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6502c7d749858cf71ba2b8467e30240a76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0462c091e3f875aad8296440b25d4d94239;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7825967732eadaa9709adbd925a3270e65f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6392d2ac819e1eed4b1671cb30b6932a0ef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha16ba50e4d4f1e06f89ea3411a2b5fdd7c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3ecc17d7837ce159c63227b9b7382a7042;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9974986aa1ce010e70df257094f21bca04bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fc8e18fb640cb5c7bce535a110404886969;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10e6e3316ad7639d8b1018a7ed8d6ef93fd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf55ab8855bb6d8cfc1c1478e16d02608ff4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbb53e300a0eaad2186f36deff25f3f821fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde1552c84ac639ffba9c70a94cf7e4fca5eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb077ddbf5fcd1f91a62afdbbcccd8a3cf60f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83a2f7a8c79a6c19bb0c765333cb499ed0bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c400cf5b6c2752ba72d2c0d93d91d4f4ce6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd3759f1e56fbe7432281f8022db94aed671;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h344419e76f39cd82795a9f46b34257915b63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11f8d26ffba5031178987b0f09a10a071d37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90f67d27e9b93fbd82de03f8411b431fa705;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89bdd0d8cbae9618f0bfc45e2c88d35b1287;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1f44c3fc9a46bc739a9bb859023da237267;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h514a92b553f849201b086383eddbdae53274;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h211d92d80de8b85f00e8784097efc6fc3bad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab169f2d510ea09c51b9a32f117c796ab801;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69c374a372141630dcddce548e0f9bea2c43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bb5b26b6387f048f83e54aa87f5adf58cd0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he21d28df2437c47c4597b75fc65f6a8d83fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42eb206a9028a10cd5ef0cd1ea55fa7685b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b0e516a266786855e4bbc9b72c4eda0b7fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e76da4eb895c8bfff2137da60bca1eda508;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf24351a66a9b65b67402320074271349c30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d6b9cd0291a8513c96fb356aeae43697b4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9e663c4650fbbe85cb4daf54378d9b74062;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae847b37507e7e12b557cdeb3053959f83fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6460b6479b9a5606e065eb489fe2d311adf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c2a4f48d4c59b8ec4a13a419bc846e33830;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h504fee98b2d772a8b5822b2a8cc3460d63c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h603bf86a3362f3353f6896ba9b4d93118a23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h559546ee34ebebabd9392a420736d01c7e05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5622868adad54b696a090a1274bf244d0b52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h961db1e60537fda201f5395c4e5add3aec5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc29270594c105e603057f61097578d3c912f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h958b5cc9ccdf9cd6a1f6d24e1b3a034334ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha051b629e78605fa0ac70b58ea95e69e9121;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h537bb0b6dd3dc2e91e78f4b53f25a973b302;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5291c9838ce7f98c8f5d426cfce85efd9d23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed17a44085cb2e9f5003ee22a4b75d5df33a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb48032a426b9f859de58dfb4fe0b0d90280;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f2c8f1530bc6397c9a30ae874662b4eae0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92073f14be1eed6c5afe496840358aac7971;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha74231eb2cbce01bea8e097d7e1601571fa7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h145f68a6ce2387f18a3d028b942b4abf612;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58c6c529c40df4b48af0cdb6da401e4c255c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha23f0de2ea785a99e1bf649cdfb28cde9237;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a569484f16080b323aaaf5031444104cb43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b7c36aaee26dc1439eeae8d544e71e190f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25881fa669314a6bc8279aa99db20658f0a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71097124c7685f4bff75e27080a8ee355f48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ab04646f4af6028cb889be4845fd1f84664;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dd70d3faf334524389c577db25452362171;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b2a35aef60a645da78633f5551a56860b28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1279a041af328fc4a488fb1337c739d6d56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7570cce882735c4340b5cae7b21d3bbc9a38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19a40e8ac6a3ee61b2aa09b88aac9939dd5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c7dc42466db0293e9aed935019ec6dfccde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e42612de6a4755a1dd2ad60f1709c18453d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f669af5e0c269f3eb76962397f154f571e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a388acf6aedc9310bb0df71817d773a7bae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29ee8cde7185e66d28f5ce93e338e7c913b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha542af399913b7cb358739dd108fc39eb7a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88f0d2c4527fdfb4900da80f370d3f45e012;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84d8e3a86eb44695fe3b3879a6b829806071;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26f48b8bf08832a2dcf9c778d87bf95abd16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h573873e79a432ab061fd64b83670e3b9b69d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf925c8c392c30cef0ebbe5fb4a062990bfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h397157fb2243431bc28e8bb7ae24308c01d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf111d8778eec575ed8b87db7dcf769918dbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5e11fdcf3def61746636f51a1ed7efd873;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a5cecd08e0a992a960de3baa0822d706c71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e9dc44530d4170afe3466c35d10b0c45df6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca71a2e6750f760f74a39a3617cd4f425a84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7cc7108b72f80d2407aa1b4880479ad8dfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he53d3bd970494a6a54b4d7c34e3e78c4254a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26e2e41e2004300c3cb41efc870469c4d21b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ed1d6b27a9aed9a3905125dca2a493cceb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b9bb1993a5e38962b09fc6bfa33e1960bba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9b7ed06ffe590d8478ef6a6bf71f7837f87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f03d09cbc19cc5d66070237f908f49ce262;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h646e3a23f6eb183dde6044aaaffaa2e715de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a81ac97fbd477edd75f5469978bcf0a9c01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f6287f84a2a7b62015bbdda2fe26619574c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cd6a5421d0786a456f3207621f4e68fa789;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c882ddb99d2d3e6db1ce3f83902a0b4e6f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73c3e1c20413877bb993cddf2822f319f5d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff0916d1848afacfa35752a5fc49e411a3d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2556f8e9ae0edcf80d64e827c9e735a72de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc49330fceb17360519df411b25e5268c93b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6f6f656239605fcb69a3a76b5c2459abad6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc239b13ec40b9d01041e83cc6fb2d162c702;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6926198bc1c6c0e6cc090030ca26ec70970;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7590a683a038650eedc1ac78d54e826b720a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1328464cf2c4d66167ecb545332e0ad03acb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44e501be788694f7b9a18a342111f09d19fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8e8b386eb7a93584d1e472d42c6ab52c18f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a1c2c452a6c02108c8dcbbb05e2736dfb09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heabc1de3df18a500fcc281a9d264491ac6b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4649b636cae6bd9962fb3e33946fd6cc45d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29f7332ccd04b096d8498103ed56441061cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24bb9708a5e2854d98b56400aa701b4f246c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4516946e1e90b065cb6d392f367542ce014;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb167d27d0e61571391a2fb5b9b4aec47d7c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bf0f2645b6a385e1fc54e7364a890ad1852;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbff026f6670341a5ee85619ae9c1d3f1c8a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h237037cfe7059155d1eb581820ea0d78fbea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14ad32a2153c7e2d913b45e2f1b063007dfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17b39b0877aabea07423f69e0e093887658a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dec7fac744c77405d6e418c0692e47840de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf629066072c5326274bb869a249e84493448;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf0674944920f8b6646382d9249d2499b957;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddb2587e097443d34bc4d8c1b65da7f28927;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf3e22912d69d442961fc286887c998f5a49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b49c3bfd9dedb408104126c9706402a5350;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89632e5aeb16dee8490382623308c5fd41a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c1280fe191c66a9e52497e6d980188e89b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8aa06cac814c970c6a95edf527ca1b19c65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf12f8aaaafcb535345c7e8050fc2e779b61d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h956a24dc8eb27913b4342b5f181afec11d08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66c6001d0272dea6daa5c886cf7cefe5456;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd01f7d988b480cb4e50feb717b7c4d0dd9b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9178b6d121893ee0a964d4cb8d969fa0ac79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c49c1393189c963bf60a1ba1e8ad9e72bbe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5173be1a815a3c1660f2dfabebdbd2a3b89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a5ade89b40e9710b2720926e9c186659c92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd089c206b6c2df2bea3b8023e7e0295f705f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb447ace7b6de604b18ccf915dcc754e97781;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1156224a6dc3d2aafa1c1082c014a0a8ce8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h334b314b1a05b2ee6b1adf6e6027483cc9ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e90fa1afa6a1c12c6617fc7e2b6c11e795b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9472f66aa191a4f1e8140c82f59a5e5c527b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeea6b9da5ad26837eee2860e35ee240eadd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8469307b5e444e8b2e99e8875f296c98f0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdef55bae787d659fa172805058eb9473a838;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha755899200a546c288b5c0d414e7f511a577;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h701c61148abf2491aa64a7b2f42e0fde850f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h549eab762c66034df7f24364583e0a77fba9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha667396556fe82de9fbe14739715762c978a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd55d592678b348212113f0482c1df130039a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a362ed90e583217e2b53ac3656bb701e1c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67cdc9a712beef3a1a3468ccb6b55dbb2923;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ca64568cf22b7ada62e471c2e113580ab66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had65d5bc5a7ab8d1b5efbe6add92436c2ae8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2711e7695abd565db76ea2773cd76efb678d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e10048b95241da8321e97bed9989dd68929;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cfead2be4aba6fa74d84782daf29a978608;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8abc0033582bc73be68f38d51cc590f0fae5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf921ad38fd0b1239cd6df5b81eac505ef0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h560a0a6681818d695d92b5a74e7fe58a7c72;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60a25faf0e6bf983a99fb13661cab4e68814;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7226f0030583de9c56f665b4dc4ccaafbac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h272a748c2304276c7156befcb39b245c4df9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79363a11b324b86bd9ea49074d56cc6589b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa3ba4f383cabd928703162c366658bedf45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18afc096ea083169dc9a3ab04ef27b983376;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc55b671df09d20f5991f013008bf446e85a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40b5a461ad8fbc69bbc765980a02c4c82613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42ec5aa17020c6715b25363231e457884b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0e52dc578a390b8c825ad341d068d1c8886;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h517d1bc8f055ce83d00fd4d849c84e9aa4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8faf542cb70401a9e8adffef046582f6fd4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff152b6fc82b545306e795cbacbaac6466a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d0acbf108e62796fea85d4da25bb1451bc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef98190b47658d7a3b8022fa95c904480f98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h130d0f494b4226616e1d78145352c0ce895e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddddf3bee74dcd7fa2648ba62d4332e3f563;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fb947e20eb9ca798c9b3ad7f59bc384bb9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8474e51441e7fd142bb044e99ceb5faa2c03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e3c5150269e32e00910a46c9e564452a928;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82926ec693323649640168bb4aef9d0422af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49a0e1c110c44568edf2bcc680ede1669481;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e39ba27b74cfd75856b471118d73b3a7d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h344b3b27955d2375328adca93d628c4b3740;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he011b1959ce9c0ef05dedeb0d90390ea2f5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cb508aeb4775f37bb6cf38fbf51b3e008b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7842901aed9200a834d0df0ebbc02bb74f83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f1ad895ab78f2cc353607e60a932948848d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fc72bab4214f91745db0498974989790a9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h673f8e673f602b22ab1b2d5afd7c654533cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9162a38c3751610cac1f5f3f9deef2d8ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6900b3bf1b4aecd3c03f54696d6c8bf011c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha02bbbb0e8b944e254be09280834b9191550;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2ca0cde3513ec96120c82d4ce026e6d50f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heed6c33e2899f4cd2c5ba4264d30c34ee0f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h912d383a940b000b7d48377ca91ecf9702a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haceec8fc477c45ba64c77c92d77e6256954f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he21528ad6e7a70c4ddebb4b734df45b30945;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c3a60706ef75e7794da05bb9df4fb5ddbe0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb23294f4d67e8808b6da74a92cc4f2abd247;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3fc1c6782bae979b24df8445a2c63294b7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha119589b3a8833221c7774361458343adca3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h420044d738e618d05a264616cf9387291582;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h160ec5edf13ec3adb84ceb71a3ba4879c204;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae9d6180bbd088823c320532ed491679cc0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h675b13944acdaf8911dc693885f0bca2c9b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98bb58aa08d299f2a8a78331d0b9a62c7789;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62170a2d3ca9bea41ecbe61373c3b832f9a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf307ab8d7f82a9896c13c3de449ff31aa4d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc2831a38f15452db63a752ded27c3c00fef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd12c71295dde56b9b74abf699345b0f114ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea3f3ff8840969575aa29cb89492ff569cd2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeaabd55cf4e257351379ab1ee1feb7a8fff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8cf4e68d9c5136843af71ab795917375d21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78b07f4298b8bf40bf094b2f41054c18ec83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h885e182f09339349fad9b72d80daacd8dfd2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cf540b6c8b1d4c4805eb7d2d29a50cc5768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d04e5deb303510109bbb64c155642f8f6aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe58ab27a10c4224adbc90db8681e2250a70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3972ad8712b77ecc655666d232f3f27eeac7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd256c24cff1fad5fff83a6776db40c2cd2f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6e247eaebe8e1ac39149fe388e1057868dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89629631a7a47b0eba8f1dadfe48793ed8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ede2e75dda7ae07efed874600e206b6f728;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8abb7eee35a23a0d2817649621610fb692ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf713ff1a6fb8840cb05d6d0401ba9e79e9db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c8d9015ca4ca38c116ced6bd976852acd24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3796c301ce16cfa70c0f0a909aaa5d4a69a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91bf26a046df1999f70c871c1324f7c1b234;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ccb14e0e400a232d080ad64c271d2fe5cd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9207ae69eae62cf5fa5337fc7e010571a71d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h437915f1115960e268d1d39ba8feb61cda75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40bb977a65b9c6dad19151b8a86a05311be6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd47fe8cd99493f7fb96b92e23fa0127d82d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60c9546a131c78aeaf0822494492fd2283ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd595a6127b667530c75828e439463ae4f5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf41189700b109636b3629967a32da21db9dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97fe22498028b6f94b7f97c4b5de137b5cbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94c558e4e0405daded8684357ea3747897d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c1dc6637cadb6a479c54666d3a426779d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf08cb4ef2c0c1683510913da278ad9300a44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92ad10425e6e19fdc5018ce9c7cc2505827d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h496ce0e2c65c594a944a0e8fa4902fc7d694;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac9ba80355a52224ba4617881afd050aecfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93ad29f0297550037ef3f8c932032967b2a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a1a3fcb1e9033f8490acd8784f4c251ead4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee7ada7b1461d0518ee91f6b2b08f74c16f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4aa1176c72af1cb8d08808b9a1440dc3f5d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbb7d451a7d340f34a4620fd4890d0c61b1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a0ce4174c0b38b5d1c685ee1f2981444e52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6782551759d61f62fb41324a81feaafc4fb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49667eae76b9deadfb753ffb8dd4211832d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c4c8d5680ac24a250c90f887a7496bd1b92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h552e9518f3d1e7815a136dfe4e8f4d9f00c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha94d9acfb7e93d0dd906bd3608eb6d5a2b73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeabf429153c6f196ff337cf3303e61c77d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f3f183ec9e8290f3ac06375d9beebd0d0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f1f619aa6d96e0810e11e30c4cf98b8ab69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h795e7f1347dae923212c7ee69b18806cd5d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed35bd88fb75f7bc25433ba8baf1c1ef7da7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69ba579f3b736d3d825728c5d8ae72912b74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8c2e6b2727a69639d03ad451160452ab058;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a92dc4c0f7b50e3bb194b7989e975f4c52f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bf071de811f90f709ad6f0327b15a21eb41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38f923313eb463ccd3a6ade8d76b3c105790;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h592f195041255601fa575d46b8b8b9356cdc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0ac925d4275b5e71da253718ac38be0a421;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ba3e36c5c00e7b663e21e904cc02935e7d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2632a2254a92d5455e3433cbc37b4e3588ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h155a4018ca8f689f84b28582d34cee07a9d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb3ad059f8b17491a9784fd124bce41104a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f4f4db2fcd943f18a234f45a3bcfa4ffa9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h240a14f68ac41f5ce83fe2931691beb30a3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16b43de8cb68e1979afefadb830ec71a14a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e3aafd6e9ea550263ad9128f7c9afe5f33c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b10b8c22210aeb0dfa15afd5ba23d525e2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c2dc00ff963bc854af26b933f2ad0cd5db9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab3e60d9f366b4a31d7e594bd8db96927b35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a74c1f497b335f0a3671d7300b325007229;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa8ce451a94003c24c32bad0e477689663b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6baa5aa71c773d6957e1e55b07d8be74d1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3677cc3829311730d8fad77b52503a8908b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd41b5bfec164585f67d191bc6a8c6befd4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b769e260f6fea11411f0bbe94eb672c5963;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36f51898c8edf64947458d227be65059669e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1f560efa9e52a5a67d8efada8b48a4d3150;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bc6924047e56614cd19fd85c462e360f675;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3298ccf4a2b6e8e1dd7a0f58b5f790d7f179;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he00b8c48db0d20bc1daefb6b477fb0b008cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haac16c43efd02f245dc00724b3e1dd2bb6f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71b042110a680818680bf6300166523a385d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d81f2fd13c3a41b5d484cb4234b8573d65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7881ee56ad8d6864dcc4c541a88d6024e065;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e9d7fb5cfc56102c53978c88292b92a000f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a5f7766010187ef656c83a4292eb8ca8706;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha18d0f14b4408cb94ded3964005a29f13e07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7cbf9f7c259dea935db9c352616080d433a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he15dee2ba1857423c6de523b9f11fdb34248;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6d9240a94d7c90bf5a4b970589426d88593;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6102bf60d7e865af18beb3b58c14a24e2860;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb8e0881bcddb2863614a385590e7800d4cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2fe56ea7f73b5a29cc202f253c3a420ba37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2dd69964a41c63a5ba6ae5517c1cb5f207b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c2a2ce1c3648f2af5eabbf43743517e07ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc83b34c13fea1c59b5faf6e842ad987af371;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf17839e87b338cf48a03427ae6cf856dcd0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4dfdde3fda1793c97314f14e392c8aec9475;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h929d333210bbfe2b5433017285de32db4bf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ca5b79ce80a29683e6629ab7e734f0dfad3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h845e533dc71b3c06257761c4a7ab655faabf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6a993767ec0cf840f3175e8678aed268724;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2afea040afa821bd48a3b41f9c270a5781f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he830da7181d5602a3654b370873f38fb2e44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h352684458fde7ce3df8e65836c795560f479;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5af7a10e01ec54cdfaa1ff06436863f6ccf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd316c50031e1f90bdccce10ae6b8d3d2c675;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e93d7577d22218e25ec11955e091b487a60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b456a4091272fbe5d5bbfdc007cda97407d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec02af25282b68d3fde0b2d5f8f289c5dbdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6970b14547ead7bd354fbf4c1e49d166c83d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87a2eb42eae8377757da87261a0fb9fc6b65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb348a0af1bb6c1be1c1d0e8c81898b4c1265;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb60e04569b4dd281050fbb4dd502d23d9105;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3939d11ac5fe20070e247f9a7025047b1e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfed707e37c981fc49006cab33cf4199097b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc53780d3d00bc0c167b355ae23714536b489;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35d54f3a36523bcea5c1c94a33ed325a7b76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62c79de37c57dacffccc2935aa5b7e41abe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd470ddc0c10c174c71b0236307fd9e601858;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h291ce34db30cd9500aa2e71388d3b52e4ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1214206ad021d6c47492c001152b37665b03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf27e5e364c1110ee44f2c6f1364179f0b4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h971cdfde4dfd0b9bbb69c012ef0ed8128788;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8787ea26eac33fb3d6b0a626fff32209b191;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hceacfa0e75674924786d2a659f80dbfb29a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he46dc95c129f4c3d534158aa63498cb9d22e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb362da5fcebed0106b867b754fef0cf36580;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf740b19c9ad3d5949989d9f86e630984add;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef34f8fdfb07937ec052c7c34a61aa362976;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h895cc74981ef82268ec2469568bc808272c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41a1802ecbd044953f05a1dd6bf5bb6769aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3aa0b43ea3f05c3cf6ed37991a4ceaccf26a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h332106f846b239ef4a92aa73e0de170f1953;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0177e811f94d8d1e5fb65eaad81ebd9dce6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46e65a096ce71995d413a991ec1e0857f4f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4975d3c69015594b1dfa7b445862c5da9f34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c1c44a6da4034341abb9daaa3a4400544a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h767e5ff42b6f7d8517387091126f1fc2bdd4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd4cabf85ad825bd89b0d32aac03829811c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf80a73a7488067a843848f6d5d8d6ef1cd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb052e9bf294db067d2be9d825d0ff39df264;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2185ce301d148636a1adbbe5669ee0a3a6fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38e8411bf490e16a29031562bb50b5f587bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9f3827e28755386aaa1033a7a0e1ee6840d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hede90126bac687d24d8a32bd849f05d16f38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbf893e2e54b4c3cf685b25b82c4d478dfcb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28b0a4094b091768194efa88dd8be49f72c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee3d62d35f2d9fcdfa061af36926e470e413;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea4d6f10f8aa09c53f900442874bc24aa3df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf8842ec92bb82bec70c645786151f66a5c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h539327410f9e8a58a4f4d112475cdaf1c4de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf975b78bef3f8f40770f5f89358a193acac3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35317e768824f3c915faf8fd414b06ebc64e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84277e15b8e6499391dd591ab3a8cd93187b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8d9043552e1e49a23bde5bea33ac3dd5f34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0d9b6e8c0db58239c53945203d05ec2feca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea64de2304cf3e5bd75de7b8fb454dd3a680;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba95f01a86714adde3b159031230734ee7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h731f411109a441613dc074e047e004c45dc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7106698a5ff1952147a726778913f803a730;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb141af5bb63f4576e85adea5c6b12cae79c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc613367192168f026407c4accdf64225c73e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb179fd3ba1d49749d005957adc1f8e760f02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1efdf8cfd244b4aade6b6511099aed476046;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7473c1185bea244743be7a02b9f72a81a3bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fc8b24f8bd389a15c4833607c252ee15370;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd124f0c957ca36cdd91d7684611d3ac2d3d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0ae276c8fe4e8f01aefb111e419b8307ca1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56ea326caee1865ce36a4aaa3173e248c92c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff0a4ac8540b7d882e84daabb6e71db70779;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he95d8ac3c0758d38eeb04c1858a098b430c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9eda6e2b3d8db69a0b0a97b11fca196aaf26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce8adf6da01ec0a2877178f7fdb4b29a5aff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c3d5778295a47577c22d6dd5fd6dac82b91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9721d629e5e6ee88fceba2f14b8597798fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b56a4e608b19f1f418318ea501cb7ba0791;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7c874a20ddb871ef6d812333192cf0d11d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha278c517875124260fc3a7b9b910449e180d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74dc408ec58572400af44267a0d842fbd1c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4ea2457ae97c6d18951c3b4cf0a715ca080;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e180e5bc832c40a88246346207d644ff79f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb55d2f004ac851e5e20caafe22dda2d75d78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc37bb5a1b6c961226243775f8718a0cada4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9501b75ae832ec8bb9e12428f1c4a3b8fa3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ca1d6115c371cad0029e8ef4340884df2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71dda0506754e1f5035fa223ffce4a723671;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d6dbf06b18073843126f48e9fc10c6096db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8efe2d26b41e5b60d0c2b01953335bbc108;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3698495170d2f1e9d9bd76b0f08c01d0193c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2c81e0752426a72dc9e80cda9954bf5934d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6157063e2f568c0df0ce51ff49057c486136;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha60ba32646f08e0aa047fa8ca3270ffd98d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d008d8b0ec94c28682a7637299202af6c6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h570ef1430528c74e67620ca7eed59117e78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea6b0e8ca9d566c67a0652b4e931c734a258;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac0a622bef294ad2136e2ba77922427c9ae6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h189e86e450209af4a45f5d201f3f1e09ee57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h182ea45f9f402cac6652cbab3dd0c7a1b7d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc2b908b227b63a377eb501956b6b85372f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h153d250c0bf56f7580c0093144b3182bf97d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2c72fc6386f1a2438ae0905be28c599fa44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c4d9b3039a9e2ec43c867b01cc1ec2f2352;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62cd35f47d75457c482675f6dca0a5e69ba7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6d0d173e13fb8eca440b0b560371ecbc907;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcca6189773446a039f5fcbb14a5b6621433d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he805e80d94476ccdfdc3915efaf01ba55724;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda7d5900a12cbed8f9d6ae0c6a9db6ccfe00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3183ea28f2586680e6a9ff542825d291bce8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h797bbeb1f0ade383b496bff1d09dcc51f1a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha68bd452ca59b47fd3d5e5293c42611cbb3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23dd3f03bb0d7f54d34c95f3c8b9a23e3116;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55d65d0d5047022f14d1b2da28603b6b3613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80c81deed29fde2236861dc4a1e4e9508535;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf0f2e59fcff974876fd86cfd7927f95d7aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5f62a450376e0a91451101c4ec497e9cfff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha775017ab21b3d398fec5da59924f2805272;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea6854a4b220eabaac53138b2b02c1d8ca2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8125f51b88ffddbc9c5c93db9271acc056af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf4cf1f5f43d0acbc6c01d749228e7cf291;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca011bacd6b8c6b599de250c9dbc83652218;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3425c4ca21426596904eb8bf30ccd431806;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8ff8abb2817c2327af93f16c69bf386522c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h400f30fec25204f263e5df688b82179bc772;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ac9f2711fb1470c92d6576f29d6477cb9c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7259c3772c689db2b72c56026e7b96a49212;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57284755a18ec07505486454da17e739f5fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc2fe5ca628fedb6276cae5a04e6bbd355fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26b15fdc91058cabf5ab6ea43deba43ad2f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43e425b6e05d88ad15febce04e0fa695b97d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e74d598ce9182cddd89ce62160e1728efca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57e86346308c5039cd3c9b8a6356a27863e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92966999d2d0ebea7ff3edf99bff1c47cd06;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8363ab19ffbdb5d38bd8ceff91d42e420f37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haae36881a60729f826ac3d4b72eeb6399e48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h328af7707cf7e6c568835e10b6f083b3c404;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde98b8ddd1a8127badd32b0b39dd313dc2d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37432fafca19d13c137ddcdc82de92323cfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4da5ee21b2bdbe927207d94ca70cb0e917b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac69901a5b0eee294a3508666c82056a2420;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1351d5d3e29b5b0998ebfa59eff5ed052cda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h946c80e6cecb1e7c6406dacf19cb40e2a7ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8c1af4fd35eb370424e1c20f278cac9489a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb60b788f1a7c2b8fe73c2e129b5849157b7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c83d8c03c25f1c923bc9741d9380c071cd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c4842044083fa076f2e140fe603b2e3796e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64e351f0355bc2dc2ff787591c5f7ecff3a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78346d8e6cc5241779b1591637af6b4813c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d4624a5a63a4ce750161e9716b6901ac219;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c23719c9b1b8286b5219bb4f2b9aca8f1e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h253cb5a553a5c9372e1de9fd2fadfa99ac46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6e831c9a92110252a8890b4fa675484771;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36b0d0f3220597cd09dfd73d17b55e187991;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1caeb325313bf47aee0f6d7c0a220ef85fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6944c6fc574e4b354bcd968bd6d53bdc5e79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a49e49cafa4fa4b631a9923b74b55279968;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h523a31ff572027a1ae49c74663ddd5b68303;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h856c2cc26c0cd76ee56e68f1dc312946e5e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2230eebd4809d4e3d6548f44368be80675e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2dc924be349fdb566a047d2f77ac959a2ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea02d1c5856fb720979ca8b3af29c36c80fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haac2ce438af32519610744c2872e3f0d638a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e25ddbb88c5b3a906d0a017731f1fa66f49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3011d507ffbc539428bbba182815152b1d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bdc98ea3c42817c3f6405a4f5379bf3105f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h664d5158a59d45b4610717e539c712300275;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde84c84684570e3dc42d8f148d1f9746850b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he591b509a06ac86c8f4115de4d893cce6e76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb293930c542460beeec37efb7e2e06c5df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e61c56fa15c5c4dc7b1fb8ee964132094a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25c809e14aa2615ab591727de42dbf93d352;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53d6c1bc40e937f3f85af12da14b1b3cb0c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89251dc33ef6538d27f71cb598b76e2591e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h940582ea91cff181504f6571c7ca0484a2a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h805a6ef17b6e5e2fd941e592b1888128e75b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd70ad2b1f3aaa5f2c27dfb7d4586024e8885;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69a1449e9c7a9175e99d9bcd5ea4854bf265;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3951b867d48123af10e7a0c6105d47cd3e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec4d9a6140b0108b3e0b019bd9c1ba93bf41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1127c2a4cea3b173dd927da2775dbb13e768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3b408111896a56b31bee99639cad26d6470;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f96f6ddbac2b05ef452259b4c7a9a5b2d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h306faac746f3410b3a174b3f05003a9f59f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1425757304c0361e7ef15581c78b1b727263;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd707648f2fd664babf6d9de127c7e51ca69e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h627819d66be370151a8386034cd146278a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec3eacdf1a6b8691346395430e283fa8eb7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fb079d540adaa169431f89185548289a4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f01dfa6c073191919b520460e6e9722a2e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb9dbff9bf54c95423ceaa347526840c4e39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h662d2be183483a45a8e4e0e9d9058c803ae2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3230044bad598e3e15c4465b119de55d2b3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72ede936feb896a166d84ef68ced75df6e66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h342e00970e6fe8bf1adfc2b6a361b36f1b91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd35b011d04e1695a5134dcaaf14fe4ef1a80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h804fe7b27b085e554898f3a6d3a1b8840c37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e2a4c7dff7885bdcba212382a2f24dca067;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h926fa00824a24207bed1c40f167926a731da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1849bf346a206215047a00216cbfd2e2a55d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha88af72e9f576287db5dad01522d15639d47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8439e1e480e5f34e2010d034efe73e32e9f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e8cca75704e633c86f1787c7e9e596f4acb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1b567794e69ea45e500f826237fc400a237;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc2f72509d53085da3c58cc055719724233e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b319cdef3df7a859af62f9cd6b1ffbc883d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cf634aad7383b3fe8554e7de5422e68e3a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9c599890a4b2e22785b492125e7ba0c20cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a5742422b1ea10e7122adb12cf390cfdf7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0456dbd1001e2b4e69a2f2f243d16627a3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59e51a4ba80e31f1ee27be8040b6c77f4c0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84cff1876f86a075b9e11e4eb4c37ac59b19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h409e1080cca87a2e9cde8c427a95c5ace389;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ee5ed66d3a19271079b043f29ead5ee0909;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5028458fb586b82bdd3d28fec4a033a8b30b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfceb635cdf9563ec4ca0a8dc148be02b8e35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7475a0fcee2a07c13d74c37d9a82cc27cec2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd081ec361cbfd9bc92092a1c301f84959e95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab8c36649687bff15affd6229c6f38b7bbac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1b25ef68846bc7f0010110d79f9a8555b11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7d47bfc0a7a4ce69d604609c3b7cc574d81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb9be8705f21c77bdff63b474315c6ba0a65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7e266e967cd20359bd1fecd7215de23d9c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h414ce663786367a516b68fa2ce46d6e4ab8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b3743f236a52e36c620996215822658acdc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdf0ac1a294ca8648c0cdfb52f758502d587;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c9e207154ef78f0164d2480456b1a5a463e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59d02614b828f84d4b40f6017f28608e40ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2f13ea3de0f1d84a92c9710bd255e7f14f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42c53f9a016b62bd51c1c06a9c246b8b95aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16a4dd0df3626394d2d9f991d6324fb8c025;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e990057bd95a815de19d5f60df876611b00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bda1d48c141c99f84af6fc619a51ff4c831;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe33ffb8ce4a59beb6584e97426da9ebacd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8316e962318300ead4ea7d843f5cc03b5698;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5190baa02b51523828726496b407f065f5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24f98265ab9db589f5826c0ee0c02997b1d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0ab3ae58415be6e6c68b6f5b2f96085d78f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5420f4b70f1a0b500632df80ed2a18969da6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he62e1fbfc42884f988599e2ffd99749b109f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e7cdeae3fb76f6bd5c24df86420e665a3fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8051901b3c2b09893bd28d005a04fbbae5a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1054c5cadd494abd3bc1bd9db007e65b29d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cf037ea35afe1e7fba64eebf34d50d638ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d035b574bc5af5e30d50f753557c3cee765;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95894fd8a43f482524792564358523ea9da7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e297955005bae95ad944a9cd350986d52a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99280ae07b3b4f405942ea193601d9cc9414;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67af21d04d224728cb2bb39a23bef1b00ea9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a961c5eb5983d259e83fd1eb3867fddd14f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4df473fbb816c318c04b411579d52bc75451;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe79ae7dd6a055d966aa4ad70848eb2b6132;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h625e0334fe08a0f3980cd27143378dc0b381;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3291340e5b28906a0f616461ac9baf72e3a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a3fd7195da3aef879ba054a2e2ac838d233;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5da081ecf3bf409a9f7c3a89fdcc7eaaf35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha07cf766ac201e21fa1ddd0ceea47d0f5c6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17c54d2034179856f72f82e77d61205192d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1d65d7758f90d53e2ca2e83e46fa9239ef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99121b802e898f1f63cca807c11be6c4b124;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4bb5416d1ea3a1eb4d1069a5d13c7c9a769;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4d4165cca6ca8251065e1f35068cb5229e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha18f94b5bac18aa5b6a2c28b1d01f73f8ac5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f37ce0549b25aa434c7ba14aba7607d2bb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc232f899301744ff5b47b8ab3276aade68f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c58ad61029cfe504bd08e6a5cd61a7779ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8fc8e6d9c6d1cb284ece78eaa52b1455e54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14a3002ef221ea64d11a0430fd8c32793dda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55b76f5346df9986be8f9c29450540aaf115;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b1fc2dcbc068f955de00be034ff63095fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b280c946a66e9186a1a4e00cb7fba0c303;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59f4c583f6ee965d514ecdb7a42843ae57d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29c85de91dc4ef3669a88414ee1f6e1d02ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf764a2db2f1dc6b988ab85c43f9b50ed946;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf797f5c32078da64c891cfdddc251cbd9c5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cef407d259594f7fca25f59a83378c59402;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7d9bc233e45fb73c8058d3ce8404dec85c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a311015656c454b6cce6955daecdd2cfe0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcbf20beb9cf47f48e66bae8500232fc028;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4eff4121c8bb338eb64c7c0f740aa8771766;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8212535984a000e972b1d8aa9dda26c558f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd7d082a6e054a683120362f309649f07965;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf30fff3ef756ef52e7c6e6cd10064b383bad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf87a0dda3262a4da605734375c1423ec1d41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3cba533c6f61dbde30f92b14b77ddd7b707;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fd0cdc9f08b4aa70f600dd316e4495fce41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e12b4ec19a8247286e9bd7f55f875391973;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d8838780ca546e96e1eaf9ed8b2c9ec7fb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23a0a2f126a6c9dd217cca13337e40725535;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48dd18b5f2f9b518137bb6b6cc231a47d6c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14020262e39c1e240753c1171257dfd728ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd1544fbf9a4de83b0ee6cc7f524b78d2f16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50b6ea8b27e67293b20da1eb40436f22447f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aedb0ed976911495fc1fefb83055699e1d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49d053fa5bc7bed95e643f6d536c125123ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha38767806279d1fb87ecc4bf8382ceb5380a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe082e2dc1b9cbe08f731e40020b71d982fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2253d657a301be04f294b282658322631792;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6427c1ddc00af9bce28ae1a68aa04c00066;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37c6e4e2620d10398ac2d448a58bad82967d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h300ab2b19855a3e4e08706aa5ba8283b6934;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habea6fb85c4d6dfc95e5a814fdd0943223b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc764ab860a9a750f119989fcfd583ddae39b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0399d09c3ed954aabe9a015c13338d9c90f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heaa187877f3d730f69c77f557ba3a91530fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fdb23524bc9798e6b87fedaed78def718e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba919ec3ad9350b20baf0f97d39f6eab7b04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39ceb0332ff94dcc7025bc95311076998e54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20fe849b40b69edce0768ef384dc56fdd6d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1785980942f1adb7d4e6b61f74819194b5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h710540e8026e4ea863f51c098bc12120f1a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h126b056ffa2cf9d95145a9037280bab5cebe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc2506a24b8d0c745da3e2eea16f6a69b858;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he21ac74557f57cd140295eeb4edba47ee1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce0478689e91fd0f995eb13184f7a494a116;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fec18418f0c51f8bf88bfe0c3f397aaf928;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1582f1f355b166f3176b50e13dda78b000e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d2adc8fb8689a7c6da4cdbcd7dca15b68eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdabb90cad1b2628ef9f5bcb97616c7ea6fd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb89310ebbbdf16ac1672fe7aafd18e771fbc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d6ecadd0429afd630e0d77c9c3f3def10dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cd22cb558ca537da1137d9bbaa7abf508b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff13fc1cc51a0cf28ab0a360f53d74be5fd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he40303370b516768cdcc9e28d093ff718da5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f2d36532a16f386c0f5ce4fcb13a46ac203;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65fbfc736790c85eba9ea8b193e900ab4f3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc336f1e7f714d7203b9b28729b47a773abb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbc2ca42dd0288e3a4534dee52a43b2a7c91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffae30c2088dcdacc1df48604db079c02f9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f518086fc5cc553946de7c1c5979651e788;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc64b2f7213b05164370215ea0a4e69da0cf9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f7c03c15132074e5ed8aa70d6a57b931e7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aecf7acd84e073036971e6832217b23a3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61e48a4b30f70e1a81d84200a8a8704a03b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f60b73b585dc6526baab65c4f24f770116a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55bacc8815923fbfa73fd48e1fd8d3c07f60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he78fc41b716406b5c4a2f3a8bc3847cd5619;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he15aa254e9a12151d7c047ff191fdce39c18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f022a1689ef7d4e2915c68fb7448a5fe255;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2a97fa2acd153f881d2a3321a5fe344d5ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13c68959e3dc0bd3e94f79eadea4e8f7603a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c55c4700b10817c3ebb44eaf24cb06d47a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he20f762c2f8672b413b495fc130423c2b76a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63cb1fe954d095a9bbda527ec0413a8a8e23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd618890a81bc7d4c9486faea455c04758675;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cd01e139eb1560fd9e9165e0c007a27da56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8bd0455e755b775b43fa81b643dd26c55a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ffa8dfa023ad0db351fe8432362dc9b5aac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7e64620fc7d66f3c99d2834ce341d6412ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ed1ebaaabae6cab08918e0b10d53ed9e5b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f5c6346753da651b2884e1684154a51c343;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha21df74d5fe907ce9e2a619a98bdcb4b935f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had1b151d36a61f5e6c4190a4d8f844a1895e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4673e4708faf173d39c54e3abb2fd1999a9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc35bebb8a42f9c6a61c9509e0a6090301134;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8c3912cf694863bda58cb9427494b8d6780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4684700b9ab9c1c6a2b30bf1a3b8d3e9fcb5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2cb54568e2bbf351173de42638694f5953f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9193499992677c32620bf006edfea07e6f87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67ae6e81551863c9cdd13692defa368f4a54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17b103cb29460a7e0fe6054981ba0b5c0f8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb212d2994f756efe407e882c9a9b5084011;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd36e6271c59b19c9b906ea3a9fb7018b13a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h882e66aaaef6e061e66855905aa2ebb49ae7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b62f9bf17ace3b03cea4f25fa3796bab768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88b7215e7daf8e9c8dfb3bb92a9107642b4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h342a401d409630921afe78a07b58843d3475;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81cbed16bd0ef9df17ed64aeccb4714b098d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha14077b4440eb243b8b50db5b3995678c736;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haba34b686b42fab83b44fcb1486047d290cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69edf38c6f84ab7170382f51ca4fa56f7681;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f90a508ae5935a0a7b9b12defa489bd6494;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2e476b78bbde0f7eab5d382474361e22b92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fb8d51ddc6579f39166e2da2177a8d5bf81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1259c7bcb24fb063b017511f4ccbbdfa845f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47087f87cd1f8686ba9eee4879fe36cdee2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h484a7035d4614f9a8e1f26b7ef31c5d2e7be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hade4ca8e27eeefdadd56e33f3836b8ebf397;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf23cc08c855e501dc6e898cc935e3362ffe3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dac50b02e75f65cff37a31d225d7cd246fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2fdaba67d5fc72cc7b2fb6bc359ca0deaf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h310f4ba38db8aeaf28451d8c6a8603bb4d0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0b9acd0de4a7b2aeb2f50dcb6b16ebe9c3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacbbf21caff8dd7736c061fd50b6eda9f3c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h559cbd1485ff2dc0b619191555a2c359a491;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f4d7bbdfe1541616b6a21ef77b689ed5a62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5abc77f54f4e5b3e4130b3826adebabdf514;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha034a8e60751814b848088185af3a3b83c7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb45b0877adf5c0c9ee1d3b6bd046682843c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bfeb7eaa9b6fd04a5db31a10b6d54e19755;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3b10e8c7e34eb314edae0047ac300b3149c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f0461a529f66a09d50bbd200ac438c3e1f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6a094dd374b74a8916670db6356cee90872;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fb5a5f58a74fd3b5e0838e9c11258134f37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81abce945727cf20f7106225cee98a78c1e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25f1e4e26f6616d9008411d114dd0843f936;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8150712d6036aebb167f92d993d0da757124;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e352b9cf68440a1f4c98651df22638002f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7932c94089a07d1ec7197ac83b1ffa83041d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22b891b32ef7fa2cc3e9adb5959e2a79a13e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fdf9301d1adfad81fb265177ac6d3bccea8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h598121bf30da82b84e856f4d699923489078;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h333994dbd803d29353bb60d5969fbf1497e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a0a63eed689874847ee260ab0658d20791;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h748fb049ad1c50d7219f00f3c73fa6d11f3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a915d23ace8672ebb53730e6148b0bfd77e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed1f480ab562591a6d812acd669785c5725e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ed678f0015cf76a962bba4e526d9bb38c5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he088a6998b0dc89b6fc1436498d654548464;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h200b411a538ce1928c14d24fc7ae159c6422;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2c091fed50532e6b727087625520353f841;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d7326813b15fdb3ea3c1593290ad0d3e066;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb28480ea6007b3e1432e18ef2ed6190a374;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dd8bf4020d8909f698d87c8c051974362e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4b414a7be5022b33f092b3d5e00feb2a03c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb86530f22b7baa3da2e36e0f2651263cc6b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e9869685a1ef5f0e28bf0a4325bacf8658b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b830e82e5fe08252b9d00bfc19d6b946028;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4940a18b9b90af31ff97fc6a916f734b7207;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h801e35425a35e15d24f64d5427a728b2d312;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a60012f3f8166c5a6101d51a078a5128188;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4de907ec3f37441e02c36d4421f9c3536;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58f16edf984656611ce61fa2514f73eedb03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfdc4a42395f0ec15430ef63c199b4b32a11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h846a6dd68b0be4a7e50e8275803cd9711735;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1deb22b854f0d082cd39534588b96298ee48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15e8c51f9530f09003f195f0e9a4f2880957;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8422090a868ed8f5f7a54bf21027de95e5b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a3b4ebe342f5a57923e2227241523b18d4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27d02726b6748579a13a469b9ff5845d3f2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef2fd0b5d42ab92692b01b552cc3fde034a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ccb174299b289d99345f461efc8f79e86ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2853f09a405601a497fb0f00fea7b2dbe27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ec7a0d1e70fc4a9236125f8b76374c0e3e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2579d2a6b09571a30fd068b3e7dcca6bff3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha925df1f571b3cd9a467033ea1185c9ef85e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ff2d2f159e8b553fb2bb60ad3dea02eaa94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7566d0dbc39722700baa9ff63870611368a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c7737fc47c3699f97ae42c18bd2b4aef855;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb17199e931c348422a75a044a4b5561036d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha80a5e5770cad96212ad632c493a269dca7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha82a180622073224b9835f25ae1ec12a42cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc21319672f72116376128dd633a9c3973a12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf36a58fe7d37d528e3c29901bc93ad7d265;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4957d0c06e565225ad632f39338e413783e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2182202870722e1ad30f8c56ea04adc7547b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b58f62dfdacf803e4d84883768c304c72b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3d2e05944220a91c6c79634b10326863a0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h723dbfe3e23df664767ba0d93d87a3fa393a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8f64e91dd9a887270bc29061bac5b7b102f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45b810f10d20c64a4d84166e93cbd260fc73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab83fa054aa078d29683cd221c8c630d020;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4f06497f0ad2a28ee4001e1462d35936ea7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he39ca22af9e7df66bbc31e91664ad1226e4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b9573c00ba62bb585e761e81ede49737079;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c6731188f7329af3f1b943097cf21f35a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h581696cfdfecb29712f39e21fc66b2734a47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h388ed1afe810b56f953b076aa0fd0ac50b20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb24b3c882179f8d77089df5f91c1caafffdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32bd4d10dbda615716a3d6b9c183ceea189f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea11169509614e30d868da60030e4e50e4c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd38282f956f27ed2d47ca971084721ca7a78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h272a92f13c92bbf7c66cef03424407b779b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1f6a16e84f12418150b3c7600279aea43a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f7a4e6660b495dee1a3f005d49aae60e193;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f36cdb0b683b8a31859ea428e9d8592ceb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h707cafda50b259142cd043f234e08f2a8826;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9836e7f3672f3a53340e8cf28ef5f043bd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5cf4e23d16eaef4a57ddf54c720ab407db6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha71030e158c255638031e9dcdfa63c607863;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e6c3dd2fe9632e5ca3bd2b2f9393e606dce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20338ae7833196efd3fae19a13780e692788;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e0d892c6c48a13c8a0a746915c5d1dbbf76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46e0353e250055735e21d0d604355fdbc9a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36a620d29ccc09f8e8c62792030c0fdf471b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e6d3a021a51b7a05deb281b031b3d0e3e9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43092c5db32ccdfa467a04b47d9848426d22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1beb51ff57e69aa90826f47f867a66680ec9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h951fa8a3316bec3cde1328c4938ebf78104e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3bf7f8854cd0915edd609a05ac39288a016;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf85d0a576f9a3ab34ac305f126d8cc41d138;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd272b41940382bff1f4779cc033ca3644613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24b2602ec7f1eb43d217688d57da24eb265;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h796a517863c99dd55df6aa381ecfb85bff45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f71683a78d97c57c3f3f4c6fad121139e0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habf80de7a5e43e45051dbbc320467ce579c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fa021f22632df2a0959aa0ff43e5d05aa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d5414af04b7aae2bef03e9fa2a098f43164;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha52325d6944201cbe356006db3881c98f68b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f9be5ee873053339378032105116cdcf2d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1720bb0877c23df775e13207084fd829b2b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4aa742d02ffc6137e50a50b14c301833b58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76884fd5a5e9b155e69da43dc9dd6715edec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaf06f00869612afa8bad2505019fe004a58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32dc197c3eb67896f7d66ac7978eb03da03b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e552cea1a26018fe07e90e7075c1f9b654e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47cb9e01c27f94de6f4cf6eaa7aa1ce20f7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffd07d6fe7f3df384c017fef11dad6512e5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f62d4f7120fa07daa34a37579da8f21402f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e7110ea188a3797aa30baf24b72efc5f4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd27106968ebd5daa023d47ac2fb5e83a89ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf867ad3fb1eff8f2b1485dba4001a18c5856;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1119a3a261daf0794ce20fe4c83dd76ce4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59adc7047cd9d5c32ba729af9dd278c1c8af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc4a8e0e55faa2406c734fc68b3e554d2396;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d71277eaf2440fd65992b8319cf33ed1e8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3910922bdaa71774096e89476b2d68d6e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7893dab88df048442f2d1f84f7782a24d75a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53b4dd52117a1c54b0af45d68113eafb57b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8db9b297058edf67078aaedb9db63135dfed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17c514e2b3368bbc008471d49bb838a31f4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h279883796c5465c62fa74f84411d98705daa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c39e3978b77c6977d4c4d242ebfc0ba217f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb0e2d764de4b113850e75374ac947e55ad8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h452fcf279c7076092f64c5175d5c9b58918b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea9ea1b8ee84d196c48cb0099ef77647a9ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf950e928c8cab6348226bba2cca29f042591;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h311913441a4d87d38a2c0b2e04d46a084b62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb865ea25b3530a68a8648182495b54921726;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb04c8bcc3312ba163bc2a545ba095ec52aa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab8e55304296febb187d8533a4276327955e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h160d07a6faa7753d87958f84249549f2b39b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h196a667e16976b99206b67d13791adae3060;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he01c088dc2a1c827b568a0169f03ede2792d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf572e5b676b2f72a606e686d516b0abc3be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb86ae8e3dcec2137ce4731ae4d1077ec652b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb05c64772afbbb93717b722f69415c5d57e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h885be56fe94a249d8ae631717fd01a5b656c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb7f9ef77eb94046d298611166c1b79e0526;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33d1f4c41a2a16bca23d2c390b662aa1aa24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c9abf8e4a24fbfc0afa41819075bbd11d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba0040a753a2281e2fae2745b88464803558;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e100b3346ac6a34dfea48b16da97e98aa1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21947b8568709c021304bd4215af316985e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf665b800e4376774f8525bd9fc966ed7637;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fa71a9f37973a91aad51040315646f82248;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2de2387ab88554f12cbb08e54785221a648f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13ec5271cb7c42bcf526bf1a13ce370c3346;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc005accb55043263ef7bb9ed73078f43ac9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5f094529aac673cff9b2fff713d6d4063a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h819cb05dbd4401dfb5d1f4e23e549abf2dcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb81424e69e597df48adcd677769ddd36b3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4288a3daabfefd59bcfc3e50f336802388d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8057808b09692951d0b4a3b15c2aa00e9657;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88e7321c9c139a1c41f513a115d9db8f4142;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h394d9311cc8f7cb9fb74275b72b3eb4f3b07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbe81c032c29dd154c6766a1856fd2e307f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf049c352f386470bffabd97183acbfa19a18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d33bdef186951368f61613ff6a93baec429;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc4cfe5906cc7ee44db7234be4c1722472ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha116c1c80ee5c84b1dd3ad074026235c2680;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacbe71a634552613f833dc486cbbdcad5e92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5001bf8bf54e30bf13c807157962326710c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h278a7b44c92b46d0da176b525ff0451d2f48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdee6fc0be17d93a549fc9cc3434a2da028fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h769bb558ba0a3b495bf74098319218dd9d13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6dcd479879dea4f1c9ab2b1cb9fd88554f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h866cbd303fc6edf2fe5c3ba5139fdd60c393;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h927b12ae6f194df16f232743f1b055471f4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd1e9b4cd6c8640e60692beb8ce759f6fba6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h558c8bf7234fb824683dc720782abbcae5fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91e2a0c55ec69b8376bf0ee0268c09648088;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b1acf741af72c3c1cca3d54845c70ded48b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52d9c4008d7b45abdbfbe79447223d2eac61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ca06be31c73da0f182f79d11c3be3904030;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2807a47883c02a4e9ac9f55804769f207eae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56b97429a78f082a0761a7ddd44c2be45846;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha18ec09546996a15d2353ae6459e52aa2ecc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f448258bc63300b6dbbdf44ba9176c7f693;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc56ea186523545962cb63a34dccc2ea50f43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65a80b05a50911fe926406d46669a9866808;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94d32989540815ee30c7afca04498a64fa73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4a81a7f24504060154440253eb56001d6ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ff1f3fdf01d2abf03511723362fbf39a74a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34edf40df34a230f9d9071c6d94ab7eea61c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc2efda9fa48ff8e0ca28ca9bd2fde4d57cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8349e1ee46921fa2e2a5d4b6da1a87a324a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e2ea278755e48d1b8a182594109a97e8dc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac61c325a33502c6373364f3cc0703c44950;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h976e4fb5a99d7bd86bcc14423c388a494972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6caac61f0977a1d7bef82733470dedf04f64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf504366595fdde6a7d897b6a7ebde810a1ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba38531d4506473d815bea774f784a262ce8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h603ac47134dcd2146894bfbd852904c801fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h769e18e47e3e47a2267bd256d7c3c90b629c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf15a737ea0424b03027e19efdcaedf696da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc83abddab157f6f22aa26bfaa2f5089e14e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h142cd472185304dda1b90300d7f06558dbaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99d234d733cb778ee549a737795fdfea8331;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h645d2b9bcc3352e9beeac2d0aa49d1612e94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cfae943ed3df9a848f0f5f6caec485cacbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h249c54d085ca5492d56901daa312aa0fd99d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha67fb940df8ed87126e6273e318981d920ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c4c2a4fed054fe96deaa3c0928a54bfa39c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96ad90068644e05cc84607e01a9e081528a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d85954d1b2f41733de839ba2958e35f2993;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h189eca5f9c8c9e0f3ea93abc814d5bc9aaa0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he86a455b26a394dafec44bb512dc5468b727;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b307d17050b9576e0aeba33e60ae99a4f24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6da8505c49fd7716f5a99ad573819caab3f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h759e9d8ce353e9f6ec4596b25bf893ffdc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3117be01590bd52859beceedb9d297fc328a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h696d8013c1559c1b324154857ac4288fecaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eac91e803a4eb8cd7de4fb8b54b443d47d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd31893886919b29322389cd961d8b535fd3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f0fdfc5189d31a9121fb1fe6a2d97abeedd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81df9468187bc648f7e89cf85fc989512820;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5a8abb33d25e9d714178ac3e7e107d303ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f3c64ec664da885d2b0c6a69c16c66b1c23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h463607f0fbee99378208aa3df12562da7b5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48a167a5384a7bdc890c9b3ff459dc85d578;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6ab0724e46f278119400f484167cd49be68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b2bb0f89c4d67d6bb2c6d79045600fefbba;
        #1
        $finish();
    end
endmodule
