module testbench();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1975c6a3bae97759d5bf2a4f9df5d4d54f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd438a01ddc35eeb86729f9365def64ce43df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h433027269b173bd056ee4ed5f8086f831306;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dec4af9eeaa2b30b6814019a35d13242e90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf158ba17fc123d5da3b96e2bbdc52ba47c49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h303896d70f9cfb86a2070fa329ac93555772;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99920845e8a19ad44b2838adb4bea1110971;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a713ccb14969d78a0f6fe8175688310584f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a7260ff2432c2f068cda8fbf2a1e593116;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had866c73cf3f501b423175ccfe6d6eecbedf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha107d5b5f7729ead21aa1dcbadc15c727197;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff8c24d6a8efebdcda0ab83dfccb63ba4c7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa83a8bdfc4ceab007f75e972576f9a97e64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h519ab9b52ad3ccf369b679072b903b2aadcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc233ce4a9df390fe8586dc72577f7b73db7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf25f2706f741645d842ebe481e6bdc6fde96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6895541901c4b98d303f647b470af5ff7e15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ea6029669c351593900a5c989e01c3f2839;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab9c75ac38384b11a02773c094d85c66625;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18925764746cda8e9c0fd49ada9bf49e0698;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84b503c348ce39c6790c37debb19c007e7aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c42e4ec6aca92e511c18784fda18a6bc2f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h135ea02c061673cfdbc4c6fea327dc78198a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73ed2d434d37a55141736b1696566585c187;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90f30808b7bc319ff3439197dfbf27b63213;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b849a3e30751c6e3f246a6ade71dfdd176f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb571c8eafb50baf773104194ff3861ab1671;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha699a87a54226b594e14deaa46237edd06da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha49e8b45dbc7b8cf525b8cd3389426d2dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he40c4ab9e2f39c91cda6b418fd69ffc00faf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b3f6ba3ed01d790761a0004e0a36947bae9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc1e81426df946a81b1502a1ef29016180d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3b8c347bc9525f97faf90198258ce2860ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30454294118da5569e71e84718599124d9ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7c2edee6436a4bf106b8804d089fd834024;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf5c6f8e3ec35c1ca9020b5699e2016cffbb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76211e54e1d320133e7742521892c50489c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2791313fd0678f4097d6710688e340e9735;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha430ff3f075f953e8a28bbc7ed3215cc83b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52d31d6fd7c51309396a8c88d50d26b3d4ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79f6375308b6180759b53d0a6d613f8e1ec6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0d8430e04aff91dc843ee617c4c0b7e3b40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2de385fdb22e4c95d356665b21d4d949c11c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9c9702ef7e32445c86673598a768461f9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb034e892a6e3d408d8eadf5bdc808c510b79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc45d6fdb37ef4fe92ca6c4d5f17e27387cfd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52595b58f28550da5a4d44b2ea7d64673c5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59d2a7833563de552881b4a3cfadd0e4eff7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ae9f7e8e23a9d568673c93f3f84bf6e7fed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h282781d883e4278a1ff55d09a4fc4ed6d00b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd29da3dc3bc239f5b4a46829ec85013155b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ae8a67beecaf40dcb512b4faf3d85b73556;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2ccc5e1f33e2084915922e5e20dc4eccb85;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h735af8d9c9fa7e64c05f0d0707a94ee80b71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7226a79f4f3ddef051363773cb53f1730c69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb47a4e99efea0432dbb54385bc7ac53fbff4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1689d822e780d43b3cb8ea1214ec709b3644;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ea9820c41ab8a898d1371a94e7ec0347810;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9765be6e4259bfd9ac2f1e70ebeb2074d90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7d7d093f3481c612826a81b6f8c9da24fce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3faa1dace0d6f517ed8c74a249eb402bf217;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hded38013bfaffb21c6aebf96147f5dc1aecb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a26e2d1a237982b3f9db62ac85042a36524;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbfbe2a4009f88f24298b3423f25ff70f5c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd97f12e46afb8a20c41a38d9b0a313a645c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25d08e69a62b1bc974d9f8320ce4b7bf8690;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6c13d3d35980f08bc09272854d35843adcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3df11dfce4df747481b61d0cf9fb1d4c73e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17bd13178e184b19feb7b65996c57f31ec6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec6fc925bf22ed09fbb0fdce2ad3307d3425;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8006ba8222b3d20aa9047f0874e1be02f80b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a7fc1c63b385427665ce32eda6a05ca52e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdece2f3b0608d323c1857ad5e83b1bfa03d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d63d99843acf2e47be6b91fab4ee2162c48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h870c51489220f2712bba994b6866051b041d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74e3700082375d32f26529b0bf59a5d0859d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9907ae30dae5a64efe2ce5934debf403736;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d3b3354a15d2d3f3505edb8e33c1a2a662e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f4d083ad8a0770a35eb7f3fd9afaaee68df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83933083a6b47ff5b224cb5f1b5621231d70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc33382aa22be9c7cc16872f9e06e0c725dc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d9466e44fbf352301a4f00c96e8dbc323e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe9976b63101a58cbe0caa5f59463a7dd7ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9694996f7ce9a19a3d3ba597f8a0ea4fe497;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65bf68ec6ebc7e827717fdee27447ed93a71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43805b26c94dd17f9f4ed386935d86d1de0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h878e0ea6e589abd83128d4ae5af965de407b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h644282cdcdf6ede0dec6be17ae96587a9d9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5945dc4d56f816557043ef42e7e31842f46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4476fa347716c55e8e43722fd887ac94515;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde882d0e3854c8a400726113fb900dcd5975;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d9aa865f7ecfc71b806b960adc5cae4c74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58767cd457f42d227331266ddb4cdd0ba9db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h188ae1e3b59b5fadb83ba91966d3236f9293;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1e9e19b328d0c4b2788bf75756e9e75bf51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7eb1c121d9ef6561897a80cf34a64690aec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h479ae35c449f011a0a032b60441f62dc89b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45a17ce002c0117276f8aa4b71508e1fe410;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a028c98950504be0fa52d824afbc825b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27990346d55453fd0ecd17ce49b6f410a4e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59c7e8efd99fde96f99a3308c355e7556663;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4301d15e16478423199a3472d4dd9afc26d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58b98eed0c740af3bc6b7e53321cb06eaad4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99e8854d728c0a4b33faf6dcec2808f5795d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd895d048e503e9ce808041ff89f37196bd38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4ede0526fc5be46a3d90c6b80bef3c982ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d873eb85e092fbd7d5b2b6bf91ea8d8185a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1464f453a21478cdb8eda2fef180d5153c76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h491f6706f95a8d123ae5bbae90b9c1731a26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6299b4913a1a845afeb49707b81e052acea8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6308e5c65b62f07d89a1bac20421e5224196;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1532d774f9780c24a29663bd30726985cc7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h479291e2191e292dea0b8b29848120af8ae1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha33dd7b138d89c07ed0d1faf86dc622a11be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h250efc918f8dc2424e5a9e4f3e489d912dcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8908bf06f00a5d7fdab3b7d45aa1f0b906dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10cdf4d8c74bffe4d13414eb37dd994f592f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef5d05b74da2000e20abb940aa5b0015c599;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ea495820eee4e10bb643d861d310d3c6007;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haba0b8755bb2002db7fc537310ecb1429ef8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h990352a73ae19f785ade24913e8528fc75dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7325aa2084e85a6553ca64fdc88b98c4b79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h693a0365d2d802c0a022120fecb619e8c7e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h187ebeedec17bbd1d727e7153d863da7cfd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf50a36092ea79b3f4b1e85a8d765be20a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ba8f944c3f5858ebc94ca3b5f72c5ac5b09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf4c2082a9cbe92d17d6e345181547a6f443;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h365464dbe4178de1769aa31d6a2a0db239d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h156feceb8ed8d7fbf218be0d1037ad0939f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc98ae28e00413c604fcfdaf3371db2d0ef83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88052a6370d2520f850a8dc17a989cb47904;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habe644d9ec3fa51ae145dcab0aa7386eefa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69bb956014eff4b6aabbae12d6d0d8faa613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ff1b3f5c5508153762406bffef572f928c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd79b3eb4d77f4048605501463d6feca76dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h664f101e2039254b7e0b442993eb548cd7d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8724860f8e53666cbc8825b1071414feaef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40dbf83ecaaf76c8bb1f05b8dd3f82d22191;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf306c840fa9811171fc1451533ecb8ebe1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31974e9e3815c97c628d57913ac1e79ea559;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3533c72af4c4149c27c2dccf9c63ef5a0afb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b2df717f5878eb1f5fb3bb2114757a2d958;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7734279b0fd1827f0a30af028048df484ee0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2791742ece1b99b297b51fe2e7dd8687569b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde9a927df4d276bd8d8a73aa1fd90cce350e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h505b36fd0b29e73f586d024403264af92725;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63199f67f050e780ccecbe6a0dfc06b43a19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e5dc3de8d0c209c365f5717790f31337ab3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8685af5fef37f730d54949fa8ac795c22fcb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11271727a2fcb0da54fa03b193498e8c6d7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3050e26a0889160aa60e3e4ea0bf3e1f9b1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1889fe53dc85e630c3e93ce62e51edac890;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5f4db5b9367f77b6f4188c35f98204b652a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb46c9803fbe6b955cfa198036decdda2fe48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h994475d906f20fc0f0a6b827d265a0cffda0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6851c1ac39a05ec1f1ea42bd59a65a996e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5f7c77bfc17e96d42e99fa1e74be4b1a4c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9268927b0fc4e368a38520bd3a4d6d7a6bf3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f4ae64df97547953d28bc0bc0c7c93727cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a4306486078964aa74d5f705143260a17d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28aba72ae04ccafa5ee39089ac2d8445cd8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9d1cc860a1a2e8ca2e273e4c223ffb2e84f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h376f7bc12a2444a74d3be4d31d767f36a9c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc29f09f6977e1c98ef2b5327fa06a26f63f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc483ff0b2f40eda374ffeb2985827dcd3616;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72aba882d4f0247d2c82a1bfa982a35d0e10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94fa20ddcddd1ca55acfa58e877ba4da6584;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc4fce6f7a5de67f64f728a865a3c46728d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9efd8e5127cba14a0e2db12939d3b8fa4d1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdced90a669d78f3eb42cd50a9842229eb96e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6e70e8212b6293e3d1c14e6ec247283a4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37e78e72255678b153b60edc082fc14fdcab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e7febccd4055fe799638cb6baf7d8c9019b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c06bda697dbcf1ec3ec1a0ef29929f46a90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a2ea894bb9f86ad928a77d6f6e9e7d28ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5525ca7a19d1a34342044c4f2141b9ceef60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfdf3bfc2f0342c5c143e04e0a4726e993d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h690b4093094ffb3922e0131c792c5a181284;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf444ab278bce982f1f4daabd34053b09dd2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h343cfd68e497f781dcb35cc9c00d3361ad61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92003c3eaf55e36e83f816410aab74a17f4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff97df63cad59176a3b277e70751e2df1bd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85b9fbb8f6531e3c5a0a87ace465389c2890;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8d7ad8e8e9d541f08debec2cf80190ae7c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc2e446000deb42ade3cee632a12e7bd361b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf4b6968262ed778dd3dff69a9527fa82016;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb88570477f35afb88dbaab89341f63714a17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e586980507d89cb578df51853cfe5d8ae1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b6b1b73486c9c50e8d656e25194e89bd06e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h645f93c8b41ffdec6b2efc588839456aaa40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a2fd38a80279e7d4b440e3000ef844e376b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h306b6a31699a719355b67ba62330c80b7d5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb04c23f8d68ba7293291d06325db3143bb12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe72d585622f12bb8d241d720d2d8b27a0c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf212e5f5a1ae70209fe1640b34ed8d7b5e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafd0aae6a5f8d3d0c37d7b8a0156607554e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h983a8e73afac7f84ef82efb86846621afb55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d641fd4b468281be02e898f83492b438ec0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff30de97a67d7cd25de522c4fddf42b9cb4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h393e96c0836fceb57a8087f04c8298caf65d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89284eda323b6b019b5ea1ac8d933d9da651;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had65f622cc00d5f625ef01982b496e85c42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd6536bcbde8d1ad90604e90137aae65d329;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9f801a5798d784a8b15bda53ed019193e6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f4c56621f1709bd65869376cddbcae32849;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b7870913bf05ccef0cd2e8a6f3dcafb2b02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he17ad6695148db39a23c1b00d78582900579;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75e5d068368298fa6d982f05c2682902ebdf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb82dbd12155536d96edbad4a666a7b6366d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31e5c9c9b2c11ee11c31a766f55e8c0d31f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7eadefc969d6e453e15e585a93829ee5c3df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c8b1f5511481de6e04446b33d4b61231229;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65f82cb1d923537f90f689cae76598b285b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21c5d503df147033c46ed61f0ac618a708ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5e118183a185dd45d7bab2780ab0dd79e5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28d4c3c239b365d276ef193c69791bb95b45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf850e03e1456437b46bdffdc80dae38f5ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34a8ae1cc9609766da4b976658b104f8045;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed771b366e9e70a5615706ca95aa20d1b25c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a17ab6bf711404b032db930ebcb4afa83b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfa016438654d7169397838c76b6038cee9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha72981988a33424658789bf04c16c90dbd10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc10182bef864a06229ae22fd1f70272b4502;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7950b33b77829b05d6f169b97255d282ee3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2506368b3b59c4e809e0669d5b90573c88f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5eedca3f60acaff15aa37974d189abd5264;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d0c03055493253fac5a67f16bd32b521f82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b54b813efcef4327497948975fd74d3116e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h595469118055e74ae0dde10b32e49a926fb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0821446dbd84a62dc4b909d5811e375235b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcffa8c067bc6d9c1805e17f63fc04ac480d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e850acac3bf0c96f26fe92ec8da3e0fff51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37bb1dec1519e1229a3a58ffe70ec963137d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d4374cc3be4f2a04ca0d953c131f72d8c48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h607089cf3f3d71a10a21029dacd6d493b6ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he63ee4b2bf71c992ce273ad2fb32f703c10d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h231b5ec749a0b6a84f2100312c50291497a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88b8595e1d62a1232045ac0b4f8cdd744578;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha78fdedc2752f87c6878d6f8ed67e6456873;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27914232aeae416eacb2d483f679fb831c52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9700d084f060b8a2d1299c5d60024aa65e13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ced4b1bc3d90da3816d9f39d7eff06bb442;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aed4705fbe8f6c69653a89800726e7cc5a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea0d51ddb104bf89887e148b780c569af33a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa57175d649014ac2663eb961d0fdc7082fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha71c1dcff6cfd1b83e3db63ce85b10b39878;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae748d7fa92c366442490142e594e46d9d7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64e802888bdc50e49a1de3fac94eb7ccd25c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f362abc75607d7beebd1a4459ccb38d02af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a79ad8af605fd3c37059626328cef850cce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed7caf9ab181011983a8b1bcde9aaf2fdb53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f759c796b1ec7f8897ff10699ca696f0f52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7b0816ca87cd75293acded1e5bc8e3aef16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb833f969a6a7ad36829bf74e4373ea4853ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87dfb9656eb6e22f577c1c85a3f9c15939a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf9716fa7b70a4a0713b52e2db72d5fe3f98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87d6c2e882485d75ac7dde875a1e4c5d2bdf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a09d59942a931bf471283126fde4afad917;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3194cf06c9d349e4e9cfe87af3dc09ec0a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55d1d568359e6d8aa69dfa25fc82412e3ef8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fcac145d3a4ed156125c2b7ba495a8a2cd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb15a1b22efb932c8efd24aba1ddd19f1960e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3be0d998e4c69625aa1bafa7d392157598e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf689d49a814caa66f8e51cbf04417ca30bad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dd976e2398474106399ff95cf488b817a99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40f91ba0f614d7c4801c6adc3f657eedf8af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h595bb5e23f96389fcf1a0487c82bc7189652;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb797e758c3eeba12e6aec259abee959199c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25f5336042f4f6462dbb76f052676062197a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h321084a8da04bb7980500459db023a415708;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc63058606b19147962bdf79730d74c06cb39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb278e5ba3a64e36694d6d99815ae8a872d3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h361a1f81242c35bde03f7692fede548d2210;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c09fdedadfdd8077b4af52ec7aa81f5e060;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d900d1feb8cec5c82a77d0ba30f558a69c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bfadc134b468f2a9a1ed09cf1025522f23d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc24120e14cf3f3cc2d25d31a3029886cd15a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25fd8671abf26f30b0baae88072ba89d8e97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bab49e8a5ffc74f364ae5d95286623e0b1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha62bc408b5279e07731b595882d349ef8506;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea7a8849f15ba256d622e3734e3a58edf806;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h333bff144382774bca3f83c8bd06d69d8128;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74d78f9103a54b52b8d6a7037a5826266258;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10e29d49a2438c505577a744d50799af3354;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c413fcd7a0b7c8cb1b007b89861e978c57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdebe7c108ec715b0a0524e79fc029a5eda4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e48264cf280f5d60f047412e224f6ea3c94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25d57a23bac782ee4167f3125ca382ba6867;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb21375ad49e124003420e25ebce9c9301e56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b24451e7b52080db77b75191396d7dec9dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd19f8c881f5095f230826ce4391c3584a6f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f929c7945b46d0c1b46925ac06d1eb21f23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf49db026fbd364036d9bb4ea74ad5325a348;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43e78782624e580089fc70da50fd7bfc4a21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae0396915c9a15c23008933e3c5d98c1ed33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafa454c51466f543ea84631f7984f99e8189;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h351f5f5721e79f87f7c854adda87763e79ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e7a93b912102621d1da92a20a57bb113d04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf71f9a19ad24e95803692bb19827f50c3ee8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha83753df4fca849a23d13aefaabd244df3df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24fd238966ad14776edae1d052027fd4d7fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h895352a49533f5ed192b6ef8b70bad1b385;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18d00a0bfbe3fbb2b411883d0741c7988144;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ee734ca0cedbfa47eb2ea5d334078f2fabf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c900788d2755ecee236c36a8e5ab4732c19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbecf9fd4b92197b58d671f1af9112ba95ec7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0c6fa41fd769d0aa908e682f6e42b61586c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d3c60af08ae8ab3e0dbe3104d3617902d70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71deadd4ee02eb1aeeb0f5a9c58168d07f86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2de9d6106e17bab8608c02235f6b76d105;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf73d22e581004fe9f038ea2dd089628ec34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bbc143f5873047cdbe8f4c5fc9b245efb53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7de3dfa937abf5315e7f836c6921996b6ea3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcc7ae4560c9223abaa6248855145fa1824e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5af202ebb2d3a0722fe987579f7b57166f3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74557d65dcb22a5d308d88bd7fb20ff41965;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76984dd5167be836ab8034ebcffff8eddf0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h309730f5aa32e2dea4815d5f40f72958259c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cb132ca98361c882f18c43b474ac3be3bad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha55287fd6ca49192033da7b27509b2d574e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59e6155eaaf872d72af32f8e599abdba114b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a1ab0b61e610b43d20b016765feb943b1cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81f3862dce6cf948173640f9c7c67043d177;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc727e4a39f6385667b33a6e1840dc4cdc2c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b41d6a868719e91c96f787dfd3472e9a45a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69d6213411317abae8bc77ccff273cea62b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9545d2ad578519f7cf229093ea2ff079443;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13b1afac36c8774c3176c993c63e78316e99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha60580b9dca57fc647075d067d9bd11aa632;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dbc0d21b7dc8836ce354c0b68c90b5bc3b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f9e879fc92fbaa26fa4e1195e3064050299;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1db9e88c1d6042f0bd33d74677defbfdea08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19d69a8da8749aa394de79e6091a1e6e81be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58a49e53b8c3e4e7edcacd928b51a34f9c18;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93dea5866fa04ab4bfb5a7ec4cc1613c6825;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a7e0b5c1acdae209cb559ca7f9f09fdf945;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a5340df5d9be3dbcef735a084adb93e5c92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6561348e8f51e6a18428e71b33a6c506ae03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26a97aab05e1ed2cb4129864f4807ea0acf2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68ad63bc63c999d652edff39758dd1dbc9b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had2991a7ab282465f7f0009d7cb62739189c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30dd3fac4d3c4f74eb9ed3f00cc1990c8a79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbec55e6ea3ba84b912dd96c7cb04770a08f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96185f951c93a23d9a851b4c4b209ffab9e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e4ef623d9aa3cf2dc4334c9006cf3107e30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfac83505ab11b78a89d45ebc615014a832ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2c36d29e76af054d2afc295554a7c71f34b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd72fde70469c5c17122fcfb92b302242c40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cfdaa31fc91b5648e220488f5a4596c25b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2a2fa9d4b92c5fa4663c3a5a7c5586b6b71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22346dc7ed491f451ddcdd705f47390192e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e2b07d9b3bb5d310d1bf1fab5afdc0a3588;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b00fa1e2cb3f2002aa8a79f75e67633aff7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h417053243431b590b8b47d646a13be740975;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3ecccec25ce36be31b9d61d1193d38b342;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c769fee252a07d6876f93090dbb9e046e3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fab2d1acf6250a849cc410464351cd86457;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe47968839242422f88d6bf640ca472f6a4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h811c490379ac946b43b0ca564ae9ad32aee3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf372f0c5d105bc228dc9e815b3f85cc5d85e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14275478dc920881666054576552e7d63a93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c1c7fa21f0de26823219285b07de90311da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf04600d0994f92a258f6d60f36947f4b6705;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79fce3f789dbaeae53f974b919b9e9b9501c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had7e4d13e921d423a9f15a30e5dbaa44d6bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fb2a8b08ae07a41f7dcaa30614a69f097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74342fbd46d005617995f83f3c88cc11c8ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd093bc310c48aae221a205cade26fc5735fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fce768a4ef779bf51335eea413c7333bb4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9d80d9c00b92aa70e55cf39705a7a6b029c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dc70e54cc3fd73dad5c89e5703028ec9fd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h241e7f950fa94071c39af31bd770ee3bcb24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h751b3534a5b417da087355c6d61e8921f7b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b3b87e5a9274634611d2f618f6925249ecb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d3774510a236b80a27446dfc81087bb9dae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5d28ec935bcd5fbcacdcdccc11e59ce7d7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbadd7540b15e4b38134bae9c11ea27d2c447;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb80328a7e55fe6461b2ed3a2f1149f7672da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8493832752f87f2e3eb7a0201c46cc96dca0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbffdf11376ed2a66eafad564246b2b720b36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d2b4020a9831e8a68e7a53ee2c2a0ed9c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f6a26c4c2fbd4693acfa6f5676e3871f4b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2ffa125ea78ef044ac5961e5bc9007a15c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc912a6ee7b2296cbe05c788ad7964beb1fc4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb6ef1198e4254523e537c6eb115ec10c3f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3882e8d2dc6062f363ffcdda3cee96edf48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee717b9ca2c624f3cd3c14ff144c80f85b81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cfd0b3c077f152e58b81ef56fd3387f99e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb90686a041f97c4dda654dec310c135f7c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e15e106f7f75eab9ab9752df276d85eb48e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1e700c87a9ab1d744f8c0038c272339678f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h878fc86f2115859eb14b35b31d816b594acc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha90d1db3b97b223f5330e6ac9b20bebed714;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91f7e83554d63487d7bbd6c7f11bbd827c9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce36205a661d8ae2540452abd5c739614f56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e0abaa4c73dac38e72780c824916068eb8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf71a11395ec7d887d8ecaeb0b5b49fb78fcb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f82cc6ddfa1cd855274d983085a63383387;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc825c7b5dbbe47b1214623ecb05b82037ee2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f2d261fe334dbcfe0a92b5e3007495419de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe480b7691131a9a5d389b3841f0bd0755f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he939d57fe0c857c43276616fb7268b3a48d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2acacfa63797efae2ec004c12aa03aa97c05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h122864b266539200027bf0eebfdb598b31ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd8e94b44fc76302cc56c659675277228bd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88c103b4a80ae643bd476e84624d9248c48c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8597adf10df6c6077e3ff15d2afa96177af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha23cbbbbe8d6ac601cfbf96dabd400f67b5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8ac3ab391d4765e36047d6b02c0cd771d85;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a795b41b01da59747f5c104dd10a955539d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2e806b34b0830ddd6ef78358ab940e0aad6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19e37e364d01c76356bc23095104f2bf3a53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a742fea15a857b9f461a41edebda3a96e01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77d784ce0cb19bbdb630fd6d53201098e55e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h257eeb984e574e6aa3490980ac3dc0f4b956;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h598755003c94adb4f949012ad1eaed0094b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h705ab3076186ae210ab7d6f51ac169ea32f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72f4421b8dc2a0fceb312cb430d1a817c7c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1267d65835360beb662621c40487096c6eb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a4336cb1ab8ffe73d4b611014ecbf480638;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8df8f5488bf6e70f463a1cf2f7e3bf4b296d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb13d0748c4960f1f681e6d32a50b8cc3268e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e84ec6b91b021c4bb9373dc7460e5638d41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac299f600022126ddede1e3a35a1d243dbad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49c3a74e461053bcd0b6f56334eb2ff2e499;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h831a061902988aef1ce1e21eda032e7eccf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70b3a422a702194d2b1c1ebeaf9dcfcc8141;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b2bd39ad2917d0c161cc4e0d6d50299b99c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hceb7b7d603bf066cf16144b171e33207d075;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe462494f96c4e148b3fd5ee434ccf56394b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39783916055af8abbae3e0cb3ada3b5e3911;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0a4352580336f293df9a7e30e2f790fc9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2731fd1a263e5749c73cb88a0ab5d6589a7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa6c7324465125abcbb3be6521c950b4b09e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d2a58a9511528e759eedc9742c02da7b23e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1502a6f68eed1861c02e4c8d356edbc8d08d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c42bd40248c2df314975dcdc3f940523a12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb951745b8a5e7eddd8a1f8472059421060c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd783fbb1ebdda19f52cbbdb11bacf7fb06a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd84010fb327eb199beb62a5f45b243407238;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h201d95c42f91c0c85f2c44a3abacaec0b63d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa9b019788f90e2f17fcb7038914160d6e97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47e20e0844d24aff6ca9a8b28ba8c343f7b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fd36e5df30f51e10b4482a3a7310c663551;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37c9aaf04b8a5462ddab7aed528b3a660c17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h899f51dc3643a3b1e0cf936b8364ed78e097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57d2a21fb6e11d0c3078095bc5758f02d3a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h692da78faa5ca5c2470d4794be2648661064;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8686c12e910926fb9bb1998faf0c9182da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he982b07057d89c656a8fd9ed80e0bd0f6f8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h611ea150b7a09097f1a6fce9f59279c4178f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ff532002654da93d2192c762dafe6aa87b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa94aee45fd7dc5384d76dec3e835a759d51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a530bdf7443b216e9d40fd88873ec2b3ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47ef03f4a9a37dd9789fe67014f8831a421e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34bef329b2fb0f51295248bba110dc9cb6ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76466b638d39121f499b64255a2ac787fef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac128d76adb00bcaf86b221378dc21dc5cdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1201192eca94be1082470068919d68a0ddb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5124473a95f77bda790db4c40a4b7b3be619;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8d61870066be22c159b3012eedde763bb01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4576dcf270e2973c910876074c65d4940376;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aaeae9a55f7f4d2ac88287e955e23cd8429;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2889bb7d2677efa1762f7278debeb1e17dc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd79a401ef7ee1462fb1080201bbf5db5a330;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9212c9536322a56756c5d5cd1e08e9b08d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a31a07523f67ac256d22667d9df2534aef6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60b459200835384f7c1a89863d4cba0fa161;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf195a44c3294b676f9b6f06c7dbf1a708906;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb073c1413d7e8955f6fe54b098d58cfb9618;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc7e7b5aaa2a27856fb9b8f27f86b0f5e6fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63f3b437adc0bfc5bd201903f662410d3d60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26122eb82eb9f1692ed928b23f32358ae0ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1def804d03d7bcd797b1454d18c8964eb4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa8ecd1d02f3069bc42298e75a91a8e5ebda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43e02e5413cbeaf9621bfd1d26afd92e3fc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aba3d522f254e2065b1b86382f50d262b9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3bab101b64b8421f898bf4e81b46096b252;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h175f9d567ccdfa5b2c0f3316c91d6e644104;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7694a482367f1e5d6e24877260423704629;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86423d74c0a78f2485d62c8f6cf46a0a5c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4938b07a796f091eeb73c04ee224421421f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab93764a6636439057efae72b24393c7b277;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bddd8b6792c9d65ca181d2bf66ef2c33453;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9eff1b154ba2f50f94bbc1ed0c2cea028532;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70a75618529562d77360050d9d53d072da3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h862656de214dff05bc8f421af3e01dc2811e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b0babe8af277ebc41b01f6622b817f2b6d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ad80ea3caf193e7a99ae6ef10b2b95ee216;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fa104e7e6e1dd352afccfb466e1972c96e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h825563f1839c381ff2da814ac8cae0b66631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf61a7f281743d2af7e974c1cc8362a94088b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f4e69f9384f318a2630187bf6bfc8e90cf1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25db2b4cd72e120eaacdc5f32f455254d00d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bf4093b6a33165418962f36fb12cc49e890;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h505e2e78badcf233360412f4324903f4eddf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcea4ceb199b3c2a37b5575bea75f0d02429;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heec1cbdaeff3a4fae35569a755e285d8357b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fd7a91eb407b536fd68082337b32dc44bf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdbdfeff02d227472564163b36721ad86a60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8acc326b84bdbc45411013669a3cd78213ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aea611165a82f0be38626d1e1b12d28aee4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2da0e6a453b1ac65ba46f5ea76edae471b07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7129e8faeedfe193f1928d28f2367ae55b82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfb1e1e80d3a868d0fbfab82bc90affbb8e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9165447f4ff6d0259eb8b94951276b685e83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5bf32d07d330eef7418454412515d0b521;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6631bbf5433ddc5fc1a046f1348747b6919;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd14cc597e51ffa94993a3b2adf79809b8933;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f898c322c32cad987c95f9c044c137f25cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2f2b8b1f6bf521d86b8541c91a5a4bcb2d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1382ee4f764f917bca9a122b1f408595b849;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hada716aaae52340837e2b82ce30fce9dd79d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74d23ebf05d0edb6776e6d39f5d37d1c036f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64f6c4859cfbbe455b8ffe3e5b8174e59ea5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d4d031eb166165396853335ecc703f3c4df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7507283a973e3fe6fd75027b4867cea7b78c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc9578ca8e3caf433ed8b55548c2b548f00e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42333c9600c5e25b75ed25b207c2d54fc558;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h657a34d27da48c2d2dc0c1eae1c362603d1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e06894b4dae3bdd6c6dd5dec1eff8b16e63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcef8022c58c3ddcd20a5e3f7a74f9b737f71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d1f0a107568e58a95b471cc1d74fadbd093;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9035500b3117e3ed5c1496a2d12426a07881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33001dd70e450eadc83f4ffb679af3da4606;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h685aa4e8221e6d55cc63fa976145c1fbcec3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ffc6763d27ebc44178d5bfa5ce740dd52b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha837223b5023ae902502933e6f2b1e1224a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f80744acb558132de0e97a30d7aa7715f00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8be9191430f110bf79cfc53490443ef6bc91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h946e84fa6c82050a80a008f1b57162a12edb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2726e8c3a120b7cd18bb474a3e538d0e844;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h885566b4508a1deac53c9cf394a0e2485485;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cd0b1573e13eeb82f41703d52a04e8cef41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b967a3fe587ca869b593b5d74791389f9a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcda7ab836b7ae56993606f4994f3eb36c67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62a4e0bec957d268a61a74cd108eba0c5ee9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86eeaec4ed814a55b3584940c811d162aa52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha358cc788cadd247396f02675d6b8db6865a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf350f83800ce44d9aba06f3873a03b830a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec62f95d69ac934b499d9b4aa576fb92ae15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4960669f6a961679f1832324b72d922604be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56041ce9493a2ddff44510342e4c2d3c778e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h302a40d1ced6386faf862300bd94b9e537a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef338bb57254750c60eefd56f710d7d656bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9da677432a8f285f69e5d3f6fd81ef0c25f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fb6cfd0088e46c369097f3d44f61edd0ee7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5cbff21d6a6938c3b8c4cacc7999ec5c12d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bd3cb1aadd5353d96bf522d84980e83bb62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9be45cb5e285093462f195721178901546eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he925283801fba57356d706882f63f7fff108;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6bffd126f038de79449f8578aabde03de1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b70346dc8fc615c700eeb2ee16e7718d766;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d769ff1a9c7e795257ad86d35df708047a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee917b31b57777364a5812751deb8e2271ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd390af275a761ba32e72f908fa6e4d707584;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1795cbf089f76c23c074fca60c7cb871edea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72061084cbf80de951b570b0d2a26e33dc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h414d79d2c0cae7560d01072bd19319ab2982;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7112b993c22402c4557e92d47202cec38847;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4aec181a9643e05536f22d1f2bbc11eb7c29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h999dc0b73aff74add529a964538c3f176927;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bf2159273d080c758354a63ff4b45eecd46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77fb4085d1cca4bba7593161b1cec4f52a9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77dd1287c5ea0d1f83178a5d8b83274bd07b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3c176a8e149d576e0265e6fa2770e2ffd47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab8aa4bc659155ade17c9d71677643e5c5e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he493913c10bff99afd1dff9878f262bdabf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fc85ece5617afa4e7d58b7504bbf75a458c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2180a127de807122e6cf2a75e739532b681;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha647fea83cdcdfb071c2dc58b95e4e912f25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7984a4eef43d001d82ade73f158a90bef3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8381ade159914eb658b5f3e725deaea775a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef435265047034ff542d0318eafbc01e171e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21e870d592715f54f29142e8291aa1aaee6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4c34fc2b27b0c88e1577b2ee902d0208c3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha515dc5e2ee448739873965e67c10c20abb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h781dec2fea89871fe1ba1d344460c9cc2573;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb02446f1408e0edbd1172fd52e73be8f23fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45c490fa51d805713245c299c3829aa1f2c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb708346d0733560299a51ffb4932c286cba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d22369825537d2c5bd0bfa1f572594a0b8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48922a04f927b6e62fd4414a718cb0a5e519;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22d73103d15ba8bd17deb7a516112b7b76c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbe29f8694c35c4631c9868a84c24113dbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5b8972055ea739d966967ee75d5e5bea96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb313500e9d2df59814f47f63edf6a07c1fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffe705fa87460ea35d932a088d796ebe7b81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1ae52e64872a1e4b1245f1fb5b637f3c383;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf84c623943a0b570b32d2f8c61abc6f56732;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7baeb5ff85e2f2c517a0b73d4c207a62ebc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fe1481e4bbf6280d996bb61d36b694be5f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h726d1e14710247b1faffdc9d60d5873cf9a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h751879d0c8aeaffa69a3932110cfac1f5fcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f6d8a83ba2d6e05c8a8a8e8009ec31484dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h708d76e52052554aa83639e4444b56afe87a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf26436f5e17ac697e0f17a782a44e87b5f46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ecf16730d8ff36b5fe5cd44a0e30c53564e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6920543df3d2b37a81c661623697ff759b5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6844044e4bed398e4972585e5b68cc0ba617;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d0905bb275a76d400e98eca6a6b3905d0d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfbce3274c9b5edd432d20056441b922940a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd9ade58ce78a1aebb65ff5a17166dfb21c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha92eea9c36f93e7b5e622cc90c57215ab8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71e1fd895fd91ae4bfdc486ee53e15d4f144;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3220bcb738f3b6476d8118e30c94ceb2cdf9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d965bbbc81c864a08f56deec8abf26b215;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a8d5779f2cc29645b47bc8b0716fca66400;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf4cd915b5633594a1d149232fc536fab314;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac668ca870f842dcbe8da10b375e33f846da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67e5d71a0a6ce71cfc712e78cab18b82580a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3419740517516c5e1b6ea1ddb6e9a8135e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb1d3fe8783d616c9c9ec661d1f780c822eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e47fb7f9f1d72374af8d85317c46988c9c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd72685b588c5147ea58e81275052cbde299e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c54261b132469f194ff0a7d6c6c560fb5ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59eb72cc907d2da27e35e4cee25d912387ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1efc8787f404ffc46a643596d419a743011;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f9cde0d9f2202aa3614b030c8caf6f4a35b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3586f20c50c468a1e5b9907c627c191b109f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h663214ce765c4cfcce60b08bc7fb13f7a280;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56bb8e6ee9d94b8d19251001ede9df3acdb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd4838c87b26b4ef69869e6c85f7ec30cbcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64b4d9c70a0ce092e1510fbcb4fd8867741f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h143186216b5b51f78e0524decf335b7001fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fc924741b39b1d3119ccce5bab2547c205c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha60e3fa4916ef59a38112562a7e9992374c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f7b85ac55fa1c63a71d48212b8c739b01ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2335399b1716d93872e5914ad868107949bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef956f8a24b514d58c378ee28ac82a6b4f7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d71d87801af51da2e8526b48ea69380dcc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c791b68df5347c0b70d88fd0e8bb0dac1b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf476157ad9e78ac896efbcf760be6e215bf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h521001771f70a024411358e4222e0346b194;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e70c70d409b59bbbe7be97f6fecfbe3722;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha59730bb8989eacc4c9c382336bbff05f82c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h369d54aea6e54f865140a218984b9b6813e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24e4aa56c447fd2b542756b7737d7efb5bfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdbd51895f657dd988806fefeb0d86878fd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h211357319a6fe2f82687b931e044c41f70bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86d3593ae9a3cc3bad82338e431288b23883;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd431c846350cff49044c5757ec53a3cfb1f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb37922789e96b9fa4fc899feea07074b12ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fd481f1e650731f5b5047325b449089f991;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa11f4b62f7332b0a06cf57ed38d66516489;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd43f588fe9077070c01cd6aceaaa95fdc9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb94c787a27b33502c10c126d2855a1d06f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf340e51e0ecc4b652b7b30976ff5d1dd41ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57786f4aa21806d72082b7a3d2a44f197768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h563b81b0dc784b23cc55f3c08a42f930d2ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eb886ec7b5df78405bc609992228f53b16d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5848aa74fcc36a9f99f4499f67a04769163;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfe007b8880013d9ad33b9cdb745ff94805b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf11927df53d53234fbc96f7dba4a1dbbab47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf2d297011192df81e2228c1c4ba93df6d80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8216888f16bf565338d9fe2c92eb2de8ed33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f5b82eda04a76e02c5ee97f7b2ad106e9bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5922cf49776ba48ea4bebb209e3c82c29d5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa76ba543f73b2f61059a98d432e7e1e03b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee981de33131d2ff11a64cdd0549f49264af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4d32ba8efcd6e9d42b30aa2df8f68a41afb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc66642da0e275e7ed13510dcb57b2aff3007;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h877a060413605181b51d91dfec5dd7551151;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4c818309c2ce6ec82527d8ae9f3ef74ced6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d6c8b598a7c113304b98753ae4bbd42e8fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16916136692b27c22ce7bb50efc869423875;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29a6a6c4767b7281d366a6181eba56d08e0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82a48849da17f09721df0c08d0a20fe2c39e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c5755d557f04eefb5828fde91fcdfd42e15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d2a7480c97e23683a886d22aede2b3c8932;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8b8146e2666707bc5651fd0c392713c6122;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadf0b34e0bea96d2d1bc949d2be88bce097e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79696b0d6555f5512b8a8595931eb7279295;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc43d46cfa1b808583703a45c85f23759a227;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40556329c653c73c3932a7996b4f6c9a221f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcaf11b70eba0c24f174cf09a711dcecb0b24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h922a4ac9c8344bf3154f32b462c57eb8c38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd75163abd567561484c86b0fa9bcf60a73ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44754a939d20f57f75fe742e7af17a1cde02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e0b5e3cc7cb73c9e439688254f2e58933e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45986f82545394a448dc25ebe9607928a48b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92bf7e26a06e0bd29de96fcea08ecf17edd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa87f18bea6e0130ac9a403b23d43b5561d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f10baacd8caed944f917abf09f62bc25c93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6f6ad7d9351faaa8510fe767aac998d5944;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h893d3628aaf81b9a85e6ad081f9ceb7f30aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96d30be1d7f78d17c4e2dc7ad793a605e3ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h711c3cb83ce7d137b454a12df96dd4050d1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a693805c97df7806dd96350187c21283f9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0049d895e7a944447aa2c4f6e7fb88d2d36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha228a34bf4457e700f4852becc43f363481f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a6a2581c15b180d77197ab2822c6dda4391;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he441f3627214a724a0c5409d07a3ab6561c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ce09d1dc983dd7562b4c6aa8ca233b68cc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63a6879e92e4e39231240557eec4693349ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5add75b5d5c21b7cc69db83bf2e9d8fa33c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h882abf6cedf46210c472e5cb4e24bc74c82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40cce59b36d2aba63d00bcf41b2e9033477e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha33210a1a8a1482a8c8c3dccd143ee2d1af3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fdc108e4227234423863c07c50252b0bbe9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d62098707c91c72c0ffecdbf5a715837227;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e55be373161a592b7bd91fbe21d7f102fd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98aaee7a15ac2c4b1ed671b64949f31b40d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h524df96251b12011cec118023a79156624d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69b7117a07a6b05055f0b02f2b3b311277b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72a9c7b7e034ba4669fce9223a6bfd9f4b90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a16eb7a54f0d6a5f8f43a3779a977bc918a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a52aae245bb88ef9b0304df2b9eba344b36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38185b4ed551b98943e00dc09aacc3c90306;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68db32ca41e55e4370625be2886c1bf350b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a2ff8b9aec4426abdd1b1ea7db36df9932a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eec326ea4008483be2f41a0ca348aa43112;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4120d7afce507ca67cfcdad095188021770;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee37642d2e1df110f63fea51a0d0b2af0332;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c11da9cfc2dfdf7d0b5fb03da265defe645;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h473dfe6d2a3d101e45976b28c4d58d629ef2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d2f6473cb1eef562d07d9ec97b6444fcbc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8629118a3943eadad577bc78d49e13e47d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h141a6701ce5f746597d4238f8198ab14feee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf92240863bb1960a542235635b3451511b95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h136c4710e4fbe72ad137a4a7f15c13c5ea42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdda6c5f1d597d9bf3202a91bc84ceab6323a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61c8d6038bfc45f80329ba528c3c70d914c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8be4a244b17afb1bb381bfc0220b148d20d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae612ec34cd53be3da81f30b076a9d8030d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef374b481004dc5f04eb9b870ad2798f82f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47add6037f8c88857e321bd4de009aab24fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd893aec545e1cb4d0f7c3dfb02bc4cf9f771;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9faae5938424c6ac547e1c1f73b766522c35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81108960496e053315fcf62c80b0d4b4ff0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h643ae3082ce24da795fb239af9d8384b6bd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c1219adefd33951f97e3379c3f4f756ecfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51cbac3bfdf4dfc76008409138bd2d639861;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h639d9e87931d6b130978b3adad918620a01d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6dfdc4232a5721a2207cf22967822d96e5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h306b0c9d6833557be7fa182ace699459c10b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa642f43634ce1ab9c57ab6212eed8a0eb3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd01d46a8e2680ee9098213d0d446dd50f77e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h293a99d9dc89409a25373ccd1ee8443cc60a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9265e3fbf83131681eb92b32667f3a6d802f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fb776d633612b88d00fd588181020e9c2fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2c99bfb19f5141d06e95798714edf5087b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84c449e34b8e27235f28bf4be0e1df812e9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba376cf1914de7eefc489d76843a5ad16ee1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa89c75a468de0cd647be379fc2c30ceb847;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he109b9612bca3f083e8b957baf9c8601514;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3e8f7e984d6acbe34ddda405ca038947437;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cf4994d68250fa178f41b987550c2bbbfd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5ebd97dd40c945dc0399ba906fd3d4dab12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8a2de5a83020d28c5df456420e17de497e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9284f4c2045a35b4f95a6eeb076af1e79046;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8a71496f14c399e5137122a335a5f1dadc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6528b69134240772beadb0faee314241fac0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6b81f6ab8ad620d3a106b0c671d06d31f14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h494a0b5eef9bde5d7d0973004d578d495df7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59d566dc2a01c2766569d552433e541d5e66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa0d620d4428cb2052669f40332492750998;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1fdded44d7ece75a561d0209bb985133e92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc1bb6bc15a5e467731a7103120b9f59961e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9ae26cb80281dbeba2197d7012cb55bbb20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d42bc13681604aeabe3779460b05c073e83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed105eb5c0e491e67446b8b99b244128a0dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87e4e0f379042036d9619b2d0d61c69dcae5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c29fdcb48c653a4f6108ad8a8ab394bfad2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50fd6d1949220db7d93fa234ab5f7f1bd77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9df7505c38df5f004be62ee96f0e7d8f9056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he741d97fbb2c59243e86ea33cb96b06f7c6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9614266d5b9b7284211a8193c7b7ed3688b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6155c738a75d12b9c79053ae13020660f75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e6fe43599bc3a3dd2da879132cfd0011f90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdcdddf0d7c9a58886b17e7353d71e27bb61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h647d05c7ad552ea287e75e6c64f3e3ccef1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bb3eca60d826f64854e7b8c881b0ad11ef4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ec01240818c4f65d00e5e83616b39ffee4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2c5d7a0779fa779e94d4d6dc5248f0821bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb77fdd494a1cda7c9d246374f0098c5a7ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h363e2d615d1a7039fa17b718e2f6a35cb780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3a397f3ef646d90101ac704a449a582b6cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35ec8ea541cec4bd064e79317fdc354d5e8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h728e5ffd4280333e71358311cf217adadfd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33419edf46fc7d60ffb7c64a5836a18081eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9875151e4e412f051f2405da4c7f9149cacd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab64bc8023a576bcc43ee79d118c8f004925;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc75f726d0df9ae1c5166fc58ef5487fccbbb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93031aa7faa311ac55532d87398df81d49a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93722665019bc5e5bddb637d9124c293e38c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3cbd6427310f05375e99dc2ed7ca8f53a1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a3a53d94128128e4f80c3394c85473e78c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf0633e482f3ee595e6946e20df9ce26789c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3b6dc578604dea45988e175886d1daf64b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a34e71bd580e293d25b67ebfec009f46801;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2e2b8b1d1bf63a9194b2c9b7ee4e2f95c7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2ddf324393d903c46e3f61df6bb9515a876;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9335a03159ddcc12ffdbf67c6986a30aaf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d86204e6249ca8d6ae8d64e6b55fb2efb97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h270b6ea0c476c23bb21afdfd48a47cddf05b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b1d19a1c994871c960db779b94c8cb9219d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h175d8473bc9b6fd42828bee482d6f32546b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha26f077b3bde4ab5f6b14a0f0841744c0caa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha888c62326f0580849feb2d0ad375be9e6f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff934747af827a20434450122b354c3dd4d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e186c1523454a95a6cbc62ed82217c352ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4b95edab7290118b6d1189d0baf39570d6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd76bae5ef605b2e3462ec9e0cb06a7db6bd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h498a3dfcb581936e295ab19c29fb924601c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haff920918b4cb3e127334cea2cfdfd80355;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f609bd4242a44219965864256ba1ab91a97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56db162174785c5b8f9714d95bbb3d8502d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he44f968a6edbfcab7620db219ea2f1c89789;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70bd887e1f28304f1c78a8d3c5ce3d70a8ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0e016e9136ed808739a57e316c76a7e3382;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60e51fa792ca1ea3722a25613bbc0f5e8a16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb04c3ac04e7bb869d590e1c79e3b0f717a13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58968a90c79a40ba10e77b81bd35a21c9d9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfe41454432730b6a13a9928afe562a77e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafe5822ffdad3cb1f4936411e7a78a752cbb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1727c4bd543e62cd6087eb5585e29bae6794;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfc0f3aca9c85dbe0783e6200491513003c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9aae4b3f9799e0773f34dbfe1167e0718850;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a118e691c59fe31c7775d255debd2222aec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he879620a336f0c3bb4d0d1e93764c15c58b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb42832011cb90dc472b271efec6246568bd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc83a669b835ef0ef75ff5ec4a49780bdb412;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf9a2a09c46649a2d24a32c8fc4c80e4ff5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22051e4e7672d6d8f28ebaa1b32f13301817;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde9fee34680d61cf973a01c7c51d8267c53b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4f7ba4a1a711c01ac1ab22fc663312abcf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0a73174ef42547e6433f6c7d0374293c6eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18543b7613c410bede947ead11ca629f549;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9288e4334734a89a12e400dc477b1eacde4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31e21ebf7e27884ee29b04a3540a69671ca1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20b571901249ca96265d3cf8c1bede6e22f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h385be72973df24914b50c0c0d7006919f972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81c8a44fbd50b89a929c41d6cb0fa5dc120c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefc3be897ffebae84d69e90ac324acd7d47c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h551dca6775d1beed3e75a04cc3b52ccabb11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe3180d267b2b478a8b4dfb6b87ae86e8a5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcafb1257b3c99335410594faf8a8f69a926f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49eee0f4fd42ed6ff55a031a57cefd51b436;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7da4d7e73b0317b34ed83b75eebba06b5313;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f0a157cfe22571ad753ce43c27c99bc525f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48b234d26c95fd8174dc4e1c455bb9717db4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25d761dac69555b5a637bd1335133ca2613d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1eedde6c035b538b2a425f903bbe84fb5326;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bcf70438446de2d60fd93d4aa75e23f4d02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccd11012f31b424fe1dff11a00339d045de2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h619e9fd6c88ed88158e9524ae7f89e366ab8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd72b40ed758604ff2aa4562951ad349f1de6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc83d09f8759c16e873e1d0c686a0eea29196;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h134257cd2d8f957f771469e633c5f557df72;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58bdcd389aece5a614a05dc1a149af562f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h978a9a82a1530bf2d8890dac77e86475c014;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf80522d7214694a20f733d7bed1caf8e3c05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa725eb5abd38208b70a27a28e7850529173;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3a21145f4a5f9a230c2c25a99da8df9f96c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5f3a3c1997af8fa8d7c14145b8efe49d636;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85bd714a399cbf05d574d0d3b592b5b3d85a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e09e183b325ff00e1c5022f9e9335fb1bf0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4cebd2857a971d25ab582af278ecafbec8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h654b8fa7a80fa401e2c1fdc8c25b6f6bc03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3aa08d55bf00728bf0c399af00a0c98f6bd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3132f1b701f97cc46e07b3ee950544c0b0fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9de4de7b4beb2ad2d0206e0df0b0a7ea2f4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h793e8a6360f0cc92670e0b5a8d6a983d235e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6720f93af447116769b34adc90cff7b77afe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a4f15459c65f97fd019f1b41bf28798e329;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha41499cee5629011d3e28b2c84b05ebe7db6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e9b473efdd90d3e789333eb298591760dc6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c722693817fe0429749969f730744ee2689;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb154ff77cc83f11b5e6b134939c784ad4b60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fbe0fc9c86c3f44f3f50e1b02de9e6b20f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb55106525a62fc97b2862a7ac1a7cc25033e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2456da6e31197eafd42164dff0689a1d33c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0d4fb300ad640c67a089f25addee7580f1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ed0860d3039d85cbef8009982190579043d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc68537a9055b18004e2b85f9d9621bfdbead;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cce7d0078e47a16d0633572aa9f5baf0c04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb92912616e2fa2f79912c5346ed8d4f595d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6caa9abc95fdc0a7e1b43b68d10845cd565;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h722ca058262c071aeb7e8f1b34851cf0199e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25238eec72df4c2a72235a2b97f8bee42ed1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd35bfd8533411e50dac562c1e05bd8f20c63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55b82691b10a11514c2ccf5a0ab5bb19c595;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h761606529629fdcc5c2fde5e951a33d19028;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ce643aaf55aa7facbc54f50a4adfe5180fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97e31dd5af1f8ddffaae7f069c06ce8c9a02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h151d19091404585dbf2a8071001849fa2eef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h889e99288cd6b2154095734ad0d54df42e42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5744eaed92f35725c5900f67399039619c6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdb2f7f5e607a2dd47fbe7272346a3824b01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha00c404f5af2c89195064b6b4e7e8cf0cc32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he144b3c26fa2b12d1e59c216d8ae9c11b0ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34821d27cb994a7662ba84295dfba3248cf3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a2c52930b878695adc67b31f560f92615fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b1ec4aa8ce86fb94ff6ffcd7685d86a3784;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52b4e511778e167e9c78f86452928eff43da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd56b09e52f551c383937d7f7b98a68179e2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28292da068fe365afc579128a0d61b8361e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8aaac42b29ead11df5f5c4af376dab1efce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0da0b4778649ab72fbb3549636e40810db6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4405b91e13b72b2a819e9f8dfd60c5444c4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h437637d76e39d24b0eb6aa70bfe38d3d730e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd398eaee44c277478d77b4cf5ea2b421ff3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b27f22d7240af931beeae3a609d0f08d9b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbab94dac10b1ad238cec42eeb01eb1abb2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa50d24637e944bb510c2525b76decc4ede2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85dbaec2c3278880c4b5eae9bb6351aae338;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h364f01d9988a1d20635c892080b7985a14ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca19443cb54de8b38bc91b0142b9f338e792;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb80a5ce72cb50e7560cb4e6cf7aa7ca6415a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96c552d9247c35efeab81cab50e22eb613a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91cd11c8e5e35cad7cfbc6be41e3095b085c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9659c9156a1959163c065c30eafcb1405f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf1eb8d6fc1b55a9f725565ba6a7535d1d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h927794be970e897da93f82612ec3a1aff8d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha666cd9bc9138e735ca6baa91298de11bc42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b0c9230a20aa6c3f54753391cbff58333da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68c72d1d7942921ae557b3085ae5fbe6967a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54d51856a0e5a00ec7ef5b2d16c84e2150c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc10ea2eb5f015b0e4f10958f96716e774cbb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36a2998c6612a74c787b112638267ce1b0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77710efa2c9e5ede9e165ccc861f0a3f7a8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90caa9c6ba034db7bacf7799863da85563f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c1a6223e754735d5b0e06ab9fff6caa703b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6415ee95c644253e2b4500a07cd277681b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9ad9a17f94498f73c51101cabeab7c96546;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45e7bf324a04579a2497eab5bbea0654a96c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd801f7dfcbf62b47a5e1f5befdde8c5cf0df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82cd17a5a9cd478da21bb1eb63a98ad48263;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8113ee642d5ff935135443d9ce898956c5a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he80d1e29264dabf0c190241a95af08d42db5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc471290a620468429e87454bfe18f2711d91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eb086abf40c079564d75c1d390fabd4a901;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6263c41c2970ab1f55c9e83795d6f9d9502f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bfe0d5929c4bfecafa585933a52895aae86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dc08f276d180f3e0c1c197e725d21dcd03f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h756e31ab803dcddb346a0d2769c2e79d76af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46250c7226d7764d22eca14e81910edf8f3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42e5d34861fbe54a4367a0b84a796993da3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbfb2aa34bb88edc445218eb5df6f9030483;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7da57e77939bea7ede39c9329ac633b89942;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d616539edd53b7b49c2fdfa3dda7a696ecc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h444a1f9a4e69a75da18161563ee8d7d9c356;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5450e1ec52233afac270bbb8e63ee1f8e00b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18a62e8ab498f4a792f6424070b2e383dd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f7faac2f8d9bfa4aab8be859211c2ddd68b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d85ded9e9510e5fc46ef2f9b605027edf35;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6680ce1dd6a81359bf3b1d0311e23ca13b4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44ac17e67ca1fce13cb44c25e967a3bbba83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33b674bb9591c90a1155e9c5dd265aa35a66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8c969c3aa021a40878e07769d16a9700212;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe91e0d80c4d2c1afc10e83e86ac024f4ea8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4ea02b1d880d67d0c8ba3e64f8bcfe6fd92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc245da3cfefa10e4ebfec5d7a6605d1335f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b64d208dc29020c95e2b46d12374e5355e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha09500daed3e9d42031d377ceb33b310bc2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaf8e7159459bc4f7cb9fef9871853580452;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c18793b9da14256d2dc712c27e86cee129f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31c7a56ad4e71c9d3b995ea3466476654a6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72b08ec7f36b431c2b4a6f462f70c0a8185d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7eba7fff3e8be11f60afa105c3f9c076e03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac11aff268551db80429bdd4475bd2fc2083;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h880054255456d9d4a7552a785175b150db7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h715d7d4ca2adc815ad8eab17389be6336721;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6db74b07efaaf9dd8ecd2de195cc6b299ee9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h285be6bfd8cbd76ae1d6e1c663026f7c839b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he166c9c860d0e9bb0762ae10d530f5921ab3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb78ebdef114f0b50bae02cfc40dc204d7e03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccc3356cb66de76cfec9912067ac6cb20b16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha64134e14d9a6e42a0f953e99fcfca40fbba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb358397c885179c0949f2b0dea073dbdee30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12d3a0325682d831aa8051823952f08ec579;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7d7854c11bf85776254d7d5ee08d8781f5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93a792781c4a2578abb0a25d1c0a91db7860;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aa54390f5da2c55de6566fe8e2b0d20debc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65047e2c074fbebf4ee23974de6c45af0f34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3926d427fc6f553d98bb4a3ac0d067203a0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41d5c8ed0e945e68858a60232723eb49137e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63f918364b01789922c292fcee04625b60d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9630a5847b7e854b49e931579344ab122bff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedc70c568daed2781ab724c43eab28746b6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeafb6a8b7f8e20e28465f42c6574edcac7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fddea89df903f794aca403a112697e06aa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h233d672c35dc7e166b0782354d91eb432c1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h225660cf1f10d8131dbce23434bec89f95c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6a740892f11aa97c67d4f91c83bf4a97d78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54b8c4fc59b5b6b73f19ac436cc609f96d6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haef46cbc259bcf3d471839abe5dab3164f9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc5faf0e71c3b4aa4830af77de2e82a12736;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b238bb59e05496aabb5902e65d2986906b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf035fa0c7af9277b30e2da298f58de667c14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37ea79b2a82e727e59a32d05e56ff0ced6c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72ad5d48679061f98d1fe0b2b5dd4add7d45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61207a9ba1448d344ec01e226af149119f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b7863d2885772fb04cd0ce5cdfd2fb593d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf41e22eb298229baff288c7c733c08052ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee28d4e23e887cfba2dd47dfead3a114a497;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70198b14f55ef9aabdcac670ebba27e43530;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf59f1de0f8fb22dec656bc9f4775e29d78e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b9506787b747ed61a4b02244d8b3c2d0ba0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb34dc3f309f6e2b8a4e598e4c34ff590972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25a637449be1c907a4cdd0955f1ee2963747;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h635e602386745df4d3d7cb3e39ff82122a71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde82d262de70fd45593e01578f764073a7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f583fde0ef9c05d5dca505996c6fba28ded;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61928b9df818d8ab020ddb7117ad1a9dcc2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1471b771191126f5e2e92893bfd4589fe816;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h919971785b03815eb2366bcfdef5c5b605df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb4a55c8fddbfa6a22a1c6204420043aeacc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcffed6a08fc744694b7e3cd274ad3c4c430c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11bf38a03d4072c4fc2b834e94a9c81da9c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cafe2b52ee926f0098205733d6451a9ea3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb74f0b74b5c05e9ce73f5ea1119d862ed6d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff673081f4c804c8f4029f03d2b8a43909f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0654a5a9d1ab9b38d151c6b5aa34083a885;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h848d0b4ad0f2d5596d232ea8fa0eb39cb62c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h669d6495b59f09408f962fd1eed1b6e4d52a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1f9b65feb66b9967ebb60e8ac8b4a59d351;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd827859c2916e01cc8de1c931477ada1ad9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2895ba4f988f3fe9c4ea2da28d8910e56f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9297afb9747289eeb657f54a60b7efdefe81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f8e3b7747af58e569001961d6238c89be6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddabd94f39f9d091a17a47d82ad87304c9f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80640dc3c5a19811048da1c6a9a614996f87;
        #1
        $finish();
    end
endmodule
