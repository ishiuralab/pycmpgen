module testbench();
    reg [16:0] src0;
    reg [16:0] src1;
    reg [16:0] src2;
    reg [16:0] src3;
    reg [16:0] src4;
    reg [16:0] src5;
    reg [16:0] src6;
    reg [16:0] src7;
    reg [16:0] src8;
    reg [16:0] src9;
    reg [16:0] src10;
    reg [16:0] src11;
    reg [16:0] src12;
    reg [16:0] src13;
    reg [16:0] src14;
    reg [16:0] src15;
    reg [16:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d318f689d8e8aed911cb4acc7139785bf1bd0a1a7b957a00cb36fac7544444884c671bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1372d524978b373b0af3c9936724c870dd10d11c5492fbdff6acef7833e4b90d4849fe685;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16080e8d2065b115834d34beb0f0235f327997f3faa83a1a6df09886364aa7f456b8c226f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14976a06e90b4cb1d2f7a392a85da1cc211cc16a594144b1b82f9ccc05f01a3b890340f34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf81d57269bc35cf6000ec29f6db3275fba2b6a9fa3114c4fb3cbce024c3dff40456437a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e91f313ed44b26371796ef5647d8b0ac46d565af3048e77b6ae81faed69d954a0415e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd88f9d558610015a27fcecfcf3ae7fc299eca892d07180eaea716f37f56b1f68af25c5ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158671e0d008b8a27e531c49e2e0852225cce72945881a43f6fed73bf030ce29c9401b386;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae6f72a767ae4638b89c4bb982453a555b7de500af0f8a396065385a4b203566d31a0262;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3712ad469f6f0ecd41fd3dff2247104579ba1f29779aa63a9ceef709475ca0a81da5531a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6d58a43f72bf1409629063681ccdc6b1774d0b3f64db35ef9e81a98bb3ac574ba6eced8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71ce7bce591ed644cf332eeff7622154760864181b6609c95674c8a4ef61e7af728931ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112f127eaf01fddc21cdc7732cefadd121376107be4cf62c2ddc564fa6934adf687dd864f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1495efa56a28a4821b7079ee6be8e259d51bd1c3803fae8da2141b5218f54eeb097b73d27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h291051ab456804887ce751444acc789d2054805671d836c1ee2e1536b115df34407492a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h46073c1bca163163ef8a338b53715b19d2d2c7b8e88b03095d2abbe8dce44dabce1b3e0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1568d98738f9fce3346d65e99e05e0e1415ca925f49484638966a338c8f27c2a69bc3799b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c797120f111eea9a9b057d8cef38177adc36f048b1459aa82c4d5dc8c6c06f3881ef3064;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f7d9aed1fe61232ccdbd6c339d54fe93e6d5c5ee8b359288e8bd95a70bd27bda9911167;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38c0b12d9391cdb5f3286b6ec7403edbb5ca49d50937116863808c45edba70454b33ec06;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133e2eb1b2c442da4da255189ddafd1da78ad9ad2f259c2047da10f938416c56e68915bae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1049f3e99fbd8d68f5fc06abf4035b233b5b8fd20a57ea0666664c75b4120e4430b946f33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19844be5a2ef2dae876286c2c59d33314e25b61f186b562ccb6054e01800fadc29cdf0014;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61aac1716ca85813286b2531a2171dc92389a3005181694f6947b1601e85d3a8e3038af2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1802302e38d12ffdf0273a5052dfe10cc202a7192a11cf7a9f64e44c60dbb97739ddff01e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3802a3f0ce7681b6953e4aba86f1f64ebecee6a5f4500226f7cc8b841c9dfaa4b4a4da8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95c84be65241a5de039298f9bc0fb7a800fd14625f82b496c6750d466e48a44d4ec53879;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1549b0b774d8a70135c527000409b687ca7de73aaf54c8a19137d6be52f47f041fad4e201;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ea4abb1f7dc7fbfb3283da30d38a80faef866161332537801767b8c3a0f85487d10013fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fcdb852f8ad561af905ed7a90495494ad06e312f5f2c3fa8a713c5f270f0fe3e2621b1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca35780f6b2d7cf6d60beb686d35a76c6eb21a160a829625652422b2c5f918716e86815c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a241f2521dc1baca25ed2c032b34949cd29f65f0b948ba6ad7c4c77cacb468824c820dba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da54466e0ce1d7ade7bb4028c794e5e493740a987ac41a22f9940cf01e9fec94f705d5ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd0000586bd06fd4e1a8d43cd6796e327cd5e5a179a606f1d6ae81947b36c2347d9c59a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b526a2b672edf245054316f9b7dc898724e177a259bf99c7a321cec00bf8a1f9277c9d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbcee007efb1694207a6527860dbfcb2a5222f46fa4efe6de005254d9d35f808453bcc02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8452d2d53dfae4ab1aaf1dd588b63dccde8d632774ae8d11f811b1a773cbdc3296a855c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c524f6497688506a5c10a099b87b4c786e5412af603f64baf68c111ee0c4f648d360e14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a828891841e0e93aab32c666973418fe383ba288c22a52857fc6debb117c9dcaf1e43b72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162696c47163ec75e828aeb4791deec4f3e8430182e93831bb5535a3e535d438cfba9ce31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca78db001c9fb64faf30a774d34fc797893b28f48aa546f25200747380e7469e4828e5eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had2963f4c8660f08ca30d6ac173edf8acaf35d4f2c86764cf86f05c5f5c20b50c1c1014a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41dbb34f60f406436635b4d6c2a0c571eec8061271cea2b252abcca3600af4416c75ff67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99fd415baeb17e486e6b3fdee5ebc54d5bec3076a8a581cae326a153b65c110c93d41446;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd0b6a483249723e2300a1cc1bb5e035d60f1ad30264608b8dfa2a82d353aa3f5793157c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3a3744a9fd8d717b5f04bba382706775c3815c45dc9a0b644672b5399bab7900b7e8eda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf940f8d5026e692a695c27e0a94f5f6e636893b58f7f3c93fea2dc383d77b00e87138578;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28069ba64a8a3bffdb918b8a6c3999903e459bd242be48685faf55cf5e4d65db7c48f863;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c782f36929d537fd64dc7f989881422621adb1c4a1d489b81b3c5fab4a09e7e7134cf932;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4f021ccf5f755cbfe708e946520f26b4c35bd15d4a24cb3456ea1fffbe3b7a09734e997;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3950059ad55e3810cc75f0733a91707a684faa1c3102b93c89faa487bc7d0eedc8147aaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc96a22c051e58581c35134ff5dd4fe89072f48d2f4814c241dcabe5fa379c2514888e5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf4cc2ab0dccad96c46099450cbc1b8131a7a110ff3136dc11f11e25c527143c6ff1e77f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58e7a65277824c6712a35c9c3d38785a465edd8964696be8f59958d0076d21088e402ae8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e0cbc01332f5d0174234baf5815f4caf3b63f1311e71c9836b7dd9d994b6278c77cb0eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb29e2706c42f02d958ff0904bd58138d10e3b01663d17d7ea06f67d819921711a7c5949;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51143e020b8c46357fda2bf5f45e67b0f05c58466a2c534dab50943fd35630d0c9e13483;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14aac696e009941cc843d1ed05c3a69c8525bc77e748afd469a020f7bbd0d02d47d56e943;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb2b8b5533e494f2193dc6bde0715989f2ee61257cd25423fd6f4bf6d40bca31afd3300e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78cbe37a263606c4e7f620cce2df376cdf4c9b959622e5d384e8cc1cceb048ac801f00be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cc6feade690d794f9f63c84a546875cc44008a01d2eb0406892788bb674de71a7f731f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce220f4f866a058574fd259bf8b6039fd6b4e78772fd337c5248e2b33372722157443db5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1521e5f2efbc2fce424d2c4583925da7960f4b312a5cb7fa98767261fe814a40132665f26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1690be488c40f51455cf220ff7e2d2c9b0a3e4e1b0b4c0e6f819facf67c027d19a9fdd0c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170980522a1d79321f8c124ca41dbabf68590c4a8f9770de4c2473a574081496e897a92cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h856b2a83c9386d54c3d4c75a59ed428ce7d7f43a1aba52b1e0a9e1bdf6801ad31aaf83c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc46b41a83c32ab68bc0ae6a26d815b6d3c2ba27b5b2b444f673893d4eef62b1894043eae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3dbd27a0bf384d14fdc77d794ec17ba0331834cf0697bc529a39f264d6cd5b4bce7781b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f3d5e5d9957c1a3cc446a258b6eb30927ac8b6d612c1969a2434ba0007baef10461fccb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116c89195decd817b24f5d007741a4b1d1bfda93eab13b05395c5e3672c019d9c8a9a693a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc31050798b7eae5e08b3733c536452bf5e548826b743b5eaf7be81635924a77156dcecd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadfc7c0a8271fcd9be88bfb4995712b9cdd25d3b1e4ece1d88949221e13467f73efbf837;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b65b7e9a997c2cddb03a86bba5d3b44a34ba83b2347be4bcc853a7354d110a7b198f111b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cb0da2a482146939961d1047f0598a3758a4e1f5ac4201f96a852ef6fdf619a2ae32cf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ad5006e346002a774770d090971d2155580e7bf87beceff75e80c0bdcef37d807d67f08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1522184d541153ad5ad5356052166b38276bebd1658a6e6f6d54f03081d491988dd768bf3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14096cb9baf447ab6c5e849bd6296f5d7509abbda4c4b2f6324f792940110b520cbb6cb32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fdb6dd410795c5ff8803fb0374dafad34a6801178d2514ccaf9bd6e300bdef8654bb127;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97911ac9aec6cfef1fd2f34879d4b9ec7db8ee82d45a87d1fe5e150b25322390aecb3e18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154c81f1678b21a09b862ba58e66b1dd73f5a7273a7fab3d0e82932dc2a1933536a25cc8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc5c85981899904cf1aba0fa8b2ce0b7a6dc02b8a5d6de63b69262df3cd7d7f705df21f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3807b410c85fc351ee3682459dbad031f65f7811abbaec7a0dcdcc8b7a8493e5f298a62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2b88bf799abd56230cf9f9463a8e6648abed059fc0d5f8b6382106eb5d7ad1d8561c274;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e2f41f04759d4796275e0d6758222921a4ed190adc9863127adf8b472fe210b42c933bd8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7434f0104c9a018cfd34dcc5c16022e64e00e97fc133dac69abdf23e5292c375d8bfcc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b556cff3a27326f7b69449439d13e09ffb0ad1409abdfbb64105120bb5700a9f38c2445;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1423a3c617bf6a059ff96765e205f2d09bbcb05b577653256afac2be710e2de3060fa9e3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114a94a6af1d4682d52132612cc9363d76182f135e762f41a57ca6ca343361cb1f3de4844;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69db246f697138f4cf514cdb3044609527839506f7f709dd8a5cddd1ea7271a8100de62f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had3128a32961523e09345aedeae21577bf9d5ea12d8a5b57a36939ff95ad27ddff772c02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd55359e6575ab32c07cdc27de92d48b0b08cf9f30308e79593c1262c02d29f651f8f5c70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6618c457efb4644d56c5bdc362bc8860091c83fbdcfdc97e462bb3191ed83bc489fb729;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcaa68c77535276bc5fa9021281d7a20e6ba619c20eed3b5f3c0f6e4379689beea94372c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha009cf963242da889a15a614c118adc092c5db671e61ccf1e6144e72684cb00f5ae8c376;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf77103063041c58ee362f7597a82e6e7f00ca36da9330f5a09fbcd90de1d3d3c4dcb7525;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1408cb6f7f278518eb779344fa42540556e595b09bfc05f2f75ad7c7510fe97ede01d7e52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163b2a1b05a918846908c418de7b92dd0db7ea2002a2fee82bdbda771a9ba70ece5e79a18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0f6418362a39f73b7938d769b24fdd2782057302efff720cf77456fe96e5066d841de32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18493a246250c3f214b7dcbd09ffb7e1296e5f2cc1ae97cc8cc8f5d554ceeb10f30ea57c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1546e69f88c89e02d849a7215844c295ce3e1b9a6815f92a1cae70af39a7bc4c4f52a1ade;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7910ced296a9d9733dd4788feaf12c74e98fd67c7c3fca2988e614573e1d7a84a9a5f5d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf58b6bc1246d35b00105d653a7d6e699899d3e842f6151c80a3d7f5662880a3702f4bbec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5bb26e91d23b46e0706afb0c7cacd7dc666449047213c6c0f9184ab7f6281398d4bda9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc421a13d42a828874d2f148da3f2a819785a6d67be2dcbcc2761f4a5bb8f9106169db18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc15f5ba2b6ed0cea702f1d54eb6eede61fe521c3f67b1a0d75429dfea902d6f205bf63d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd50fee71c3025dab6789f6b4546282ebc8b130d881f6dffb3b1b1ea13823e6d243e1d84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he97f982086dec64995bc561d737a057e722b74d75f0e4918bef92b0cdd3af1fb6fece44d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195a17e7acb3617f897da0aaebe971a2f792012e2e9636c45f2f28426b72374d95fdf02bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd93847d113103afe6b074a73f93100f302230655b236541994046ee3285348abe836437;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he0b60c336578a0dbafbb82a1b8f53226d81edd6c45363d3eec71751cfc022e0500412e80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf95c0f82116baf4f12cbe8deb0364e1d06404527473bdcb59a7ac3e93ee94270497b84bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9dea88c9ab27523f3ffcd6d4ade1567f8f65a6d4f8000d37f1e6695fc6b61afbe9e56855;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74c55b143fffc1830f6b95f29b6b280e71c1bee768ab3481c4eb3746496cb1bee7e99f99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b64968f8afa1745e45f53a97b9cfd59cc3772fcfaf8796d255a1799b813a4343853f65e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h851eff6467dae11637ee814b0ea856743b8336d7b5a6f47fdf5500f494fa6c1082aedcd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3c51e69f5537c75dcb2bffbb5d0b8cb1237abef0e116768a9bd5d1847fdd3b7f6b3811c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he62f88b21f6c552ba0a8ff8b40812a6063f7a6a61010c7aa2746f91c119618fcc3c37297;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha74bb4c28fc070f6d37d7f8d5df42c5ad856839d1936e87bdfd1162323324cd784829a86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fb427d1ce858df739e67e481b21ea020a5feecb8fa2be8ae1ebb5ede4ce6b5b60a3d2f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3131ba60164cefd16a41f62f416c800318ee67e74d9282736b2e6bef72ebb6ab6435b55c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h411981f1f771f465cbeb1bc422114c3f95cb049f16051bfb70817a8b9c1e2809f2f61e22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19afd9c15022de3210159443e2a83d34dea7d55153eae4e6b73bdd8b4b9608aa48afc20cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha99eeaecd319b0ac212397dd91440b20ead7a3a3c5c5345e912c4f4d5ee9cbc0dc8d6592;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e5b6ea6b325aacdd1172c85bd6b33ff1084c2ebe645870f7df87d8ebd57f00128bbca5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h470c5b73d0128991770ca3371561bd408edb8b58e39bafb0bad470d94b07401961083d29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had5fa4fc5f41681e63aeb3c8e0a0439208e649f7d8201de807e66adae1aca4a4b6077c36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db38f2c70f78081ff93191536546dac656f869f60f26c83d5b527f049766f41f1ae13652;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf32991964cbbe6749b7c95708c7858d64bff558292f3264657c1933c1ead7fcff54fa55d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3d35070f906397bdaae97b3f00bc8f2a02547777f182b402fa904c68c534c26452c1a2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1088fc8bafff1339c6b746cff7131708f444a0c07740f20bde417cbc0cc464a3c1135cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d784bcb2bab7f3b8b1a97d1cb6bfdeb7e41e8f8fcce145710df2eec3e52d9778572f25a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he551652258af42be209a48d7f126b37955241e7348fff091f1336302fdf71ed9a40cb3e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda86dfadcd8b2a7027d2c157e23615532840b97cc850b14fd76a3b2906ba9248272d2a7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6389c6e024815ac70a76d82506ca0bf7a61c6a90dee5e8da0976a840480566df387fac18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef716c9f76204db8c5616ebf3fb45a296488a14af2b8269f92a437fccf0eddd65a32d48d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1767638a7e2cfa1f837cf5934660bd07880c2da8594844a17e896ae3c04cf21bdfb5dbc48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18578e1e556658802addbca7c04eb81a70adc02bfec43332460957a9745d8cf976880703;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55d035782cd28f4f41064a7e46efae7712d58acfc9799becb360ad4e9a27f507d0888d22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0eb0e48df38d50df9c79bd3fdb898cb212adb10175d376544b464445b13d48379e3dd4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d442f47f52061317cfdaec04f39e536a0a1623739422fb4c154a08088a9490c9c1cc0fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6057ff6dde1c33a0829a51fdf14a986268dcb2dffc69a6b38d96f6200e894c8a144074d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a7d20248a71ba5d75411a11ee29380fa4b3b26cea5a4e2bf062c85f1b7c1060160f53e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19be87f8f92fb30a4df5bbf0e0ce3ce389311eb367357b32248bb1f7049be6af12b9b5e7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf7308c092d11396c505496cb6a33ebd9a568751a74dcad68a4049b26642c8a764e4131d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb294c1e8bf4233c65a77291b933711af680b1d02daeb6976a73ed42095429da07cde72b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bfb8e472e28421cab45afbbba400623f3a3e957420fe4f7fb52482a59eb2440a6f8c9b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122f31374a496825f8963112960ccced98c61d7449db0c5dcc11cfbef4c29c6c32433a461;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e4b3f36749e59d9b4e9f51fa3495ecba9c6ee76f233c71b6464d8f5f73977033e5adda6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115743612828ef9fd613c1406ab4eacce38c233b652ef29ead0c8e3f30114a77fdabc4cc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb68ce8d3e1582b29e06a51fd965834fbcf9dbbb11faba1730d0410db447040ab68a1486d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36874c4c8451f91523145ea8b126a9ca302f91b3d2cb75ff65581d3cf9340fdbf189df90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd272c0ca6c937823397189554d5b7a0c98e4481d4181396801384ff731259bea87138a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1008d4ae73ae32fffef50c15c974d8301606093f2a36a494189f1d9f16dcb507259b66222;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6652bca211af8db87220850bf03e148227d537b50290dbe924498a3c5fe1b3dd94523cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17dfa7f5c90d8ea78654a51ffcc5bfd85c9593e33f6c64f930f98fcb4da09ba84ab2672fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1846a19ebbd5a73c2851ddfef100c797396514b2b014aa3db9deefd0c624911f9a2003de0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18512d6e88fa6afb282143a5d3178a9795c68747f6ff36355e0ec21b025bcbc5566e33779;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1365e4e4a1915a3417ed778a4b682005e732eff94a228a4c7d77b1937b3c0c34cb6b9f72e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9418d7c4a3ef51ebd34f56ee2a28410b037f40c8203ceb285e4cb7695c85a8320450c59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1056e6c0235169000202c21df175377eede507ad11def70d3ee327e0cee2c38829593ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e28aaf6d1b442405d8279f4ea6c8d05dc4fa071a2eb240d250aba40ed87d0d6c2dd89dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d9d1cf095ce81ea718d65d5bcbaf5ec974c1156dba5234b6202c1d0a159d41c02570975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e911b5eef7e99702f6fe1062cf3f7b932078b87962aecd4ac95c5e31fee6c9a074e92af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha56428aefe89ff18afca8a3028984c19e91763bc978c636378ad3f5651e5ceefd9301bd3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf077bd0616cc507c11fd6139da7384a1479e75ac817988501b33c0126baca45921aaa78f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fadf4fcda1773455d6f33221e3e4765d989597c7cc3449abdd255c76649d88475992394;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91b0bfc7593298a5b5ed09db5955e4bf3c6a98962610b1da1ff64b7510186a021070b6db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h983d943082b3452c3037913f1eb923334a35eca56716e2113b694659ff353fdf12a85893;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12eecf5bbad69d2ccbcbb43f2061f44eec19da3279ebba6ca1d271cf2ea17076ce7c3397e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e60d8d62b2be8591c025af55da77bbf787d85dbf2e070af0bbaa9f47b2513d41bd35ac8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e27ae20b6fbf85e58f7cadd754fe840a7d1536ca2793965b5d101d4aa97fe75f0f40f62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15adbbd55442aca9f9bafd623774569a5e68a4eed255bc253638cd69a83c89b11b23bee9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2bd50661f9d584a0dddb9a1d04e90278e2e7ca8c112b9fe0da2bbb2adc2eea21c181278;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1366fbbc463af5280af8fa9813876bd7cc9683172fa4231c2d8ec2e09bb97b906ab886311;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1100e6938bd6ae15ee102cf5d85babbc51003ffa3fb5b46604dcbe0fcf4137718d360d51a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c51abf7e86916b251b0344a368ae1bcdb6cf5e9afc2dbb3c6c5b77d9b99c3ea58cf69f4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h231af053992b395a7b5836655a0dea8983087056f18455351176bb8ad02b32c9ad625386;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126b355ce908163705cea40d1256a643b9295fb8e7d0ccf459039c34442a8e121bed3a016;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf53bbe0b1bb94c1192867e68ddb188870db7dc49849513e1b846f5de26dbeccb1165bec6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b02559feba54c8466dbd8bf96afae5a7e2bb4278e529ba79e1b3c0be7431744bd8e9138f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195722a6c71de32406842bac9c1b6fe81b97e1ab1b75eff94c6d87bf69cbc5376e1540986;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1b072408e95e4c5471e76978c3a46780b16adcfd6efbe2071049e2570ddd151d0e618b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae939246dfba57269345e1b70f5c6582c9834f82bce0abe84917200f87ab65ca6b887f66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4b098db87342596420c1a8b67a2610ae7f20daac60de2b621abadb93ea30142421ee833;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfae1934d7395151b08d4c83b30518e6ec62ded31580fc4e0daf51f6c0d00c88e8c47c43d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1845fc69874d508a37605dd846f2332b77387cbab17a6f04788c868a09a66495856f38c69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98218d9566fe45f69f7829e1305ea61b6d1601f4f78efb1d615f656d93ed0aea06bd4385;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1881e3c8b162e8f9511dc21cb5c686a75c431a8ad80e88934a77ad7ef5d6955fcdc254986;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bd6203c75ff98fb054934104c3daa87a1534d455de72063badc0d13910f1758726d634c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1002746732d8c3e5eb2ed8fe4ed51faa163eec26d578af3b0d45d14374111e3fae659c604;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3c54901c06cea1201055ba300278a3d78962e357278809f2c4c3b49150eda500e910da1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21edea9df50c5b9c57f82b47e6f4b15f21ed1bc7417f1de2ab46df84ed4a8671cd703c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f8715d9af04df52a718abc01a2c0bfa04c9845a4cd084bd144bbdaa1c201fb30cb84307;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15586d87d679aeb4dc674ae6245bbc915f7ecb1c471afc01fc2602470826851ab7fd5fa3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11af606e59fa2e553108c7fc980b3b84695a47cabf1ae3cfcb097ab085fbdd151d30e3286;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a43a2d8670bea92d4e1b1e79b86f48cf68bf353acee28f9e304a524673bb401b26898981;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1501e3bfe5058ce3fc3b6c6e74da94629562c873ce5b8c66221112c0765fffd754a814be8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76a480001bdbafdae76b77bcbc80192b8a1df7ab535df4745f8a4e5f34657c545f982c94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112e56b813ee5b22b17e7d63bc86b304675d40c6637b040223a3dd9b70132561d609b3273;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1901718a33b83e897859963f6cbf43825681883e5a3ccac882caae80c4362773ca0c0b848;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb5d9902998081c0d1130f9182c1b3b8f838080d3975a47b4558e0b51323836eb5f8641a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h382e02445d1903e0e856624fec20cea486822e364f9f8601838b0f0a8b411c14b4899bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h535aa3a35d87e30c35a68347aa25b44fdece3bdc7eb707205c9689bb4f7965f46fdfc3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha17a599e19f38200114a18188dfd2157da85a060fe4ec96b25c53760b01ded0f0e7c7adc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e305a8989aa3e94847495c062c618707ba14f6210a1d2b2da922971fec2c456e7c40ab9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ba5c3f19bb7b95ab2cb5360c45a6f74ab07e899e805464fc59483f52175c9a7e6ff186c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h612d9fd0bbe285f27f380fdfd0c2609945778272515b20618592235cd6fe7e5c1a207773;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e366e57236967e0517d242cf1656e9d996f4bd44e0030a909870b78e85d52876bd438cb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25b77e692cae520b2022ce2681d513ea38874e1b3f3309ae91d55a67a5b4623101af09e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77e774a2ec1789a9ced164f526648ca1f0c2d3b99844382ab2e83baa017c34bdbd1ed4ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h662eb0ea567a0d0d05c5db2ea04942b333a06f714a33151819acf643ba500667e46e13d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h167b65c7f5fa914ee0e9ba00520c4f49b678457ba5db043ecc91bcf36f94eaefcda8529e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16570d837fe3e3fb067e89081c242eee96379fd5b41fe55e15b4ac8bc1eb621afa4109675;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fd07f00d6050040e52fa78f6fe2cbb0a9996985d46904e777d44e2bb8c3f05c7781b1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132b6cbcf0b5fbde50863da38d92a37000d7b0d59db324646d9a0acff0f493f6841fc864b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16af06035719595f5962d3b1180f9218e7574968da0ce383ec12626948712e4a75b54893f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b0a3f09d1bed982125fd2dc3c2e069074ea20579c5f2359cb6bf4242f643ca9db5be0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f26c333663f221cd975df1c0f26c0ca508c5efc1f7f1f32eedc1c5f9471ee5a60a44d9ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f1db9fb12aa3d97b9bda7c38c0659dc59f40e4b92dfac9925478d446d5b8501e65d9c37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hffeb50427023ba6603b6caa03267189560dabe7f624de0e52d5ba855cb181c5261038ea9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd58655da5bd4c5e78a15fe84fcb5fbc0af665c5231a829a101e2de71ca15b7ff6cd63fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bad54358e785e046136ee84246a7885a5f070e8ab124f20e21ad31c758e7f8bc54ed6c26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4775518f8c9b82f786328eaa7d4769427dfd1348c744bf9653cc8bb4306a930a416c71a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1a1383fb2b4dcbafdbfb6dd0cf22c67844a5d97c8a13adc11a90f3f4067a88521a52d7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14dcb6618d96d18fb30580c5385ed9fa12745fe745ca96ed8973ba8041615ab03399efdbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf964f3ebd702dffaaccb67ead307e1a982b6eba167e4b93c0429e6aefb9b863b0150e7fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c818f05c7c331983a711fd195c113c4c4eb2411891e3b5ccf530e70e948fbd82199e5c73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6d9949610ce57e599fca336204ce8a384f23494982600633bfcec47ee533ba48de1e4c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c0fa1fe1f40ebba3fae5e112c5ba5796305d5f150359504af0d9f06346dfa1d1423de66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22ef473dd0d91611a73bbc466900c9c0cc62110722ac093245dba102f73da02b53395d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a61d57158dbeb83bb477a23155a6215642ec27504c0e43cccf262702ad0c1d43b8ea6033;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a711e38f6507c230697f934d7d01ade3fdcce38ee31cc75c877915f357d9e1fbefd5abcb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e2c6ec636ee0f441868ab48a6765474e3663003aa8cf90fda9add394e085b04a098dc7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1313565e65b57f43b131bcfd5991b54a47dea935a31fabb2756786e1cf0ad46bddcfa959;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c580cd0201f3fdfa0eea8da54db90a44ed085a24ae257eb2fde6623fdf574878de9b8cc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abf0c29c6f61c4cc082be24d6a1382bd0053d76a955872f0622b7e185e7b8d8d801a2fad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e00bb89aed6d5dadad2e5675d66ed4a4afffe97831c43765af213c4df109388c36603f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fae07e3712314a8cdd088f7da80401b353a2f069bb830370dfb08034b2273e82d4fbc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3b21f3062e6ed6547d5812d3b3133deefc9624d67f3c1f38f6c3bac8636916b2d1d4e8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1941957b6fa1dbeab5dce70d470b64c765b12ad2141ea5131e8485399cc8d4f16b5ca6ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bfdb82c99a09689491006adbeac817eeefd7876500811e57794f14757520bdfc99724a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h861c7b3e6f23f06e8b4fd40e3cc20a69aaa020eed77369a12cf18d5a05cc1c8d7e89e911;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f6b0ffcf528542ad86bc208e6d6b3608760cfdfffd4921260285ff783a0d28ea7f8bc47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9710b795598ceee76028abec25d6cda6ba26f9a477545e7e56e65cd8b0cc9e623f0ec53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc2ab41f9619b66eb128be8b914c7dc5dbb4cbd21f9a2e55e57ce5ebfdbeff7df1727e61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6568b7f1f8a0091aee6b51f03c4cc2d69c173f154d8f2f6c81ee056cdc20c2e4ddd9cc25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha60ea1526b330fdec061ad926c3dfb676e3ac7112ba265fae0bb66f915f8b06b90fa2e4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf590063b1eb5de314689b8f3d51d396419d7c43f318420124fdc72ee3c72f309b53b463;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a097150d5e51c514dc6375036fbd14f1a04dec9988902ba770f2114237858db8c900c2dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119d2764427ee13801618eeecc6b80ff7a018516184f7a98470bb175aadd25160b25d251d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd866a97e49f04a212335be7b6ff34f159676cec78ae79f4d49382bc777d40adc9703585e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he96fdb1370ab3d98520ad6364621e652ff0544d64d369d556f6cb0b50d63e842d231e23a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf96aab85379fe47902418b84645d3547ddb5ca23210159cd27a72f4391c9d27295a0a13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9c771e202df3a1f0311e613474ceafaab0d29ecb1626061fba22317d89a8235a4f2ae03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf779ec9ccf95447c4284d85c6df9b4119bcb3b56f0a9c670cb3d324ac54c32d0843676e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32bc8072bfef0d5919d8e0a7ff924e6b6558d937f46d2b20d6591b4a48e35e6af6e6b246;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f91e42c3c9b3a9afb55a3ce271fb387873809928f4832feb7bb6c0338acec52ded5e184;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f294a0ef92b30445069334c62e8b67db88a2a0f1bb70c2359ed9dbe456da1569a88dfc9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e061f64a22f28c3eb3d5e7387ead5f9c1fc9fb50395dfde871f49769b66f9d7d28107fdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f61545b6d7b87569faa56ea0e94633736a3be52debdfea437b803c2b11e25e1a43c3054;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1deba0c5d202f9a611f5b636bd7f8a59e5316864eefba95c1527ec359708115d9faf0944;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d91b0ed292f4b0886a12d77d893ef30b024a9f9e86597aadd9e01f0834b34b9b6a6e3362;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23d0672777abd55beb14809bf99cf7597fcfbe9103739af5a6fa32d5cb2129981a9ba529;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f26d9e73dbba16b6ee34adbf547e7f078601377a304604a17097d8e156f97c5820b00a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1129a3abbb3aeff6d0856f2e13662af82a6e3af3aac47e86223a898c139b77296bde79799;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158652f3eb8ec6fd6a9fe70d1901c0e33a9212663b1505633d6628157b1f7561715246375;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173dcf6b4691bea6155d79ed553bb8aac95f25c650df966570f70db3550dfe054b7b0afbb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ab5ca9b2ec98436be7ea39b390160268099bd7a77b467053a564b431896c7593b058330;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9a871c4071a2ddb26a5b0e081ce60d8aabba2bb39714f35aabd73e333dd9dce8e0202d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbf5e32301e1c15d948a235b5055431ece53a0da9ff80b36b41e7adff73e5fc6b478805;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd1b7750fade7d5906a6c966aa1799b4012628fb9dd35158eac6dc46cc2f951fc5014fad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e2e88827d87b922f00a146407fd53df4facf199e2326a13985b7914320d61fb8925838e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffab4aed0f6299560c85a6ccac9b4d63d1105afdd1306316c1e95772b7813e6ec65f96e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbe3526fde478447e94ce05da89a71ed8881b4261902e293e5f688e7a3440f844089748e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h645fe83297f0f1cfd531096b91b9bfbaa69402c64c92a762bd5d01c05868d8aac6f7d73b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2a4d098938dafbec13020370b93cd87cdee3a0a519580b94f6209ed1e7cc5b353ae66aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41b60648f7dfa4740854df226bf5e4ba54b54b1da1c9d1b36fe2ad18f38995073643eb98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b016b98ec8ef5d5e946a85e4b318584f763b4482f963384cb7c2dd235aaadcd67244cd90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67e3d32cbd4fc8f90c4f08f61b1bfa8449c7ecbf602c82797db1aba8f55ae01d419220ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c8e285fff10e7e77ae1bcfb9c9bcc57212acdf0f7ad35b362383cf4fc127ac26a6a49b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee5a15776a98a08e0a5357d3005c71e20a21b57bfa3e278bbd64171867348e529e045c0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1914e565e71fca4850aa682bd008cafe27e57d538d3322e3b0d05802d212f0e1efc69d1ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4758263a5bc8c46c19558bbf79b85dfb4baa4978314db60bf3cded6e1d744d08fccf4975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c2f6a3502047f6c9c60688047cd76bd6867f68418b9a8f16fb8a89f7de1d82da348058b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e704929092894535767f2b6f48cae36cc4ff10b36185486393cd12c743d1db15cbe69e6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce4488ba2d222179cb31272271db9a74f857588f878d07fb04dc6c06bf9f35935f478a6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2d08b0bc4fe8ea089bae96d44c804b527601ab0ad76fc7e44019dfcf320b3de07922ce9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16bb5086a3b703b9cfaa3957bb8aee57038a81e9bb4fa9c1e7a3043cf17c14740610f64fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h650de834987ac38e96e2cd6f2a32a0109f046555798ea82f429286ce4cb488e559d2012f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177ae0175af7639f18ba814d13f928f5cfe0cd873381656ef112880dceff3966570608718;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd23bbcb7048ae38c417becd759eb6ce7f70caa6cb56f4b5eac55172e08574fd3941122be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aeb60aff3699cf4fa19faa67891656ae26ad06ae077dd431bbf8dc55ad821a7a8f018faf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0866dcc2fdcdabe17b0f109d93d65c46bf1dd509242cd0d0ba93e98732e6a8e5a44bbc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1129d3fec2551645e9b414a74ce83b67e778de369ec97bb9e4a59945c33dc4a996b5d24ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a843392bb989499cb12460cae231932bfcda39d39bfbafb5775ad69e585a874407c4c3c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h972e27f2bfe2cfd5bb7577d1da57373dd5c2805b74d88f6aa862fdcaa20857229862ba87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1343b83b258031ac053157dfd0cb22a025a51f77396f06b712685b2f3a3fa4e26c618ac4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109ca0055bd0a0986e41efd03794d5a16bb07fe2fef07eb73655bc4b80b2b0215b5150d41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110042cf9814f4f90e4108b9d687829ff4f970dcde601c590211f6a68d6a9732a9d55adb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d615b0039e7ff41e8f8649d4d72d8d7ab7957b02288620336a0a7298915a1be36434dfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdf0cf4ec9266bf5f4effa894d7b56b20b8e0a1d21b8ec4cbfcfe8267dbb9f772009bdb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c75a1128407ea456366f15e3481a21cdab301e68dd5fb8a1affd7ef8cad46cd46ea47125;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12209cefb1de52b1dc5076cf263ee057db77f7ddb4fd2d0a8bac66a944b98e7baf98389fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he49e15d1a5376d06103e14ebeabf606523c77ca7bc4f92b11b48d0f415918b9e00e08c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fbd1da9344cbb0272a15f30803e39f6c0b0c665fb7d915d0fdd166984808eac61e9af63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ee9165213cfe9d6c92a4a698a2ee4c5ee46eef31589456ab13cbb588401047e4dfb891b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1802591ae135b8632beae8d9dd99fc14d0e725eee79b59b48520ee0f28c4c07ea7944cad4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0d7e7facd024ed242c51441e597aa8de62eff97432332c0a696bef4e0da1fc3f02260bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdda98e950752797625fa93a7a5aeb873c832f0b87e12a5dd1f2940673a1588e7b0570251;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2755f46bbea0317b434984dfcfa8dd65e159e7c062539ff0056163135d6f1a8647df6e80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129c047e6e51243c42d263bbdd7c006fbc584b73c9a3e949693ca7e8316b84da1a991b934;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1642d6dbc236ff049193d948d907c5d3220ca804a20c9fd0630f8653922a0a6b09f180536;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f0772560deb6f5235e5929bd40d5b3b6a41deabf53a3c426fa9a5e71967fa32b92045a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c7b068b8c47fac6aa152409d42dcbae4b8fb5e367e3b2b026cf80a84b637423d184bfcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59440f4602c3dced993038d1c3158e3bfd72bed4a8f59bffbdc47ca7163c7c78ad58d4d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14434897e4757b4acf07ee0cd53784221c0eb0ee3124afc5521b4b5a1f960b03edc3b8526;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10186b2796aefea23ee88355edc8f9dd5a817b99d364084976345afe58682459aff972a19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17672288b62da6cb16d50b83825685a4d791c68e10c883b43413f16f46111f1704f27e03e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118d634041f8344a8c063c715073c491444a5a5b44df7dc66c002818392aa2700c17128b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114109be452b792af28681513e47b90e96ab9de771989a6450e127eeb932720c00baa5b57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19264c3dbd343d95bb2bed61078df6605894491b1abe05754b45caad32d90605c60cc5c2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d3a743d3995edcc1888ff58653965216788d91892362ec3c4e1d78b23c6872c0366cb73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h820e0b5a141431a0d923e4c16d6fd64546f98fad06dc78ab58128b194cd9868a3bdf45d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2fb5a0ccf2ab3b7eb836ec21d752067c6b6e5856f7beacd90c8516360a5bb51a7fc336d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7144cafaec9a43f64fe2e8bf29a72d6260e6784cdef0b03c1f884334be662cb081440d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd6d3ea792d556cae945f2d26b29b5af3ff159c547fc703515e73df0bf23bc6af1e8d5ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a72dc095a1a8e38c99ba80a6073d2f36dd5bfd0e3b7ec34c8eaa76f8f240bf532f3e93c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h794166542ff3d59ec23a46d8203af85ef4bea4ba913ed9357c26a14c338a2c9a02450e6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h892da100f6438428f5e258f74d931a3fc0b63ea0a9a4346be144d321d976f481b53197b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18203f1b2407d28488915d3c8ee591aed0dec60402b6cb55ca59eb07d1d92dfd03b2e339b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ee1f74b457f6af61d299ae80a4b2ca87f8c6fdfd310c759eca90bae7dfba6abf711cf5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3fe0211c7ddde894e6197c8037ad0053359f74c5af2e50e88f6a1dac4320f3438bd290c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce58bc5d030ff03ee830ac85fb2862e4d4e5ce7b5558f7ab7fd9b162dd67737b85e50f2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a9e43f54771d5748c01d9d1cd4e5840373cf952188edd0243f4a1638be0f3832ce8eef7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8be7d5e6d24abb4bf7bbeb8e6ac9a45a73086dd36d7164a7e478b6c993ab35b88abd0eab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1b80e9718c8c283cada7e7705a0871537e4678342adc284ce63258b9649c58c089339a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c41bf369873f9eb1118fced96e233f3ebb8dbfa40f08bac755012cc87c35ca42acbcf468;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1928e8c00b83893b27e69735b120bab4b058c0e6cd71731526e8105a702f4cb484d8b88ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fa33bcb2e1091b8511259f89ace02dcbe054591698453b7c43c96a6e8b9b178efca7fa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf25e5ff2e366261e37c4623a227e5a0c7bb28cb74a800d131721853ae6dc8b381afd169a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b8dacdd4cb24094817c06cf5d20d05d66ac3cb1b8946293e6d55d24621e40524ad3099c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15541aa12a4eea3d2e88935ad84b6b2a71ee0a744b5029ce8076abd06012d3f93c58a8226;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d96030c4c9dfae847cee520818d8110b4fdae92ce2f13e0314fed8888c554a3b284c62f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d35979c1dad34c315a2b68e217c3acd76c0ad540bc6e757bc5521be3311f23bfbc734354;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f39fd3e99bb1d0b3373085a1a49873efdaac4b91d9d4d78d35a2b187bd23183a6cefa4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb64d56ff2c31b1547cab9239f12cccc6177616769f6b1f279797c4af4d4e3f403c26c04f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ff927a7255f73869466449425ae21868f531975f24435d00e55de8eb22742d954a1611a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h253a7f0044b7eae39401c799a42b22d9a416ad5db90233361219a7c3303bf2fb3ea7556d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10961cbca4ebbbdd9e4c51077580de422329075880220a5fa7a1ed10ed648a7dc5bde96ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a77481cb9305770bf297b49dfbb3c7d1df02291c2e8b85380072bb3831eeb032337ccb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70539e80a0b61c8e14fc23aa19fac23d4dc888c17ce90ca96bc722fc192fedd37f40b93d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0277d0792d64598ed14bbefbf4666d736f1479ce574e6d4d004b816950e7f92ab1e72a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a665f52d833493d229b0cbb7734a349858890c1fa3960c501d42c846433c155bba831c1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2a5fc4c41e8b29979118e19a0b3a668721ea85cad44b287ce5a04d7a8087b324b3a78bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ea1c931a05d8924d0d11d2fa9227f5b19cb5106d58bab4bd6f1e30266bccd7c69e174df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe67d572c6be6b30a4ce3c0d36fe14f11a5eebeb5b9dab9fbe7cd5644712769a43b1302b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefe79c9a5746fad7a927fdd4dc5acb5cdc235335135c83d9e9e4a718c4349307e86c0b04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h92333c7116e10e6a0ea4a709516fa34cdbade933bbb9d3da51a183dc1c692da54bd215e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d3ee3215094863e0d881ba097b8c209e55031aa70c774dd8d12dd89e16c50e7136a3dc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1a7ab2182fe496a9f48440655206cd338c2a2ed891c2f24cb9bc84ccc53e21ed893f9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6074e9fb71ba6dbd3ec9d4d62c72afacbfcb33c61dec231a7c1647f534ad58ca897954d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d4e464ef32050ffe3aade1f9ee9b8a26df7a447a951580186c2f69ff09ca272819344bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e9fb8c15a0cc7921556b7a7adee8274994842cb6044d5fc82704a421c822df6bccc17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7afd6f7af8ada2f87483fa4b93bfdd7a06631673f20b25b86c1da47bea1504506891c18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31f94b6690dcf51f06a71a249117d59597da9c27caa1dadb8f830eca177e636e5184bbfc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1856ad7401f1e1782a03597e8c95fd6b2b101b7f4b1ef5baccef2d0a84038208422745270;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ba0203e7973f4ca48cacfaac62117fdbad4a7bc6c8914111da05e596a9d2902000a12a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12942528f036c610f5d1ac3e4c90ec7ee7563dc17bfc454880500a01f1f83aed81f83c9b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb223222e5b71c6ec1044513b1c4a3ba74f91efe6b8bd629ccb5d75ece3acd9d53f6689a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h815029a6ea18360a246662dfa86dbcdf72022561193c43f2e15068121624d1e0985b6099;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109ccc7266e13bc5de828ce65c8985523b8450e38a7c4feec814bb48084f97f7b8de34908;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h554c1401810c8a3fefb4010ffd08b3c78e15c99b24eba3d41d8007b91277a0e93cbf7168;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h204a1327d48c7a98fece4dbacf68ec1f0c30233d407ae9b3023ab77cfc8c28854df0f560;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49e242cf2f3095f832a0440c28c9a7554f2dc3bbe9efd50ea9c21816294f686d82a55188;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80fe8800653e559ef18f3248b4f4c0ad8624d424ef4515a6ac8424e574d9d224f9586f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183ca4571fd6f78c7fa6b6df4d4c0e0baac479f35c8eb6063cfeb5832829ced8d87032fc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9de3e3049d1e2b1f099d42d18773212c8dbe028ee365b711b89d5be3ddacadcbe0c58ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc96212a3f8ed2f74f3403af22aabd18de006392a1cb2e05b6b83ceb78c53904fb4864181;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc723a1a0ebf2211b8220047d4a865560bcf771f0a4adbf7fcbee4a9915af07d73dcc787;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd7bbcc57665d1f32ad569fa5f15aca3291e3a1697798c33ac6f8779bd8630cd01dd0026;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10104afdd3247f18279ef918ee352bfae84b64d9297bf867dbb1fdd4d8b927597bbe55449;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5164ce73aea809eb43bfb47064d51602a2d5c79cec9303936f08dce048f56ef11e088eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c4bc15276eaa35d0f500b1f06ceee551bcb74d120d31b7024e1e0977bdd3e7b5cd8e79f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e5790d211579620a2b5354bd60aae157aec9af9913a33970bf53f7e9fb8ad7c8696af03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0f43fd7c283d2936de2776f0b0171055670bf6b155438a3c7dcd907141927b0f2ab3a68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a33ffd1f08ca7741471d681a787afa9eb87c2dd17b02159941508f4fc26a4e32efd5281;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52adea45d67e0e8ca07482cf0e0d9b607ab2958c983bad5130f70e733f28092b58063569;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h435564c4ffb0c80022a05b8043e8e6729ca2093c5decdbd7db4ee637fb8245c204c93d01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h942a431a4db8f121b2ec84e0f9aad99998288579af8b582f37599459e065c1f32c34428f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4f29ffd29d991734eea1a9fe7c3e408d23305f78a27e8fef386fd1433e20c14c1cb073c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1096413d51298bb57a4d3151e7e2726b6bfceba34c739adb0b7128fada31ab5329c0aade8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78dfa435b351852b506e8f9fe283f36a1690fb1f38bd925ba5b68432bf4ed9d56562c1f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12655c175adcc3e2fa3fae8ecb304d7bd71b764a8e574a55721a93275fe542fe3e3c3689d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc20e03baafdacb185a115ddcfdfdeeb5c7e43a9e602f68cff4e895a1bd9d83655488e3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bb80a231934a055225ff1d62d046dc5d6a44a50aebc027f230a80b53d93b9e345fbf37a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1b4c8b4783ab6bd954190e7d922617a8cec119abf4f42d4825179e1e5a6395a69d5cba8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7196f48a94ec07574798b2a8e64a577a143a1e435fcd5c636370bfe7a440ecf69140742c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec9590495e0367098ae556a3b47432d9c33dc454b41672e113aed136059db9ea39c9d111;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h794a51d3fc7f15db950c8ae7a504d6d405d76e4d0fbbb256c34162dbf33c4f039cfb3208;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfce6c31e9b9fe502fdcd3bd93c88dbf461bced6b1eafa5f3dcfc7899076bec19f1011e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c27b4093c5c4aa19c4fa0a4fc75036e765e1b5c9f7d09b7cbc300e3984b0d9e76e285ac2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a707b9ef0e3e747bb630a7732ae484042b1f278d301067c6189dc86b33445a0ddaf80bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d0037a74280211bc562e79be05f27b4605b4757afcd56b41543696b98cadf97d842376d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89dfbc17ccb0baa066580fcb2116420627d393766d0d6a4de9ad604f55c7542c2af57ee2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15adfc8224f64621fd5ad5ed394fed1d6a895dde24262457afb7e78738353c1f1d1ad4533;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152a4ac1b46b659b7fafd213172683874d99246ef56a62f90b4fe59b7007fc26c9167de0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14264f51bcda9d60ae7a35ba799e3e25b21cc15c4aa75b7a339b9ea523cb2254b8cab4132;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h256fb61771c2d95f1d5fc8e63d3476bf62b66f7280bb65c3ddb6eca80744975821059c9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3968c1f9a45d7f30249a1669a05fe9368a4c79f615bb334d6c0b8b6be18e513197eb9da0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103d0815627cf9efc6e39b82007675598fbc916cbae87ea5903aa5f6e55b8a96bd5d7b82b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7dcfc08e7f0285a5fb4a8e2a455831d9c67a776c41a79c81b1f1638fab9a414384cf1b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5afff042b2d7606c72677486eaf97f9d0baa854381e5918d3ceb68600b9fd6de53e3ed7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ea513dfaaaad8e3ce227118567bef7ee9f511b6cedc19e8506e2ba53f61d27d0845d23c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12500c2e6f694f2a3ca3cb12e68a61ee494149b36e7221ce76e075806881cb5c82b1befaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a07db1248cc520c9f16871c6f7f54e005ebd229275f1d71eafb08d602538ebc3345c1b77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d5f079c739b4906698f0bcb4b892fb0c44b9057b07333b3b6c86d9d4ad082d6a052fb3f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff732edbf635744b104badce263316806fcf07ca0623cba61f7336cfeaa9abb374d9ef0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc31d41826a1eb74981147a9ec72cf2b0b1c03f958efb4eeafb53710cfdf0ff59bf3c66aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3292d92543485270e9517bca8c018e4b1e4c3df019a395422ee0bd100fc13bca0e440625;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de236254bc6fdd0ebf110e88fe3d42b77a48474297897e0fbb1169d97728f2003b89bfaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fb8c2235a4c450cba1be612f04288e0772d58f3c206355eec09b0e38499e86051d4987e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e342e7ce7c35f38a3dfb7fa7f016ae08c5dfc090568a79d3e1fc750a10eb13a0f5ba6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fb180d001287524bd7745be468f53071fb200f756ea4eb47e6df58aa44678a7b302302f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5dc363f2a80337977606ae1eaf349fa2054583ff9b097b9ad02c84ca9403561a5a57d3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d41fe5fc81efc95650d5db9194991fb1ba7fe53019341a0a7c7d1831d8ff2a7f3091d4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf5b12b09b52113c77ec657b357a789c8fe201a4c96bf0a07a93e51cbb9ce9a8df520691;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5122a3eb0ab42216422cf3fe6aba19b238c3e084d6e503838ae1b79c00779f8b9a31bbe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6b1eeca692fc51ad81d4d0ab84f6f6faaece50cb376bab02ca64dab2d023744e7857964;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f06246c5f7d87b60086eecd251e40d8bb6d7b6943d1c64cfbe3a1c30248ee3c0bd9771b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfeeb5889146576cd5366375773b720f730f32010306722ea9784208bbf095ed930976d71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6147aa8db3e874199198ef52fcb1e46ffa58fbf6223d9b36affedbf24a7df7f8095bd07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9095cdc9c8a0c077de964f569b8d03b356d6195859a4a79fbb7af2244c78c66943561548;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bf842e2d0e43ada19bb0627c7efaa03c211c46bd82d518f35cbb2f080b82aa5fc05ad38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111c8145c46c6ec0f84171b8a7bc6e119b765fbbe807b4676ff14ee38fbcfdfddb761ab4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h816a619c9951c85e3eda717632d6ef499b01ed8855cf74459355a0f3383a2cb6441d65f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b593d2db06784417aec0ca6cbaf3765ea4f0227880443211aea3f8a8c4a88d7a8b5f8acd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c08e49cc3890a55af6983a8740f838bfe13e7cdc031bd75b599cd09e438c62b554f3b6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a868820c64a4f2744196cb4585db54ea32837bdee9090e1cb981b4682fac7a5e3018a142;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22c357bd5aa9c8a6c0a612ff8e90d46aa85781bc29a2e97b76ffe1afdc0b7764b3b257fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fca50e74d3e91c67eb130bf80cb715b10ed684c951d65de4f80d0ce9f308adef6aee26b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf84c74e1e9abc67c89e092606e421b97739d70f5289658f18fde7a6b0aa41c058f403896;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h921ecabb70daf2fbf47d879bc8d27715aa62911b04a8c9ce6d210aa9610d620a43257c1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73fc67b1ea0cd1047aec10344e4668a43ee8bd539b73c5020bf9cd0982c75671c114137f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48cafe31d13b69ab9bab5b86276916667a374123b47a937f63f8801bd406313b4857d79e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98f4667f49c49da282acf9dda4c7d2d304255d29b52e4ba0e02987d6fc5e7ef4ec368edf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6eb1805542e6320d8af619ae3d8b08bed8608a835df869a7743ee89ed54393fc35ff975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff8a8ff4b2943cd5715ef32950631f404f00ac8a3325c6764c56f2196851a8c6a452d4da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf3fbad06457e64c38d4f451b76ce9ba1100bd01abdf0343e722a2803f0eb2f5a2fb009d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab511d6582ed7b8c285c0fff96946f57acc4b4de9e69cdbeea87b22cc981880a054297b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h609c7f948f2fd57a2838520872e0d2e4f9bece9b2003cf40d479764304b4c1abb860e8eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae848eed9af25da08f4cf0d9a861a3095c2bd53cd1d42353b624fae8547cb41178302155;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16507fa8861d830f0c01799578585681002fe894caff19cd0e579c986b088a9f98e6010a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1341975d286cad468fc13e17ff3f86ba174773bf15eeabb251559cec408b34a7b9c4d10a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4dcb3246b7c1b94f0bd38a833fc2bbc4ae96248b79160e5f02761fce837c8deccf0e9701;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80a096528ce54315c36394d3d8fadd661a9e8cac1beeb1254cd3c3bcd54abd416a72d995;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heaf40137ac39165817acfc6ef21289197b8c4b16a8eb855e1ecb91415c933416ff8eed1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa70f291186d9f078c887789d8518431301af5e0221b7593293b049d22af89517bee0efe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h944a32f0351c8010bdfa7116a7abd6490da5ad11354ca1acbcdffa8b4019bd2a0a1aba26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7788a0619e1c9b2309d433b90dca0275f4b3151190bce0fa3b72bae0f7a86aa5a804fdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157cc6e6d8633169983a270be695185a404547603756de76c504ccb03c375e9a102966b2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h728f4902fe59d4846f94eca2169134d8a89b2e2e59bb79bdb2548d695aba69067c71ea89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162826b13aaebc710f7447e1a31035e4da4aeb3c435d4b2ba3b6eaf9a38cbb9fd91cd986f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b728e2a301f0a04b7c1c71353e9f2a5a17e50e1036c97018e79506503d1919ae77e7ccc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h912ba649c277bbe2e8f98aba1445631ffbfc233021af84230b51b69bc89f86c9c9c360e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15580cc5389157ec80b9eda5dab841d849eb9a0425d58dbb232c006fd5b95da25c113fff3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafa171974c0f5dfd820c096eb2c1b38eef996f940cded89268168310c9667d00b75fd921;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e346d70a1926a99a673f16bdf10ac91f4631f67a721ab2c5de0fb922b169a1ef678e4a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108d509052271e33b849001fdbc45f3445f961757727df9d6e9f2a35bf95171c0c6df7b04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa3e0e0faca73fe109b6d6cf36b94c7e6b356cb4ee4dd84e5946f2fdd0ec28954fb43161;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee4d661d19ccb939735a3d1571e01ffefb0fce093fec5b216c955b2d9cc69e9d606056d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1136122061a01c6d58e8e59fcdb20acaf5a4ed07a7f04a18c040c4c29f66d3e9fffadb782;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2b41e6a44876d6c3b1eea90993368f2e72ce76bb68cb02ae4c1c2279676812ff89dd5df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h128228befed58c4a152d71ab4426932a3331eeb8e49935907660752920fa1078c24e1e727;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf689cf307c0046505bfc65c36031e71d73e792f84981938fb726e4520bd6c56229859bac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h608e9b29ef2b394b748b15ae47fda4041289a57c3f6088ce90385a98778f9a07b737d901;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104fc343a700401e9ed220f78f8d0d1cb120d02cddeedcd4c634e7d19f64f1f3b8b81b9a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacf8f92bab5488319cc65a8433a2b3c26658424e324c520a9579d81a86fca14099a4a9a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4147d4a776bd399f8a06d33d4004f29268f03a3ad99e88580ade109f4fe6acf0b92c6ab6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63ab766acc7981a1987112c8df257ce872c525c7fbcacaec7967f5138d2c2ce94e08b653;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha20249d40fd9550084f98e5dadceaa0b4a7e810a32ded14180852018355a7ab167a83d71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc3d296c83e1f27a35c1bfef2b300342425a3e371001d3983856a36529145b2b3ee4bbe9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1826569468cf25ea5e2f30cfab503baee6a1f176bf2895f39c2797b25cf71abf50fe801e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135577e54259030da93eb59f98481bae4ca95409e8be2d527ce7c4c75e3c200763aee0469;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131d47a10c744511679fcfd6273400b73f1e667aa6acaf4c5ffadf0d28cb4d73bea7895db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h377ffa2aa857f02adcfece44633ed5b9043c93ed97a42cf4d862ce0c6529e79c503bd82b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10dbe823831b21f5b7ccfdcb51667f01c7bba637c9aa7919d5ca6c5d3e6d427ac530b87de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5ead802b0d7c30f812894e8511f21d81f0e1559873071a2e4626bffcb1f1165d36bbd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150a7c507c3d90c9c654ea9714355fa56054bc89f6b8fff70f2fd46c609ca7e39a6801291;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44dac210be776acb9012fdc913bf0f286486d329049792eb7395444217814aa5c65f6496;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h879e5651ccf9c2816a45807a4565a52ba91c1a23f392669a5afdbba1a97434525dbd7e55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4d76dc5b2e2a98d029643bb8a64264d19934e3a6a1466599a2b7e105105279084792f86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5292af4827ee99b942a146e115730cdb364aa08756f5c105137bc9400b333d4fef25843;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1442df51b0beabf2a014cf4bb8eb2007f7d4fa9e0827199ce36cf4501596db126786902af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f5fe38dad945e8d21d98a7f0343ca8b0c337e7ef739bc581ae33d5df1f106328a1502;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha561e3441dcd20a6258aa5a204468c78832130c658a9e3cedd39ffa3e88fc58ff3e474b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5985509d34da1e81b3f148e4da45d09cf42de018fb0cc36668117dee83ae1e86d985e71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1339df300db756be2c189eea81ee4f63d8fe0c7c4058d3fb61e799f0a55c50d41f0e75d29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce264f407ba364747b98cf81256856f572eefad933962803990b7c02e8486198d3e4a0c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf237e07cc6a0b76a752924b39520fb03f66788bc68436cecac69c9da0695580983d3abfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h693bd579116887c6630d8169cbccb58b401e7d30d695e07bdaf3ed4407b69c400f0d0616;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h347b75090256c9787ad6cabc4d85c0aca650f723ac4655633c38f3a690f5cbb6c01d0772;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180214812d9f11d92f230797fd5961cfa5452fd8ba59d5b3692e14d314e1f2078f4528fa7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda139cbed033a98a15245601bc27ff410aa316737820a6fa46c193831e38ad89ca4d2aa6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1effbaa334605c957919514f4a7c2ebdc3cf187c6b15680587abf89a2497743e7340ddb7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1036ec8708f094a6c20107dc928d4dd41bce82880360778fb93faf02c0617027e946b81b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ad419ff0509e6485eb2e012a957089b49cc625d65456e8e2c9c913ba55b1ff75602d610;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h929b971de54670acaec742851605b764199a25809ec17086517151c9452d5398ac3f15f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfa3f18cd00d8d000bc9b88466b9ca19f046f0b01242ca2cc358a99a50d8ea15c2a2d176;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7d1507633f670e2365f7116b144ea6b3e61e6e1d6a4127f36cf1b28fdf082d9d5caee6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h969b89ee576065770bb74dfa9c021b709561d85733208d9f9dc31bc8b49845d357c351e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c922b9bce9e180195cf52d4553afd9650ce7b9ffb2d18d76ab2119ae9127d14e36abebf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1209d4bec6d3d8295c8ff37af8156af82ea21c0053ec86a000c48b3a08b863380db8099a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1847783f336b0b72fb67b82fa4b9e5190d426232c5c889144d37b7d354dcbcd089ab02289;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a4ddfaf5db5a5ebb915e2211abb0109b33aee4b219f9907a974a2e0fb48a89c35c2d37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0163a738be714db0096941419c635a5eb7ecb66ecca1914534a9ff696bd760acc31bf92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a69637a08d7d64d95c684b39474c2931ffe95ae56910d48590ae4b75f7a64b38e3bd301;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119e801959c4eaf8e3064f589d3021f275ef44b20be9529087340b804d634a68c1cfcfc01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1519dea5c290bbcd25868537dd54ea35f34979952a600b1d55a8331a8d5979bd8d52c4e92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44a4a50ea16d1e35467f192b8526bc0e0670f9308404a3fefde408b077df7843a17ddd3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6b566b2443fea3a92cf5163c822db472a58bb214ac218346984d29aaed441def71a7a46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a91ea1865506a929ebbc9320b26b331d137e8c1997d1e51e59ac6e5dfaae282348119b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefc47d52908fd336c21263e8c2baff377eb4f5196d591dbc28e0525eb2503e4dd77873dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5fe2180a316feadc2093d353f6dde4869fd3a76b3b578024c889b5ce18a401e90e65e59b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h897c99f749c98b35eab9d5b692215b4055d10cb6a5870d30c98539740d21693227312e58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a97b34b3304cdf10c94c0da86c2fe2d5a47ec0ac24b13ac67b8f0541507e9117712ba8b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bc1d600f059ecdfa19808b8ad206e402c081d2d2deb4acd7328554c85055204436f5d83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c2cf860322110bfa92c2a1b6e12000eb3e03e2116a76e8d47957059e66cef53295d8ed9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8b49c6eed224d159c4c37bd7d9d90ae34a8c893985362a16b76849b6d94b9a83915118;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff04e2d365028ebb6e756ab68583890fdc23369da7e45f2db76c97c6b7ed33d70ba9be71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6466e807be6e6001b643ba1b2abd27a74e4dc08599c7a0fc97692b6aad1d9f697eb4a0e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14167fe74c7ec07f471fa877143fb4a2f91a73a7944ee370a69cf363ee7de7ce9de138151;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4baf15f1277927d2cbd154bac50f8cf61b5b652ce6bdb1b56892e1cdc6427e93b8244b6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fcc2baf43d828e0d0ffd79f6bc6fbe03d41cbbadefd8c051bac4578af5d4ad16b630cc69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1071ec9d83a70540a185d75a0349d01e28a130285c7bdf0614e0be43cb53d493b286aa2a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6d6d2f7d4b823cfe531b384f78c0b9283d3cac7545aa1f6c3f4b5b73aec7085e8786371;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7798eccc6e7832c00d2a360f32feadf23f91b4c1c615b8897bb049c8dcd2151f0c56eb23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cf6b41a5a4d144f174338143ecd986ec9439313f666c3f4303173b9c7fb83f51dc08975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe6f4db83af4312ab301ff48919992ac5475f6742ff69877d8380d96cbfbe54482ab1d5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h556ff6cf715be291419c8b906d669232622b34642c5146f7482d993e912fce614f5c7c39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22a9ef4ee0baea3fde33f008424eddc5e9c868239d93d79c2e55e82203e5d9d577dc15d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3d83ed5356e49542a0e4442c441553cb86aea1e3922c078ff1fe3db2860c880fc0c9aa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb8605c78589c0cc241e8cfc3e814d544f3f7b7309d3288b57469b9e27f940d10291ca40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bedb1390af8f44744ed21a400a2e0f461075b84f89411471797a69374e8df846d3a4472;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78d5336d6409bb993c0d3faefbc6508f1f7ce4d77de324208a75733196e5bc1a3d738044;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f84ac9f592e7929fd1f6e57b20f349298d4b62f67456bf1526912b1197446d1192bff0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b597089a9f6ab8a79267271b2b2ddb1ef4e1f077d81b6829ed0bf5d122d4ef7746c9aef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4c0c8013ab284c3dfc660c22d705aa046bdbf978f4d563b60e42eaa79e7c471b8b243a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a513e180612847e7dceff58d6b9798f0143036b1f57ee3cfc09120271d810d55b8cc653;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef8dddacd678bda61705c273d06520dfcd92d0118c42ef595ab1c1216e5d60ba95b84a7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b40d44fad871005ef57bc5a3897d80f6dac3f2e46a8fcd34e07e0d2a7874ead665fbbe78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c9ad8d97bfa7b0eda4d18240726c0210263011fa26593e3b2fdd22c4727db7d2f49e895;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134cf4aad24413a7d5cdf5efdb30307b75dd0b4b4758fb49961b9018b95e2fa7a239a560c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc42d58144359bebd1b136e044ca23e9cd3e78f634324bd45cc8fe3ff1460d341591d5721;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b70467c42406fff013df6380c45e257ceacb1d6f2303e0029cfb8946b34544c691c9ab63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f1f390771704c97a0004a579d8cb1f601a7fd6a6e14543e23a63e53d3debe1344709f34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f64ee15cb76a371b560ace0626ca911653084cf25ba026784344feb4cf42a7fb6f6ca6c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h443308ffcad8f0c0a2ed762337d4fd641518d5d42e43118ae7d5b6b79a7d6a4a01b2c273;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b5fc90ec48335c1fc9f7234c9527857d1b3cda9b77d33b497599437d2a7e3eac4f4f5b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b58ba13b20b6cb73fa1a2f794d019d17d3dee1a8b20ef6b3bf508a4d8f3a6aeb5c0f3cab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c5072dcb9c90340f493e168c3497b56ab320d21faf66a38cb42cf11481bbb421517c4ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179646dc59d839a664e315b03ade630af71d49871caff0468e23e789e7a9232b63ec14e23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e6f54b259df31f334e669cca6ed6459fc4d5953afd2701ef90e944a17e40f6119ca87cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b350e3e0577d9fc74eb18561e83b0c35c3db66a77d43f8d6b5be0294d9b1d8b8d1dcb28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1accc96f1fd16c7498a90ed89db7642a9c066df7645ef1ab5f3a4e3f2c326d7143b278979;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145bab5ced615dc354d902589573abff2be6722522563875cf7610d73c42714c43ad0e1d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4dd897f4c6a14c6c05d11c025d06f5596ee35d450827283d23740890b14f445d4295229;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60fe82bda8f243de9aad56671d3eb1551a8a7eb5c85acb7f2a40cf5371587084db012370;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c8fef28f967bf77b6fdd98926b6c53a17d75bef3f080198f2d4e800c1fab9f83e45589;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189727d8f3387d3df61ec260cdd2f34db37d631fa34027dec37565548e8f281fd7248c47e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f7fc3b7fe1ce66bf4fdf1ac02b807dbd487b799debad4793cb8c7547a12f9a2be8a945a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2845bc673954e5cec1a906102984ab4c1293b21a0a04edd0ff7dc686c9e08685685cee66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1babc7c9c3d0cd9e15ca5f7c4412bf1643dff4b357354389f87ffa533f5ec715591fe5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146a6170465d0bc2a2877a8c8cda405b9340757546fa8108dd76f0d71c439c9c0a19a7245;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66aabb52b33d4c386a355b44cb197cb7f090523e1e1dabb2f7638beac8074e129506bd41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a25ec30f8e2f25bf5a0367f9444457163017cf77c57b2ac84e839f9ca4a93b1cfae5553;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1386c853647fa5d7ed18521b9462ccf367b588273d1d42e45e08c3dc28f6715bd883bcfe0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4fc1a3c088206367b3a959fe8b2034b253c8cb2f9eb2d2ba9e9c6b1be071f837e187129;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b8a620d5e39e8c5b8fad3454dbb32b612536b4e9d172baa67ec2dd58499097c678af35c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa4374e210261b7c3cd22af47859811ee6fbdaa60a6bab177a10685e61a19fb83028a035;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1754a65826554932b0a3a1f6c2a2bade32b9bedc71fcda00fafffa0c5a1e7326911ea409b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e86aca4d37b2f03c50ab7a111721b2019e8eb1e59dea11bac5ad3cb7c489d4899e9470f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5545225f2c707dbe6371af09aed5ec55580f4ee23e09303d8afba4daf21284a94c82a33f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132f6e77fc8666e15f7e11e3034766cd21e77f1f870d8c63ea347e6096f39ad64f229d672;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cde83db06cf8bf0c1b8fe081416f17cc352b4196ef44fd5762785b038a9ba8d0795afeaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h855958cabfc177622c71bbb5d76129d757fdc35f427eae9f40aeacb4a2743151bbe9479d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17373435452c7ee2b866ea50d75062d8ebab1eb74c50a4dbae762b877c2e09f38be7c42ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h780f67fa92db4462c22f09cf437eabc2c8136fdb0945607ba611602dbb8a5dbfd57f228;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1388550717a2d390d6a0f35128e4a1de145e3b2865318a215eb14afc11b8189e60b0354fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb886a3bcf6e021d7a8be909cf4749d013041235974287bd96e369616c0a14683d40ebf4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6f3e06378d93169f099fcd594efcb9aaad8a715be8f18892905dda752d419f8ef77499a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefb9fca206e880ba2d56d6df4d09d12c500d0b45f728c82d4b938a99e715e2a7339eef1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ced4e3d88c9ae2310856680953d5dd59a7ea824854669c8eeb69b89012709cdf79c92c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h275e35a82f89e14e964087d6c861c3aad947b3d8d62d713172d3d745787f2eaceb99c74e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb27a498ef23edbf9ad2bc79e7023856853743393bb4e132274c03b74c0fa0dbdda640f8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8e00dfe6991251a6f498b562bc5e020d756a5829a2f8df95a72000a00121b9e07ac11ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131ad0950f0dddfff06e1c22a22cece0d56fbac877072daa4addfb585256258d691060c0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0f58903590787d42ac1570f117406708ba54a04376ccf35b118e3e83d5e925b856d9d7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h443a372c0d4d3b8bbf1caea64f596bbabbd079864c2b651a18744f3b1a29851234824f62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h610b0c3c5782a519823d9b895c4ae25d95e021bc1a9464781946e71b5b0d710c4b2e18fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfa7c5fa2a12a4b262d58e73379b4f1763f0072b79ebfbfe4e9fc9fa9fbd3c2449f30914;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha42b88a11d031216ac8dba432e612d063c37e4d9a5d5e4b4023cc03a99f02c65a463f44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6bbf308973d4c75b253d5814ee8a071a318a32d5f9f9924d77e79b8fd4a4b6eb44fc930;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100e85a5350868fcb96e9a56989f9a58186ecf7eb32019bbb57b9d46d22719cb26c9312e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fec0dca6ff93f90db2137afac73228c5baad876bb6f8f9697c40322cad36a1c39e0127d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196008780f02e088cda980ce2bc9ba60485259fa7d9504e5bd9e5b8b671941c99b27c6e59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6f203c48cb519a7761b43f7b7c0619a9ddc1265e17f94e8ec098b5e9f80e381509ad846;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146835e2cea6c1512f639aa73fa1e82ac0dc70d6cea10848d6f743f237a0070c7e1d2525b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc031a8c1ea6f4dafd6007f8ddc020456f9e0d386fd4b4bb3f24f6f5828fe8d65ef8362f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120579d56f4c945d17c6849c94301f13add92637e6aa203a84f2c7aeeefa161bac18a4407;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fa231701f4b44a4823a32751a087a5f8b1f7d7696cbd612349c92d435da8967ccdac03a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144f91216f5a17ae4b186cd0022911fd17ca0d98c90ae4453b9db04965150c3ae7417234f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1787c7abfed3170501bccf77c11381d67a41289c2d16cf24980c26b1d35e046edf1db4ac5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a134be898663d65d83cd49a33891919ffaa8ab6c8ad4b41b303ceb4f71ef98037b4559b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1471969e484a6f8a57229c0a4ff46aa095a99cf95caa556a655a5d85b85316d57a5cabcec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e942ecc0828165788c1f75636d476015c565d1f979776c43e9a05ab5954ebed91a73f41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f6e6ceeadb2958bdf2dd85215ab02b04b343b61ec1a0682e777b0eb019a39a9d595695d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19af4b1512aa36530bf15826b0ae3924fab67a6185d090e1f61a1203af2739e7499d42086;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbffd4bd43a9b369bf0a06fb0d5d429dfd118b51ca3f6b67974f079cee8ae828e671a33f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he10029af66d2d23a3c722ad562d9bf4c7a5aa6371016049e6bb5299b1b45257a8706e778;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h566c8d6ca2f6eeedd6548167197be1feea0514f254f5ce5f81fbbffaa6d2fd602cd02f72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f6d1c5174a2c59da3f5ebfb934cd9730e3ca67ab298e0095cecb9bd730c7cbf92e8bdb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d44968b060a61ec5dd58d1b3e0fc1d657fd2951591601b714df9980fe4669404be7513e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf13feac7bd9883b0670d352752c3910b003891a9366ee234f14ad9052e1ef92f57a939dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a40801e51ccab319e4ba2b35c85f801f32423acabb79003fe1800878c748b6f211ae8c2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9a030d4e293f62155e779726c503f80615f22740b3264e2b721aa14d94e0eafd5b26747;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b2c4168c6a3582fb795e28e5f5598f5540717a799fca250fd6cdc93f279baa0b5812e24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15acc1cdfd6bfd472ef5876f99007f042fc3626801e744afede8a28fc804f10018f699ff4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38f2ee0d311a4c0b6298d8e28536c39c4e2c65e1daa1da941eac9fd23b748d3720755c09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d624f7162bd27f25b58eddff00c7e9ed751d026c4ead134fc171c3ace4e6df676f69c7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he020ab6824b6f6683562ff9235cbc5109e3f22da0532c97897331d2af7dc74f2c27c4fec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f302f6b23959b2fecdc99378d1382a50ad1950423f93ac0656c545c25df0e3ee4feb9a7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d16c4f62a191da210bde28cb3ccc870a92d03e29f322ade95650cc8868985e6965ff742;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184bf96f2564c4d33aec858ee1d9ece2842508178687198b000131a24c6949cd014e94647;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6edbb061cb68c968fcd8e69e3f08a0cd20281d024fca839f663d6fc4d31685e76469a3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3d4e749e356276ec1c5b5b2228ac654e6930121a77d5e11965187d8486e1c9e6eb617cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b24e0b683df57d35fc456b7b2aa8b423b2b6d5a97adc2e55b16a45658e88a433486971b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f5f2644e633c7ecf703232cbd35be0e4df72be702e935daa3519934aa7a8ebf1f7d3628;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165b530693e6ee9747e809cb6da596a74f59e27c27df7617f609949fb7549f2ce065e120a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17563122bb8f934fff6c445b18d7170a4ff2121a8a16c058da0bd6fb0b5aee3a64267dc5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb94da94a87b6858b22699d04bb2292613b1271abcec6af5542c3bab218a4520385262e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d93973c864a9dd94d16bcda17ae2afc28fa7c8e05a4b0a305b074cfb60915f169a04960d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101213f98ed973311b5cbb2e1c53c19793f70d1732da14d96e88df0df3fcbf120aa752a9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f535c288345bcf889fa211332a6487e0f251b8d60d896bff81b7fdcddddf4e41b2e997b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75727c712f7d870ad7e251ce4c42f50eaf5d551bb548b11a223c72702b5217aba4bbc6d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0be94f916f4336b748c925f985d21e5426baeca4130727497a9b7f92f6b9aa55806c0f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26e063e9d2f18c70e656faa99203cd1bb6d05f008fa131b1cd6d7c50db273a204a1e8eff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4795bb89cbcc5d51f4b1f3b728f2fe203b921a2ad3676aea9f7ecc0f038d2236996d6452;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27cc8ff641d45c54f90f02eafc78487a0d6eec1158872032ae6095a692e6f094263b04a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d361ab011a8722239df539cf8c3b7d3967c1f7cc8fa74b91c192fcd14f52d6e86008c4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11caa8bd6fd4447df3665beef5a9f5e2fe23998dc9f9d988435972ea5604be9a53244977e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53832c965d288d6c6a1bedf97807062964b6fe5fb30f4dbfc10c46218ada780194256076;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150ee1431af35bbc732a2182edb9baabc860404cbb35a4a4d94c431d85801991409f9e6e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1474c44d7eb63191c33a3c0c56abc572a60d675af85cf94138ccf4d05eebecbbe781033a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b99d60333af3f49ddff3a952fb6a3ab6fa84ac7b804b62d77ff3f77ed09c4c0dc6e8f19c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0e6afbcc05e4350932c688a851ec03b04592397b881a09ef447c64597cca7eebbec6c15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11776a3e848e4a457fb7ca7cadd429ec4256c7035273b7135531af4770eacf64a294d8d9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bf88aa7ffb97ccd9d30d4d63c7ce55838ec96aac82d9dae5a6ad3568484bf2f8f7d72ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a778f91bbc76daf3f215a98b742b999b3926a4e49fa4c3034a41a5c9a6c7bb30eafd874f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83c60208eda40feffede9a435f8618b7cad12edf037a3655c0f5e3286b54f2f006bb7ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc774d6b5d3495011ec8c72bcc0e184b6b563c72f66b2a35da270c3fb9e7b739600cec504;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0e7ee76c092e04a856b006fdfaa6eea405b01235a60dc5303a19d03d057d30b8eceff4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa3adc89cea4b96dd8c51397adf56ef229550aa66b2bc5ee7082444c4f3b18fc945dc034;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f78979db6e1eafa86b8d17ff1d716b5571d556f62591cc5b128cde965e1f9fbd34950792;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e067299db5e26fc4257a572cab3099d845987434e37e159b3b33f2955b499d64c803a844;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb7f99c79fa8296b5439582852443c864d07c01792f442b2fe120e27818f4de7dad0db37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d545182bc77beebe5d1b4fafb69f7e4a15f33ff737e8deeb8a8c9a078303e2735729902;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e643ea3d698530a94344f99ed2ac5a5450d527324a75014a5c0e82346801b9445ee089d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10917f4182ba7d8484b2ebce39ee0ad39d722524c8beeea41002d98f818eb0b37014620c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6979062c53eb69eae6a6b2d724c23045299b196a2470b43f1c64565729601e09de29b7d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h490f552747e0ed2bff355ef00cc89f755ca2bda751204c1dbf5b59f3c1bf6ce6ae17f42c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a3e664344b75baa8842c27a1de7173cfbb6c378d306a70eb7dbdd803415080364ac9c41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb85b4b8798d1f75a72d630fefc48ac8a31e0b7864968dccec711fddb575a5a10abac2b41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1fa859f04f7b006b0b671e9e92dc0099560d15a9913aa13247145ebc8c0ea2b59dcf0e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113f51f282848d812ab8312437355a53a78be4527f44fc36cb7c4327fae0bc8c0c86c1123;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f5541ae7c21162701b30dc7989e046e597d83c0c90741f4baffa46536c41da9c4420920;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132f2c3388d2e74276e507a247238e9c664c405a9bebbe0e938ce7cd4b12cc1b73e2e51ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf40a2ec8c1206234d39a9beac9557f374230e04276f4428eddf471481c74d76e1161baf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7eeb343faa5618a3708d9d685fa97b8afde413db4b80f24975a3e8ce5ff3689afedfe949;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1097e899057909d03513df52ff24467f11befb57898903895ec0bdb274144c4a73e064947;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22917ec8f3f0624b0c8ec09a8ab7573aabd72beb0997f9bb6eab4094e3122793419e8959;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e6108ff388e4229d6054a2a434333316d7822a0956740c6cad058f6ef0ed6a096ea495a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3acbdb9867beae9a395c7d63c6ced1379103aabf62d5231c97355e6c54e7f2090d89b64d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d0d194e398d9e904bf9db3268d201cc6a91c2dcae14a14883b7f903cef7c4756f7551a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacf380795a49720fe2c793157d2f139f20f1600b36f45e33156745ed7946ed46d2e0ef14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a9ab861a6c2a3059448d69e85e63f74aa8387d25b493ca7afd2f73af2356daae810aa4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa621ec7df4d4551c83e5ba8806a3a96f01f248eb6f6a73bd49e6585c1379e6f9502a993;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb452de9892db953f8f291cd8f7cf0d267705c1df5e456a88cedc0571f0fad2bbcb65ec9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fc504a2a96b11a4070ae49f66c214e164982c0339d066a57954996d08b1ad47162c572;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63081cb6b57b87309b893bff1505740232de35c0aa7f0a3eb95e8425d83dbecace85950d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123de349cd64746ee57fa75ca5a5510ccb0910030561a8bb7ec22a2562aab37d3000ece7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e9361a7f316a52799b8c3c03a110c5274ebe91253bfc288b0f6cdfd0c655958d7c4271e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed6ee6f730c4826d85e9340a59788c6530e395f4d72c30bd2fcf5e8491dbf44662f1c70b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2dd6f0ace42c7895aff0083b183248c69175f23bd43cbc38aea6d6dbaa41100cbe62be2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc853ebaa7fa3556237775942172181631a1da5adde0136fc50ae5dccf926606b2e6c4fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8fd34b90344325cd7e6d32dcf5407b9cf2fb562ddd233185512d1c107b279e7a9c26739;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha45a926eb1b7dfa84e4701e620523e8caadd40ab36ce73e70b84f9b57141df7582cd7d77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111d61d63a924b6357e9e484392e6048f4395bf343ea5c6340170e5462a34c3bbfb7ac504;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151c8126391e7575f89d49db4598210a8c95c9bc0f7a4a7d367a875b33904119ded169f8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d09c0933900c29b828cfd2743115775ed2720a366c9d27de647600ff821fdb4275b918f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155e6ecd0aea21a14b160e26865996a2e0862a71f2260c75da6ee57438c797d5bdc0944f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca51f34d135befbb51904cdf1164f399a78b7f995ee30c12e4ee1764b538b5d0ba98ca46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb04bf58a06781ca49ab8eecfa20e851af537406a047cb4755ef3f098bd00eb69a0d284b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca3bef9304ecc6c2ea6ac09172fab28749bd1a5d5bf4041452b0aff1405f146db5815561;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105422e08fd1289d51928d6ca3fbc7c22c7537ae6b8a86527c6c0bff1c32c855d971ec74e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc965343c8795d1e93855edd5d83ea712d03762286e0852a47f3440b08627fa7b7374e148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2967336fc574a83ed7f37353525de6d817203f092bc18340746c479b256a4617b1a6e62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5be07f7e786f9273a7fa4c56bbec4ec34c81f99ca90632abcdd430a9f3d28383e4e144b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2a404173446d463c09abadafe1ae7dfc38db51b6b115c553445777ecfaf15f32b8488c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h224edc2789e6a96ed49a2b823455bd61b22e3bbe0d7deb63d548d93f675cd1ca4199f95d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b298efdf08e506ba591207bdb6c7c75bb93b0924272fb4446aa0cb3d5f8492482ab9b81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c78a7db2d4c789263e189f5b1df4c2748664765a3c132ea9eb15ba7c0e79903a16f9d9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8f2e394b0490dd21a9a36b22cfbc7c1f6fc76684ed709d30d25c811271eb8e7e87c7d20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1476c322fd6d0edb8856ac4c5c2dc1a2ca791bad809f908017d4665f25b8df1a86398f71d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87101419c19656928c3587955b0ad5431c48725c2779b90f70df66474ba76c01114514cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a75cb477310efc5ab2ef3cdf049fa60819b65f5bad9aba4fb906658714bae23e602f2ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ac1840059a5e40a8e3d1ab0587d199e044add528a0a941c09a815d3bc7f7102b988652f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a8a85f3cad03d85b32c98d598cb798ef58ab6f5b53beaf0a35adc7c0372547f9736cdef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc257371eed1194a199aa4b1ebdde8fd210e11e7fbf545fa00c01eebf4955cee64d21ef7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfb40140197ddd1d4b80f0b14cd0af2aa889ac92082ae042cb310bfd88985b707be84e0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac3805d09e9b02678d23110306eef973ebd105b39cef81dddc510f55c2e3a2de31146018;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb74ebb7112284fb4933a7ecc13ca42bf72543d7948d92887040d4801ea27073b7047bf00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68923481284e8deac9d86db4070355d0a2023f0db75821e35c08a61787ddde961bc0c7a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0135c6cf6ccbda1f622fdf0a560f4d6fc0c5320a25d0e97ee24a2590a10c00b0f55a4d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98de53ac700f86adf824c7013d4efbdca016c15803454755f3329f4a32ab726ab144f730;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3017f258c38b34baa0c4c93065973de1533eb0a8a126913e8ab49ee5eb9d0d647695cc09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha84dae6977821468aca27e7cd0929afe057b338f625321d9c3da8ca3c5e95915126192f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b389f5308f0a8d90a6f1e73b441c0f7def3d688a5b96e3612d18532fa737dc21e6ee1f23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3341e5769f82f103991bf781c8be5b1a80fe26a3e82c9110de9a9cbb38a52af04c73fcee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9a189dc93cde824d2e9106b93d534ab2927a3dcb48b0581793e3198f3df3c753a05009a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h910d62596391f81a670128f01347bd4a7458b73a5e48bfee18081aa5479c71c94ee9a5f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e8ca6086984f1cafcdf78b7ecae7e750c28f17b3fe6c01eef07775140a02858c73685630;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f5a6cd67adf15e82b99efe5cfe21f4abf2670e6d5e6b19c3464108b93fd52b339cd2ee2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12586f664fe68e9bbfb5791c38cd1962e541423362e6155642fb891796527c313f385b33c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154dcdb90be27b124de67cc23a20883fd05f1849a09b3212d29ff2ccfa1353d355ea28d8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5a2f4077fc3fa488a9f0b4571a5c56ae085d6176e0bdb795e5872768d15c9b488be04ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab4b206a6c20e18811279926ae59bb2ad4f56ef9e098ecc96f0c77c463d616e1472de4e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he916afd0e7ce1660c6fc0a7e42efc2240863b22de5e46344d9b4a6c5f406b0adade0429d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121ec0c85783c2f9fd9576c7fdbe55bbe897a9db0a66b23a1eb6af17add89f40c66e07f84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79223eb5c642e8de82b036d7340f90025bf11a47753f4073e6b7fac71ac564774c0a503b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111d0c9f8e63c0e23c640c5597b5eb3eb3f8b5682507dd096a6442119acb5a87388136996;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142c3bb8b87b40cc74177ecee0c47207e347897e135b243c8e3b9e5ab0ec5efb6e4f6214d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h611de33bf85b9c4d22c6678ab685d6971b16ce44736a1914b30f9ce67b9d4a9c73afdf4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0b90a9d476659e800b94d6b2bc686073ff0be4a5c0a67a052263253e006bacd4750bc29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f193f2227141aef6dd62919127f0d145e397143a92e9391971a623f3e66f840e3d8b9cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bdcf20e977d96a1a60e5068ca5bf75236435332759189a8a388a1a7d2b52450e4cd2fc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a40a1bef042f5d079312673c4d930acea603f14aa2061dfb3e26261874d089bbc9c69d42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h729ee3b789c816fa88bc89c2bacf6fa64319e74436a819cde28d9fbe860bc652733b0820;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h558578370f6de9709a5e83b1ad1603fa6b9c054a2b2292c022e722974e73de57ade218e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b032ed12504b4f92bed307d6faee9d832d2492dfc07984967ba6e8ef40c165af8486d253;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18df275b970fd9d378bab7310c56aecb0bc091c0e56d2081a6a6e837f7f4270f77d68980;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100f9940a9956ff0e85070947e6f5b47eebf33ee58d8ea9cd7e18dae582c8d1f84f74b3bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fd47f894e1f902bc5eefb1004cc36c626c3494fb268a2b4e057db1a6aec7782e655e48b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a7369704d91d73b8e98ea3cd3e8aaffeb80c35ef40d886dac781bbba05f71cf4430a517;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9e8552bc0670479c34f35ce024c6ddbd1b023bb966cc901a05f8bb6f635a767561e43d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199990a3fe6c26219a9d0d97e73dbd062d5d678cdb82b765bd5f06b04776a3199ed82c367;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138fa3aff8664ce0ddbcc69c09c4bfbb5c1a60690c25fadc6fc28e4075f3a157ffd25df2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198b3fa47eeb511e5d6a226d134e79d9b469ec49ed8973fa490a326a5dcf96f7ba4b02dfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2bfec72784cf8293e65dbcc6dd55b3d3756efe19c991d111fc6d3692986c721df03ff0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8618e0f223b543c0e493a1abc7d5fa2b819119725fdd5f3a7cb86919c0a0d5abf96bd792;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172522c9da81c927ca579ecc96ea53a28f703ea91ad35adf43b050dbf3771cf1b8b7e8e72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1059c7ef8fcb747148411c94095a2f57c15569edea118a1730da7cb8f57006ba30332f23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ed4f562b2f50e933c028f0a2e017d8af10767446b6b8990351d1ded6015e53c8c99fbd3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21634674c9f3b6014a8dc6df69968798000839f0a2e57288f64f754e6b40d5f26444fa80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162f5c7e5a5215383352468bc307ed0c2871170891c5eece5d7a2aaf85f48bf9bcbdea889;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h351166ecb8ce1cd2191e10017558ac7fa95df721774ee31405d9ce1debd7dda7f9042d7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f1872ba8ab63f01fa3582aed807274add9d69fab77a4dd4053d88db1480eb0254d75496;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cecb60ac412b4296bd836cd956bed37f8dae944a788794ed48c3058fb95583396c79070d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h702a670043e9ae7515865a6f0aa6dfbff7554974bedb0368f4b51c4674d24139f8ab475e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5c39116579f85412ff2d781e09f6e3afc1d6a88da1acca5adc9429dfff0531384893d5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b663cff69ace312947070aba3e36701cc80635a3b12915edaa5b8cf3c0b2a744f003c61f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fc615cb51b6359b8f9bffea85f4db5cc7d07827c1371e4064b493385ff3e31de02e6c1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5cc8fb4238ad262f14b5bc68aeebb680aa9ae2405f65ac5bf011da780287f13b292dc62d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9370762c4d79c3c0822df359d0beb53a53d00e8b24aff99742ea0b46bd4e3c9638dbd84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b769abc3ee7769e88a0267cca834f6216ea486a69df129f633c99009434efcd4e2f4684;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af1fd442e52afc013d3d00f83dbd2b4826cf6a1481aebfffeaf31d585076cfc259e8e010;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13078551dc6217455e50789d96fa882aac12f1edc2d4ffaa10f76019763342242f7c31bb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c5b353a3962e00ace435a4899d92161b16b01a516b34899c7a30eb007e4738a31579a38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11dde892876221010b1d450e8c3f5b9953abcd2a985578e64a091f935e3810dbfc8422069;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1581efdd4bf625923b6f8ccd3371c20d83c8578f54d679f4cd60e314ffd060eb94d327fd0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d0571ad25538abd807029e6d0cc7c05151148637ca41de43ec957f9fe38d58e75f766da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1194476aa8274ddbe56c18e257bf4ae5d6aae871538dece7199f170e070cfebd09dc9b8c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb457487178ba775f0b52bd042a0df311922addb80262379a2dcfb54c4a5ff563d4875a70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82eab44d41ac755edec133e6e0a17c5ec758f3c928d903dd6744f7f06d17281a6cd04cdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1976b85ca42ae34fd3b6fef0d3172d141d247aadb655ad94ce0544a40f2cdd83217a014be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c3f97a8798019e60fb77de22a3f4bb3f67fb8c4d7518191864e6d66da2d0cc668c02af1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a35ad19150f90252b0195c04dbfefce5e89def9523a4634115460d74ab6aa2a4734cbba2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h961964b3580dd8e884ab8930ba21113b26900d8c00bb6c7fad3c6c70a4b34a31d55a746d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h421fdf2b4bc9971abc44e7c6074714685305beb311968cb937f6dbc24d82b40a9d0aae16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdb43e5fc1002b43e63376b88a298761435bac8246e44486416334b9e8dc67d2cd475047;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h406e80b38036427a72154af00699e0ac63d453629cf3b77ef579bca24a9610e7b2cebebd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113e2f767f9a38d142ccc188ae68af467dde2afa0ed9dc9ba554f7720d1b090558360bba2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac8f3d9fd10445b8080ae8eaad3de29db5b6435a6e7df3f933ce5c42c2a486eab5f3233e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1406792340a5ee5abf4a55a59bfc44dc9171cf93ced68b6bb513ec04f2cc65f82902472d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140b8198574662a55ed445a607d8b5bc8606cec4edb850b81263aa831363fbc0bc09df952;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89aae319fe37c08ce1d50fea71ad8d7ef736ac259706436fc1a4f6d35c849985b5a828ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a4f949c61b9a3a5a2be661fd0f52c67a7770d72ee7712f9c1a7b638900882d78fe4be90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he38e543be6cf86e76e2ae50bed1f25a64692ea65719b76c1ccc642784c1f32ccc2ead902;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a018ad1d558dc74fd885649efb3a5421dfb9de6b8d2a9efbce19559f2058d41b2200435;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137b4288cb46b9cb9ae08853592d41a10859e640487bfa395cc338cdba50a579c2efc92ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169b6720d5df6a2eb32ca0eba00903b0200d279a16f2301e6b496883f1bc42016bd2eaf77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82d5e161c01dda2de08f63b45dba1b0dfb76af99df06d2aa56f8a8dec4b549a0aadeebab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168ed1546a146cc32931a18e989fb357413a58e43f2e6d80685052d85dd7db2d352edfefb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha88022cb9cefedeae4cc01f4fe60ec0a89203be4940eecf5028e1273a8f9b44bf6227d9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d47d3dc0ff320d29612b5fc597e1ab15b950a66c196155b9c7d70959ee4cde8a9cb51d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71dabcd4ce5c2dd067afb891d0655220164a8adb381438701d3a1874b527a62a75d080cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180e287fb019640dcf43a5ca3543f248bc47bc86a40f4c8240fe7327fb4f1061fe8f651b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8280b66fac44549c9bb761d923076608521128e66f7fccc1c036947d16cce0f50878a42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe9a52ad7d879a83ec196cec40f804ddd5e22715267834c7e1a0c2ad095a9d4d3f169763;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6f6d832128f9d3960d3dfd74940bdf77704f5ea25476f49fba79904dae022015916de69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1e2979e5392a8878130ce115066defa99e66c2033134b696c7ae6c52d9cd4f886f1bb3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1ec37830f0820bfd7814c21a6134bbb2febac16d2a7a047e689ba84d26a1279049132e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7459543f315e1b954a1310bb9d232bb3ed36ffcad04496a2f10ef135345d4cc3ac92179a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1796363af53ff91a2f61a881728a742455d5829ff31bdf176404391c560bd6cb1d14992b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0e35b4f8956e6fed545a2aef9187f56b64651675b36715ae72457d6eacfe80ab9a15031;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38a50693b13bfacf3d6068c5bafb4d8b50bdcf28cbbd3a202464e54ec773382ba70293ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2508e0a6d581525bf90bbdd2667ef55f97164450ffd3baffa611ae1152ef08edee29638;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab510e020040d2f9cbcf66fec8d15be380b38f089c0bc7609de1f0ba7b4395e1545db7a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h364ffaada0cc7d7aa681976186a40276017d16e52342a706ba81f6bb768336476a046d1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0273c703b447303ec7e53c4952c8be19989d716dda0ad4867358c4ba0be67b540cd4aff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a5f393e196547e7af3f1185fb75ee1b14ff0066d5c88e4f0949063eedd28dce2abf9249;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162b6346ff7d75b87262c64c5f174f7e50183fdc965e6444c1bf02ffa6d8e816bd781ac3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14754d93aa456a952854497c1f0b23de1e5b9ee89ef77f47705791fe906101425fb79d8c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a03f4ad9254faf95eae6b478c8b67fe36772e1280db27aaae1108190b72e50d4165b2014;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h712449a8ba6a968da16abe6c2d67d1fdfffb321c4122e9b88e0ca846d7113b4add69310;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c765b9b450a5bb481719634799597e977dc37360596ba2a52cf4f1ce642acb0c8efa6fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ac328865ea2cfdfb1afb4925a1f603f06c480ac34b972b8e8906e2a81fd2717742fd44c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fec75f4fc877385689c63dd9964d74b5993f3b13db15c174025e14779cbaa5b7d039c15b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b144b13de4d808ae440d9976cfe5b63ec63cd974dcd48924749441d30c5e5fd292b1d75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e70a65db7cd61fef3d7ce9afaa328ef1fda8ef510bffe51075020e32550d69a7455bc18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f557afc1804d06a1fd8da94427a4280d8388ff69377f11adfeed1158c125d69bec1ca82f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb09165a8f495219ac52ae322bd8fb911357d77c8a9328dfdbc2c116eaa7774c61e21bad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dc3e86f7a46a347619f187d814813e8bcd50052f5bca0a3d6e1275602594422804f2568;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e0af5099bdfb6c9e30d0f8289fe20ab0b3fee4fc1b353c4eed6652c974fa5f60c58917a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185b9716cd563f5ef3ac56ae6ba9058446d42979e631b7f031a2a6b9ce0c6e4cb99257266;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2c16e68fb879a511a814bae9cfd40b3a0bf79e953dd1347a8f8360fd76f8f1ac252e1e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e3c28db391ffd4280a9c868f9ddd696fe838885d0b8eac8f40dceb1b6535110fa12eaf3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca162bfed4cfa0a16edee6bd7f3bf402bb54009323ee78dc8b64a2a4736c76addc98311e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdf1e17c910fb68d115fd47e6dad83c27469fae0dbbebcc1c656a687a4f88244ed595497;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18624b5f414c1d62afc9b047282878e2c4f5ab3a6fd5fb27ce07d3e4081b8662c989b85fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3203814d2071d352e9feaf866ca0ab559211fc4e8f81b70410a1b9123ba53af7fa138c43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h707a92b34c9a971a2516211d60d9d2b6ae7d1653e1024539772a173ba568aa7273872a9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b13e5d6d45836cab38b3798fa9a4d011a7817257305820e82792e6848c62e816635b211;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb041ecb3e6085f193a21042873d42ea2102d45952484076b6e92c1633ce8fa4d0cf40783;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1a9b4045c7a9e2673e95283189df66c77e899a50995eea07525e733326c4ed24fa35927;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6aae3b656ff1850d902ce6a871e74d1ad540a324667629470ae6f225b5f1aac6edb14da0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78002cf05209e3b8f042879d502a44a593cb830560398d3761ccc16e7d535ac7cff648e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdbe75321d7af959be4bddfdf7f58fc9befab1921ee98ffb2db3b22e73294c3759c0e1a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6761a76cfa728f7b7e78784499df7f41af260d8889ccc2693f1b88cac1b081544494c21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b6f0d47fe5f10c17fde3518a6915b5aa93e59830f6910a2aa89b3ece4cbfcef196007e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10338b3c7b7dcb89c32b033637cb960bf8b74dddf0759cfbec3950ba33ca0197e44aa335c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52d65bc4aa640c90ab17537b39d6a7b7ed307233fe50a05967ec276deacfca749c1811c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0a82d896069bb9856766d35d9cc7d60f46eec3fc9c0f77cd53f06f7a295831de1f6a05a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116a19eb4d8095293f6bb26e5d5b78038771d54388ba90c63a6a1eeaf96d1b18ef4bdd228;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68ec6970c342fa41175cca3eed39ad32999e55709984893a089c16063c876816eada3007;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e743a671ea706fac46dc9bac5ecb87cdec32de1fdedb126c5a1bf712a0b71ee7fb151ef3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14595d310923457ca51e765ece5d1e4f077b975263c676b75920a53f81d96d62a2f5e9277;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11069fde845839c0f9652413dcc4111cc40fc05d83c60839a84c7f9fadd62140cd238803f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1857e4a887c94208a5e566a9df5e59a3e6cc2c44380cbfa2b7245ddbfe6b71bf6c4d23a79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a4b7d0ea5a36e54ade659b63e48b307788377ace9a773d7a96f4fd92c793dafef42e553;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1baf8db85e004caf50460c1fca694ff422b1f2a2459ec56153ee82e8068db9e3bab4dcdc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c02c3bc86beae2f7ab1b2d47f8d9edd227c096fc61da78b9ebf23cc112099a7338b9c58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15442c986009afabe4e1ef7c59670fd9ec9b4e20a842c13846a4633b7fd726487092960e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d1a32277bcaa84b44a7cee4c3ed3b8c65abbf36d90be245dfb72ea9e4f9943b7efb268;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fa5f75a17568cee3d477d0bc8f4bfe5aaa07271190a5ac80806df6ce2816d7ef884ef58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1143f0a99c2fb0f95c68dc83cbec084bcf9ec5f3d7ca9ca57f1ca7b51e7f9a866d189985c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be3e3d99da898c9acbcefef998573605f7397a5e56f29e339029c83fa12e65e0747c06a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1515d7c1be34b8b57f4a400aa3720228c352c84d982faa17fe20053913d9606a8742c440b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8575a666d6eb1370e6e56d063a35833a68aff5f7dc4e706bc504ae76fb950354d8f432d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fcc351b6e6734b013068e05efad2cf5fa080779ebb4e2e4f7f4a415d26111cf9ea3c41c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188f23ab071fb4578fea2688ccade977b6ae4d261b7a9c971ee876b895772b3d99544c199;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8c51e8686cf120ce8359dd554729fb7117af014ce48347ae4b4384fad47a522cd59f83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139d47faadee4c09825a3f0a4172db0e01a19be79991b641082eb491dcf538e5b47247ab6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191dfea292dad84f98ba552480dc5a2993b7bdcfde756d28b0cf0e64f49ff699d5e7fd464;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d84aee4f49700fb6d0d7cd0dfd0894d56cde8c0fc4d25be3284ad5dd3462dab23cd5362;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac0b0aad12c3746bac1da96867d5ede69c266f4e74674ca322b177e5128a41808c9e4886;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11129216c26c040b6edca50be2c1e72d1d6ebdfbcfefaf0ac2a9839c3a938fb7158c7620e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d5414366a436709ba6f7914082267c31307daefee119642b8e63489f85cb9538b882986c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3631e45c1dded83d69818b7a2272d8b6b98965b99a5f5bbab25d318baaa2c6134329f44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha64aa12a3d7336a9d5f881e41fe2986df86338151030c86fb7ddf4851fba7fa92b9a6ee3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1f176f40059164e98370db40e05ec4682329f7a5e7d78470bc150508d3c3bc36875e92b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cdb7bd714027b1b933a6ce77476188c69a43381c51c6996257e5974bf9504348761d4bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc7a8ad1e60af44bbca64ed9cbe4c5f72fda6e1a1b48ae5838893f3f3cd72b609237f263;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1787d0b0c91098b6d1883cdb789a1c36f835f786a04f93fc5984389a80a6d3f6e05c6a24b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7e38c678cd2b04cdc203768b4f9e694e4b2f7eaed4dae5b90a8c5322ff8b41653ac2522;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135d94497604796735ddefbb56c6c47eaf873de1657f658a61f3ebcb588d8f28de3bea821;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdd74c9e5f1861a15f743adae33e3fb132ed1421b409ef972a8e824dda30a3c0255426a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1f26a5a45a9a34e4c90e87042dd14b7cdc013d88a7650ceda9b63e9d33744037b8662ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f323b2473c0890e5412793bb15df6ef3a22ff78e6afafa100f3de1d561c9c2d11f0f5be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25bfa3b46aeb49ccf0f2baa876459bed693befbc2768092c5a491628266048baeaf33c0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbce59092973f3f525817fc4a3281aaf6bb48347d21996885ba9acca33c856b9a083d2b90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51e0fb38ac6848903916015b7e76e8fa02470bc60db10721befb58fa61c128caa8bde8d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h685ccd21597934935968a51b774efbdb82000619e86773e34b94d9e97cf56b124255a266;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf20bec2d5ec51c07399a249a88baa0e4a8d3c893459529a0f1a6d761a0b7919eafd58691;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8717d90fe07308483bb4fecc9e117488e15f7a32eb91183c42ce493f222952357e5eb12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h287032ad00ab421d2ef2a025ef31a28cdedb15b82bb9bf56ac6fc2b32cd5bc5f0bd70368;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1d4e8996365a5829cbc394eedf64b98da2c680ffaac3cacfbe5afda867d433cb545b76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d432893a86a810c271a85295556daf7c392824a4fd27da2b049f3940e7c19ebc7171aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39df8f0dca326e42614c4499598fc735de2db8e134a7643883ee66495b463531d5d6feb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd1fad1f0dc709a0f33ab90d3a40a759038b461751720b226d95713acc6bd4ccdd5423f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b6c464c7b1d4a056ccfd6d7cc9cb6d0e9918eb0629adfce47fdc7ac8a0716ccb9495295;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb47c49571eb6cf8dcb78889f95fa11c48bf8f85583400301a9ad3f765c2a27f3a34aa4ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cc97b79f6949f0890a64fb4b6c9b4ce8a532bec2c4e455536ef8b5c3728cf29ef4e6b9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee962e666b1889d634bee1ab663c44ac533bfcb31462b5e649283b2e4cc2d9837920f216;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1226cda52c43b17f49350cf5ea134596dae373e9ca081fdd6ad516d7cba9e3a49eaee7206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106a6880664a5908d971eff1414cf15a6353f2b8af9f1a28e1841d3edcc67b033c6d162df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50b6304e2632c004c64ff6f860bb4971290b52b625e096f0660c8cd003ac8e29429e75dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88b9bbebeb078d7b49c0e7ba2cf16a180249e5de68a5d70e74bca08754860f891cbbd2e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c2f0c951482c56c45d503d0d5cb7c5be8c75bd0c874501ceac934f7fc14a52fe63bb046;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb84d0b8e32675bbc0f9b62c7a84fc01c609ce61f68b2e008954cca7775df620863e981ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3aa07e54604184ed0b64ee5518045d7ac8f0e4318ad7bdb8aa2b5d2425286a55955d15cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9cb45dfd94fb790af795e6343400430c1e75c3608edff9db5f2381d0e0143bb9254a5367;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac836308005cffd4c5303d6e8736c4b467a85e042fb70678140d819e7a4104f08ead1921;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca766f184a60aea6ca80fbe7675cb9af74765e1b96105edfde378cf25896545f559ec486;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h335284e77a689a4e610f1c3609de4169a1237e0cb8a282371eface8aeaecb8d2b28459;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c646291db7c74d2407561069536ac9c5bc3d7d93efc65f1fb9dcb2f8b8c964360c77c92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1a1c428f0174d15021061db2154d3dbffc8b1a3ced5dad6907a3c5b2e55793ff61c8019;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a35fcb7ede684e2df26a073dc4c915847149c13be1977d7f95fcc1d91035730f3f095e75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6192ed827eff818fc30f18d5ee8f897136c88299b32bdc6a517a021628a5afc4ab053309;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5eb7b2b198a56871d48cffae1691f2f44e1667850d503ecaa350e514672222ea0fa52d23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48b42671d3716bc2cc6734aa5c3bed357b4806725a56e1488536bcdeae12214d41ddb75b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2d861bd3ade92acdd9ef067fa2b7930655ac8ca298b1008ffeea82c1af6bd6473d4f82d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1186a7c3e4afbfadee251910a1dbc45fdfedb2936b6e6bc461310bb872729fe6c6d0ebb61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8d75a9b3aef81f4c60974d1389c954a742db4b7d77fe9bbad592e8d40f66176588dc492;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd0a414e1a8e1a4496bb09d2b989ac07ee44edc77b2833782e5f44b871b8b5a81a0a3ef8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbee142c9978ac037603d7391200762836571a829b753fe51564bc8a7362a2668efd38a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3706c4c315f6a9085f1620aa9a553853ab44de5a3bdb4cd015baff672d329559f71a3943;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9430e97d93d9b121a2de991f4f0d71ad71f4149e2e0dca70b414238c611397189e8304f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f88381207f56307066b368a727928ca1cf763480e5bcc7c6433e085eb40f1f782ffe34de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5194c5f4e35268942246df7ab2c010e4d53ab183cb889c41f4d787d4b94046b0bbc42c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he36a82ab78a906a4939f2d2fb27d86abc2fd1f74ebb3118c4be25ac25da5e8e1291276bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca71440adef1ca632b81b0cbf4932b77d1c2de1a74c762b5e17f203cd72d6f87661856c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h994661e32b27ca68913fdc83c09bceb591bc32d15dfb8cf0f0eedcf52b6eadacc99750e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1348c22f3f846761ae121e587e6d92271b8cfce9ed1697e9efc66264f64bdfaa9b4f3f6f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b302c5a46e6c83fde5e1c4622075afd8657e95467ef3033133fe0941112bd4aca801124;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd014b37fc7a183c7475e466dd1e3165a4a7ac90a7602b1dba96c2348e1431485ff9ad012;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e14d2efb5246ea64a5ddf6df92d2bccc93ec71f67957b2bbce75f00795889d5722142ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8dd98424e64079922cb763237dc796a584af2bda7ab0218da3ec58ba3b7224a2bab9f467;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db65a2c1850033294ecc4740198b68f1d333088964765d7c94fa4c2787e9f8f16cc42c00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1295dec42105645138051ed88e1ce9cacb62c22403ba5239ce99a66f449e02e41c197735c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6013974a08c0cb793e776f17f0e23e91f94313870d2f9dbbe315522d171dc043f8436456;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112a2eba9cbdcb3c9608b5556eb1a78a9cd6dd420a9800734f4545124fb29a08a2ff9b0d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca359474da70f24fa5d16d41a8e4623dbf46c538d7d5f35da66ef92183a27737e546a76d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81d3664f7ac5099d20cd136b4218853c5294ad6dd04f7bb0dbfcaf2b43e8c797592266b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b668dc375a1c2b7033dc46287efd81a056bfceeb085a4c76e08137bec7056b4a251ffb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1bf33c691db2d959502c2ab9eb1c77086e6d0254c9c1bfbec11b4522b3444318bf9a55e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da1175491578c62239dacb34930c89e0070898bdadf3bdc092c5b0d16ef377110c58ec6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dab789607095ded37000726f9036d01c3e3e24b0e9fad47ea685861839a6fa6c6141aea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0c890c27b09b450e3f611b534ccc265d612bb35c09864876bf21f1690b8feddb2342c32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f987b0984c98a629aef86d6a7da5ca51d4f984408019321884fbeeb37b8168f9dc7d05e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h862356cb505eb2dd735e903d91bbf4e0dc190a56c6b3a682646387d4304d96160c582a98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147e5afdf468fefac26fdf920967d52cbfc3db2cc0a3bfd8b594bf2e6c9dc0c563db4e829;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d2853e9e86801cd98691d457af5eb37034ce09a894310962c279cdd6c59e7a0da5216d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a044c41942c35615a66017d4ae1b2970b8a8cb1c110085fd274ae6ef4fa81e579293f3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb5cdecdf36c30f9aa953e8bf43e611039f26f6e8ff1e2d594ca51d6d9b83dc0fcc76b19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h455672928b390e8cd26acd23d62be66b95c1053cc59f9fabfdae17e0447c58071fe78c3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11044aca122ae099cfcb94424df4b30521c2aa97f6572373b558e888135f2c6e6a1afe24d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba540a7f7371987f0f08cefa4c6e0d92825689a310f6c27db0fa4d66518d5cfe83e71362;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a76f5b9fc4ac2d25a7f8d3af1c1ca6b663b00324204333551269ec80520d37786a440a42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71eba7787da8d8851eeac49fa99d51c8305cd1171d839b552beb444b4524c580dda629aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8914962809129428e9e0461941acfe0dcd4c132f30d67566eca189b75656ac0d7b3fc50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f6abf70dbe290d8a7d7c99b056f9fde15bcc8ad006e1af1407ababa96dcf6eab9090f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc51c0e4cffb3af36692a69c676baa8e3b265cb21a832a08e1de807043dd13d31e2a16a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12232bee77f728e508e641c91b1845f07a3226172f4af9c844b01ae7e60190d2a302de36f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43c195fbab91fb763789acba962312ccf6151ecf07aafa4994cb6afeffd16165a5384d8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43b1d9c5f23115fbe5eca0e2b7220084a73ebd11ba368b59a07ea2400d7b9e03ba97dd99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135c4f9111b23e3cd729db26497181b539285d2140ea848f80eecbc31f3394b9dd6bb400c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150bf3282d0c42f5cde396854b9417d60324de1480044317d8617084e7875b828aef8f57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49d5bbe1534885acf155be275f44d5281fb63fbfa18740a3564c71e8d0c0a30775c61fed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1355bce0c5410d31262c257870dd32c3611b8170de64d19d06e640dd6a3d62c00f07d22c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d3158f74c152ff02778581ef695cc2a58c725a2aa2cec5b6ea250e26a38b9e88e2837b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32cad420b4ff4d268e35850590ea1cdb01d203108b0c08ee1e083b9f1d5b1643c856df10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc564d5fc94e6f3534fd3f18facf1b3978ec25ba0bc9bf534e34ae7a256ebc603942fc1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163d6cfefa9893f7738840aa90da4f2009c14b47808e7416e54f2dee632b869b9096d0423;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1291a99a442006504bd01d4c52679308b69ae74f33d1bd65e8881cb5448a114ce08fbbebe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da1f6c5d1a4d28e2a39c81bdf2fb8db6b1b97fa6ac0f252ee75fd05d3653aaf6ddfa3f3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a08de58bdc1509535d6eac33933ea14a8ee08eea4dc8f3115dfef42f8a4536af4ea5df6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6d98caa75de81ba1a69e313e33459abe361d459749f72b80306c7e3d0d189ec92d86ff4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6d129ce6d02cdd7d61a7384fafbb01fe786dd6f135f14f2cd0577da3c5b8075055d985c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38ad1222992d4f6cb497c6118ddff57e72dc5a5b0429b835afb495c8cc5080dee627b1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3d04e5416c1e3343d66ab959c7d9e9b660f9f8c19d3bba901a4f556fdbfbe2a41b0b052;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108bbb319c462fea3a9893312f304565f13a94b615c8c6152bc5b137c4de23f484fa793b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dff7b26f85745ebbeca43a5509c01b4e1537020fee97e36eb5f64aada4e08bb48ddfe588;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e8ce8dfca2a6b1b9b54fa50862def804fb283befb26429d348547004ca2f0d3e1c657fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff736217d2feb533b34427c833400d9347c8fb62e01e6b4b335cba3557cd57764fc60472;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h235ae014406d8ef7cad322bbe5e7b7b9b9d7b6dd3e4a4fa69e43823daa328a38429f93a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13616dcd6e11091cd5e280ac522989e984f913f70ba78907af77d088295f8e0d11fe2b78c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a9cc0457a0712d88febdeb991f6a81f80d3d36aff2596cf0e27092653ecd8ecd274cce3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13534f603d076e23dab6676968049cd26eb8b4c64d76e49fadd242c45d751076d611b5580;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb919f9271ee4273aa7691c7ba3f354b18b7368cd8ae691951c7cae89744b1d5141d54804;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1d39934193230ea41a8fd614cbbef4e4bec183819080f1ef1d1431e072fe3b114ab8da2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d71a161bd4198db9b43e55520920620d954d0bcd0cf1b52a77b9fa7cfd8a21ced158e14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a10d77977c6a03af7ca24e0072e66b0db31f00c9e277cc29143a05156291612b40da3a24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d413594ec8774151bd0e2bfa201a5f56d5a62082191d4e2cbb02cb2c61657a90c47b6b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84177621772dd6236e59cb229cd58d133e7e6d1428a98f2560289cc056d4d231bd36cc7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bdd19f42301f7917b6295e420207e45967199ec7a16640298269fc28d13a3fec166d81d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9240f4fafc138221ae137db579d370ae8cbf14197caa7731f6ab54255b2a24ddf4351859;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1d5529700d9dbf52ca90b82195d0465f42d23a09bc847ee8b8cd3fd43a534ab8519423;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc4065ef6c0c84528ecb53767515f8f6dcbb8955649d5289c8ad4035186f1b0febdf70e7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3d0e57a3ba30dca08943c2d4adebdb3e505bdcd1ac33fbd142e9570dc9218f5b5e52bc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h473044628dab8b0e94d91d0b3205d8d2e411a27111ccd17fac9699612eccb9a4e91e41b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cfdf9707d645d02c6b2ca02a7f4a806f13440e1bb15691b9eb71d9db3b723cd0631b0a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1670dd0f1ee7719ac787660138b26d9b1d876d54eca9eb21813af1b358c02812fd0070881;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fffdad82b9a349c4314a9b773850c962afa571315688b969a0acf6281a45e7c16ce47c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1858418b9389261140d0e9c2643bc5e3e756c425f3e9d80ba8ebf2b38b7828682cd9e34b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8fb78f5350e1c2a8935d9af4cb0888bbfe3d32df2f04a1a8fd1f9f7f977ebcf110abfb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafc7c518cedcdcb60a7146f33371a043cf9a6bf4dbb0dfa5f6b7d2dcd49ab3abacba62c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1359f0772db78963a8721d2ef87c5423145346df57338248c0a092893d2a40404711a62f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cc8439019965d9de1baad55a7cd6be4c27f8881a5ee061e5befc84cf949e11da847cf1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143a584e8a805cdb60c4a2becf98a387ad258bfee4fdcf82879b331e4e547d272d2c32c91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2e00d9c89c27d4597cdcdf8bee31ff40760abd5fc530b2f02e6225a03875f2c193300e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2491aec6178897ea6223d07544e0f599bd8d68d9e14acdc787f1ac7cf1cf5cc72f7dbc59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcda13fca722faf8662d5aac535a7f8d2452af11a38da865d453eed8f48a89a70b4b39a4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d19e11654966cb5e062ab416f450cce94c0504286f1898a40f69ee8c0470f3646fcf03cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9296bac6303a0592b5f4bcc2e37478bea808ad42188fc03632968d69ebd951324542e32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3e385a9b38174e16a2a6e006ac1fc45bde89384b13d842c1c788e50c67209b744c9ba1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab38e92742ff20e1dc05442aabdf39c6846b7bcbaaa9ce4766afe2eef3b6cf04a1bd7bf0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42caac7c6299ed8d1aabf844cc3062e169337d4d2318aa8ef2b8ce2c1f43b72b2d03121c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b267b8a62a9dacd5d6179192b69633e1930d3e3bdb542029c8be76287dab0b9cf04b642;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc92df03b87449f21cae79e54988387d9804d70faf3084274171d0c4160de181323d0d7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f6a9c07fd6a44179062ae6d7a09760a2f8b61079b1c8d5b6a56565b36c040885616c352;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9011ba24546dda66ac03ed3f35aa98b44bf6a90949976333a351030bf4df471e8fe4e630;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb35e994549c8733573fe5c40cd7f49613519ae039e5c995e50a252362e1552fd9325f091;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190f369a6b12829b0ce8b8a5d91b58c7b063c0245cb5c0a797f79e24e28c90ff2b94977e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb2bd4ac06204e68e39b2d16799ac356fd44bfb3a431fc11645dcf328a8ef738f237b827;
        #1
        $finish();
    end
endmodule
