module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [27:0] src29;
    reg [26:0] src30;
    reg [25:0] src31;
    reg [24:0] src32;
    reg [23:0] src33;
    reg [22:0] src34;
    reg [21:0] src35;
    reg [20:0] src36;
    reg [19:0] src37;
    reg [18:0] src38;
    reg [17:0] src39;
    reg [16:0] src40;
    reg [15:0] src41;
    reg [14:0] src42;
    reg [13:0] src43;
    reg [12:0] src44;
    reg [11:0] src45;
    reg [10:0] src46;
    reg [9:0] src47;
    reg [8:0] src48;
    reg [7:0] src49;
    reg [6:0] src50;
    reg [5:0] src51;
    reg [4:0] src52;
    reg [3:0] src53;
    reg [2:0] src54;
    reg [1:0] src55;
    reg [0:0] src56;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [57:0] srcsum;
    wire [57:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3])<<53) + ((src54[0] + src54[1] + src54[2])<<54) + ((src55[0] + src55[1])<<55) + ((src56[0])<<56);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194454d6ee9bdd5f7b9b41811aa61bd1e35513b32c9e5ed6949620df95f22eefb701522a73be7f676735cd3cffb3bd83c2738bc25c36a76963a1220783b2b11d1be89dce02295bfcd53ba15b997922fc267beb11af6d6de4345232a52730ce38c9af6ef2f681d27b951;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a1fcf3ca8c70f9af6f20e427cd7f6517ac597d38d2440e3d4e8904ae3cc45f523054ee3a3b8c8bf6ac2ae6253a20bfc713e42e354cc933e2cd83fee178cc5ad4970b9975de08674792b2c94bb8601ce7176a0fcc72006e3315145934c4b7601eebcc2c088208bad39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c66c433c4d7c6007de405f8e25a59aa51129b367074490db95be84fbcd99e48acb28c1c490ec8dfcf157e9d230e88abc878426f02590c6d9a154ad85aab602c1fe2f54500af3410277b60a633ceec197ef98355508c05947e8d73f73f4a55c82d47b3c98a8bd015fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dda9f8ec5d546da1411b656d1ad823eaadf49f7f752ea29e65a014aea52e1eeeb7949e406646a3a19d742b8b817724c863c25078b6a2a7f6d323bf8b0122b755df81b1a88295e49a24bf203da985995a3aacb889f962ea16fea543c1b748070abf90b1da11f970a07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177fa06046a1fc404e00ce73933fc843149090b561c5fa2968cf247f42dbef327cc7f00bf18e61f3442c6a2b21706383f5290526c81493015505c62dc717e725a1f037bee24e46be89a2b780449abadcffc20ff0d706509ecdd5aff96cc8a0c8a107c795b7ae1d8489e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3d33cb449417b167d7873a455a3a6465a37a0c5a4016930368cd3861f2b942dce231f71131ff93c2e151646d0f2b1b09cb2b15011fbeade749dc0058945dd1aa7647f75784c4946849d8232541307ad3edbbb5746e11f899a849d8a3c896b72e005f1f57665df841a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1893ae3750088fe5e41bdccf07d0c84a4441dccc0f25b7c71019d4727cd7e16efbf602058a902aa37a2005b507e75d176f403b59b0bc615346465aea698d771541328334a4af8929c7211af83fb7405e94c338ef55dd5758b45b033e12c56e71c06c31f0b2b3b85873a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f874f6ef993a2b4f4cf1f8008870ebd37c804aadc93db30637680cdd906b62f620a251020fc5bef67e16c75a9287aaefd423d7cd5e6edcc78f178f63ad3de0dd9e20158ea563ee2d5eaa6e0ea8d36ad9a02c0971efec0bd28aaf9b95d86fb51356b26d0f2137973a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75b22bc29957cc0598d9f452356a54a40f7254600a84d0acf35f4376db9d1e6967180eebd29c32558da4579ba5c9f1ec7ca4e22a9a359236ca27af2baf43fc7bba8717f643e8abc88ed3dbe5a7ae0c69b84c2b1fbaf4c6dbe12e0d8b06b7b7a751c117e4f40a4350d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1995b7b291590e2194fd5c76e368b00a5a7f65e7cfd29c3b8f278bf9248faf015d09d09e96851d3c908cdb17d32284944c4c55344da10d531e212aa4abdbc82fa132cbb3954203e74f7be193f412d0537b4eb6d87c8a319b5d5b9abe54983fe4396986832dc890b9456;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185b10a3dda8835873ab1c56dbede8ec84457f97da64a560001684a8610397ff8f36c6d091666d593efc4a98dd193050abbbf4f218cf5d59e0b8a72385008096fed40a3a604048a18f66e496f39eb3d2bdba48bfa539ac879e2b67fa5af8608f360f758173ac5be2bd8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbcfc549fad734d3297dce845c37af302fdfa49a53a122c97203fbbbe06f00acd6eed5731f2fb80344abcc2d496feeed03a263a6f8e83c3a7c38abf793babc5dd4922b1fed8f5f033e6e0e8798954865d17ff195f194f3c43d95e5e49b59399c992c47127e8b96d279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26516acdd637d2e561eb098581f7ceb614fa307ac01d628ba4d1a160c4f79e80a97859cf377d523a9c2efdc6c44e238875c736de6a2814fbd59294876bb30f8a0cf85487af486b519c23618fa1d92a5dfce8c1dd947bacc930a0cf6ac17dde571f40d6875aaf4df36d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b01422cb1a4b16890965881ee3cf58e6b638a635215a2261d625d7a19a0e816a86716535e7a93ccf8d71224f813ee01d3511146507d1ad8cf3c74f4a2ae3a390a508ca214deda829b643c45085bada51ff07507acd9ead0b7944bbb32ea9aecd495545591de47b8f60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80adb2f3bf974e81d469cd046d3c06564719903d64d411e6ed2cc02b728e7fcdbfa08b997eaf789c194b65ea6692c32105ecb98cf22c2eb792b17bed32e03cd773363f3331b269ce5c460ea67da94764a395fd5a34ad99de4903469b356b3e22978bb08f4781fcee26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha923ba7c0d7ae00a132f0999adbe664026eeb13b850b78de06da5d1333ec9df36b67465bab700d952a75d592a42464569fcd2663c67e57017928626da86a762fdc53d67fb90874ab89b078e6f94a6b5a54e7d7b0b3d5d0c17b827241dc2e554e4bd859b15cb498d839;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6232e0c027d735ff8ad9e261b9bb9abea71a289d99bb1f0269498799c9d88fda318533e73c0bf034d97cd084ecbc5d743b9a29c0686e5802ad8cbab4fc36c8dad91b7e8481108f14a38ba79db27181335201e38bae0d438f27a650eccb70bde6c8054e15cb4b87ef98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c2aa334b71a163329ae6ba43c462637e24d42712c35cd626476715ff6f196c874a9ca58b862c9479cfa96669a47f57e5eb378ef45ff3d613b173f0f744f3541bc5e128da09c37ce7bdc5a1201f4e9856a45ebec06e57502d350587e7e274b6d4a804babd0f8d392b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177f42900380c434b0fb75df76b35d61a4e9e51c8938199adc457d09fba58e264725aa4e2868ae75f39cd3bde9d1359019488bb209f6361956cd4895f031d9c3538191ded9a4a5cc49a2d485118f743d14bdae3f1a37bf0b0d654eb31554890500fb6a408fe27c73071;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dafe2d6da9700ef2c69d2cbf750932a264f2793e99c70a6f59892b304f169105e8c5f54db91694f9f7f4f35d4e565622407f24c2916c8b6ee637556fb8715be477f561e234d572caea2f76c9066aa47d7fa0b4143048ce63b896cec28414b7cb67ee120f1ffc9f60d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f67f9b0a4547c44000eb54f1ca82b843b1ab77d2a4d155d91672893de954a45502ab43efc40c70b8b580d295d46d8a62160123cc504cc9d2b9980df0659221b6e2a0c6f5b3e2e42130aa25bca1358d26e8ae59d46bc18633f15d613515c07c7b89c72d4ca597e72c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec86df1c2f8f037acc955239a2d851a3079da57240f33aac6c05412a7c50539f4b80790a66531c74dd8061b360e172f27fde65d7b47fff96f58d97b786387b6799bc66a69149cdd5c99f622dc4cd5a6b98579e9fa28b73d15f12c08393794215c9fff807c9a5bf000d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b0d5d227b7fb0ee27cc8b1eba30174a6e785b62c89b2b1f41a8735457c544bab6ffcec49c68b883c1871fe84b60f36525398da567284c153aca3fd9192ad64902b86077db4c8deb05be1de090245c54d404d3ab50461efa28f379878b79393f8d6a84a03eeb96aaee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb512e6aeda6c9eb910404c99128e1851bd3c07088ce4b326d117c06397615970ae1538346e5d782fe38e171bad48b935ed4f171af46d6cb426150f28cfa458961c44d046cbea0087576209f3319707a23aefeb4c8cceddbbf7c6bf9bdf6f3be1830cc69a299f41e3d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12041aeb2e4fd2da0f96d1b47974c7a31191a93e3fa0af17373d41c05586a984ed2747cee31a0f59f33a8afbac0ec0a73f8fa0099bd3bbea3a1d730a49234ba2dbb6ff077159e3d05d2c6778e8a68edd106c8f7bab56a16568980f3212c459dcdd3e49cfee68356039c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a8038feab5a4fd6aff1025dff540a23ecbfc24e8e925d8900a4281a212c508b628e94a68dd471514a93211e65a8e5f947358a4aaef0b8d7496d04bd848942b0f96a4465aff341ea473458b839f6b885b59a25245520305286b9dcc077bcc02ced751c387fb9f547af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb1d811a05609bbe7ca641ee5673c78b7dc89e210d4a6e6c267b8e9ba225819082eeb6dec285b4b671eb2fc40b11ecce3997cb9866755db221965932888420ed82c876db896bcc1d297653a742574fa61c519b4173040dc5a163ba085e78f4f70218d8e5d0a01e886c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7005ce79aaa19d9fc84d1e1cb2866900b9b03bc418db859b12897c54e50494b2a6db3b4167daf665b1c12c857ce07dccbab5fa4065c26148027d7580ad7b0510d5c6ec04e16c4ca15c3c7e559a8ceaf4301a3c7da61cc32120c4e9ece27abaa1a9cd49a5843c9239;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40c85d5654b81cc0cf602a3fba0dcb40d1f1784ee386545e30c552a0956f40274b002efe544925b870b70fc5a2f5776f61792205b9bdac5315a8f182460db56d8b9b35ef9238c8655499ba87732b37ee4f94a688f7f60c3f198bc2eb9dd80bae138789a594ce1972e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de23e3eabb5ac78436cc33c7c5fdc1b042c65dd5ad2283691a894ed116708fc1c471802538e29ccf3088af87b9c42d70030012f2c1e8af530afdf0fa6b58ae5d5c84c1ff0cbc6cf007e613f07669f363bcc5a561dea3b68e4df9cf4840f126a23bdc8978b0c5652bb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd4c843e4c2289e80ba49b7c1280541a058191dbc1e1d714e29611b5c3e0b8ad279ee1dc5ca7184f5ad2a534135e8a94c3df275fa2f64423bd41acc2aefdd0c53eb2195f86b609dde96e78b5ae3e84405cd84df4e0f04c5ba268756e80551eaffa06aeb029d9d9eff4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1657f92107b37b47b2a4050c31b8b7983f05663e820f67f14a55b692fbaacc3a7a74e9f4d01948ff6f19bcb49ea442fb9c2d94c202f096b7b0b24481a1ff66101e847d12c36629b151f2b74174306d21a19e268312101875339d90068dc712dca701e35b178fc8ce8c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1650a99cb157144f06936b703bc6003d1ba488e11fa5791114aa191dd735dea9a7ed71662a46b8af8195a3ed3588f6a33026a3780f42df16c95f1d9d389f4638b178ae0e8b478bd061a3284a265629ee9776b2fc90c4f63ea4a231a6be3d1458c599de8b1674bad4e94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1719d26cb49a3c370588cf89a3dc93adce5ef1c392b1f4843e8dcd92203bef4cec3f01ba34e24a6d327dee6bb9fe8d69cc653ebb3684056b49dfc13c8b241de3dd3a515d9fb0a67c12b5a87978447dd5b5ac9f80f6190b0a901ceb4be11d680d9bcd4f8da34f62eb0ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h983ff45cb17d58c751a66d24329348a6fc65de65e92f4945a5a6adb830c2ec3c76fc3c8724e5b5de3facd8c5538e94b25598e126101c0411d9f4a137df751a2cb93802227dceba6f3666017fba7892123717ca17c57c2b80535a33d76bc278b90f8cf0f2229d06115a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8d911adfadb44504329f56bb063d9d0ba877d33ff97124dea0b0856a41c7364556c3dca4124e2d269929b3452a1b3217c4a8c9553296fd493d397fb24cd2707ef2d6150e8a3784e11b0df62bb421e394c0841dc595838ab9a1cf43c1a74beafaf723f98243825a562;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108278855abb09fc795ded024f398cce023e2a99012f6071de6d69efbb44740316555411627d80071768b1275dedb67b751eef3e747051077a9b0b77965fdb7e8999e459d6ae69d1c8b63163a7ed43cc8f20e830eff14bf40cafee2c2b307b89962b1dae7527eb66110;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1762fa1e1386b5caf84050d1425339c9c729f6c73f47bfe97cc52477d4fb66319e15da77ce262d8e428f2f8f17a51656f9a612b2d468b83b50c4155fc1b23bc15efb026add1cc85e3916a6fa48ca414a520cb7345e3804cb38c9de216b7a6d8fb3ed6862444281f96af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f71e28835fbf5b42959526704bba5f346dccedbec11502054721a9aee8412c8c5f6dbaeb15cfd7fb7e84c5db820e2cc842feb1240f8a18f0fe2691ca5da97c84b1198a7ed689c04ecac94d7513b5c2bfa0a4bc814929f386e1823042c15805097ea98bba0c833d9376;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7585e3c5c3159e2de5fcc03d9e6003850a291725f249215efffd289236c8eb3974f07c8ebe67f91919335d484a9e6879defed3b69404875355b4f0e5600d7362083c684273316f2d9b589bcd8919b34d37985a4ab56df7d8c2c84bc491270ca95dbf96df724115ad12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c6d66d6e4f639cd6b70211a9d3a7f619026295a5419009c2f136854ac6b7899fcabdebc2ad8b79d854c029192b4a2eedd5575703fa9c6e2f6021f30bb32491bc473b53e7e44187e3e84ef57f532c7198eb148c3464247f05855acdbade67a3e6d86ca36e12db25d7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a590d7de0a6560fad9adb41ad7be06337fbf8d0b7ee9d39eaa89dce9d17389dcad3811b0cdc9b9fe7061a10228b2cb67ed5fa9a577b4ffce240a38a72da4788bab04f51d75e1efa4adbabfebb3ba49fb21a75d50e74574b3b3cd301f6b2b81dfbbe2e7cb52775c230;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d96c21a6cfe8bc38533942185b08adc2c3400b873d15355d9eeb181bf9adaeff271a27c55dbad4f77cc8d7de473761eb6a05fb3f1a4155c815fc5445b0ba56b04ced2afd4068c81c561a37dc5b32568594fd4cc3a51613fba858982d44ad340ea6533810fa7be75e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5d3e95c7b2a76996352f3936820b7b54a7b46fa3d80d45f03a554c356ff5c152af50098bbe8bdae25135e7936dd676be956b6a0ed084368b98276f722a5c7c8d4e2f0b40ec7085d30994b8b17977cf84a88f7fb890c7e56280b8e05734afab5388562d4e01915cf7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e28a65d2c90fef5b8db2eb11ffaa7683406a9228f3ce02cca752451a39e80ab87b98d10566bb0176cffeb92dd73a355fd28e2219276e519cf9c37380ab4d062f502e45f3df8d8ee236711ae742943410215ea0b18c5aeab0fae5a7a8eeae0379674df45ec9935a910d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f0b822322d5be1c33a76f82d207a8ad24b59c7c236c4aeb147a32d60434c9ac1a29346a06ad67ff675f5b0572efcc353717c75ad81d97b1a47459fb0e0f6c8ce01e80ca74f6e876ce552548a793f7c18a06e314675ad0c27684beb0ae40596a56fd6ad364abed33bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afd0461d24c4ede37e489b98b79f42b252ea9bfedf6302109a6b48fb1ac7b77e716393ac86d89d33aecfb121c8ebe41cefc8df8887fe59c73a721dcd2c0a1002c8606788afdca88775fc3faaa243f4723a35203cdca651bb7a96fcb321e878dea23337e59421551366;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f862476299d39a1d414b5f9f0f19802970b40407251fc853c19471590175fe06e907782a4346ff6eb4f8cee76cc238b10e2c10a3fe0ef2d84c2fd2964f91c407d170626a2613c8d43db74db9a79806a07c90f40178b95a415dd5c3fd58dd43480314e83829cc85eebc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7aac220971b8d13f3f39abcf685a771ca2dfefba82b839a68a6333fbebeb0bf79d474a0ffbf4ffa6391cce546a5420c20b445a4dd2d9c88fa946847d8338ca48798a7704f5db4f56afdb3b943cf07f310a15c0bf34215313d7e047cf310c847070712d28f5f1cb320f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a269c4c4b71ba9dc6f83cc65626060b8872e48885a940bdb2f2f85f9d7cd79d3393c30b48b34db2eecfa8cdd0c7dcbb2a21bcc7f0c93307baf467aa7003ce8e26e2269895c67166e9a95ddbc9f5ab24e7d0da083b6243759aa1fb4dc835f95b2b3daefc021f57877a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h873a1d5f8e88317dc61f2eb736c27f284ac3bc9656b134d67d3ebae4b508fa1d18ba3d931a23048e3f12262072a07fbabc8106c60e2cdb34ea537d8f2bf2af978d1f5d8d772d70173274c042f169a404dc3ec6e6d103973e497150076c509e06739181e3d4142df084;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd84a1f197997bf4073d4b8f8f5a7d297285a48013123d085ed9cf28c4bf96336f385075f0079033d089ed882d095816e82fcbceebf0f245126f81d7769eeaa3948f0f82b5e3ccd4fd82e3142a29e9af4c25a1e5dd11efa368ce8ec20bb6498ec86fab799427e68ec28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1838c80bdbccccdd6edd945089275bf4fe2816aae6be6525b4637589812333b3fd4927abd0180f2dff3302d45107e4b7a3baaa7dce971a7fe266cb97e5ace0335fde188bd55a7f50896ad29613b20f375a12b8ce06dfac8adf45203cf87f944946839a0adf4e391ff3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9abf863f37174b7cda88f887fe146233329df3bc5b4015e109672f650207dc12e69ee6d9821be9e950c093b4396cba02cb4eaf4ac973d6413bd450ddbe7421570593739eb6c680ea91d5d5177bd38db5fde38dbd9f00da353c33db848cf0425c3e58657bd5d6e25f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1203599d62e3c7da514fd95e542cdd4229597810510cd3dd099ceb2181e2990c2e4d03926a55b315188e490c965d785651f1be3a448acda00ca2700e1227c162812308147f307518c86d9494de3eb7e73e2e1b527226b5c7e1c060d59ba7da791fcac19ad69e955062;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19967f66bb14d29ec43657cc873158ce8af3d5c743cd6b3414600c98fd1f4c1cfe6123eebb9faf2c1598e841dfbb4abe4523c43b0d168c575999188334507009138bffd4755c615cbf16451f6dbf03954f396b425313a9ddf2bbd2c688da9e51d019ae9584e0c1cc0b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h958430f2369ae99225ce4771384e94497079ecde2c9454a2c0dc36bd94118fc5ceeb0422628655922b4c0499bfa9b1a357b275f096b18d4dd359117b7e5ddc850e01b6ad2c7317775eb3d4476db3fad373a5d549a8dc216af4ef98110d8aab776e914e18b44f34a742;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb09b1d194b8f87e2569d6e4248225474afd3585f8ecd1823e79f99678e1f77160ea0806d0a6f0fd9a330f4d6b89bc1583e80eff01a7985268b2b6eb9d33f7d96cf54ef2aa25db2b17a922bde61de179d2dc6c64bd001428fba3a3d1de7c87dce7ed762cbd391993c5d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c9466e0b1acdca0e11b798b24e3b6b8dbbfe4649eecea2d62ac55f863e3bdfe9dc0181077496326debfd176995ca9c4003acb4f532e05bbf88abdbb0ce2f47c9e5c7c83e1e18a1ce08af90c550c7bd3fe2d28ee2e5dc4e6402f13310cf844dae56d6b0d414b87a5fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134e52ab44528ccf1762d72c87e590406048a23120e833d4d17f2f7ded9fed35f147730caf1bd23b25717e0b6c3a5e2568c8375dd0766cbb554f000563477c2819b2dec2ecd9fe91ef1c68eabbd6637b19228b7ddda4ce31978f4c5dbdf57b29b2f6193b27be9e03d82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h724f8ff6111e0cdcd5caf700aea54a317cd3954f076a89002a81b6c5eb26eb36b73f8e44f6a7bfac0346c324092795738d7391e1e2c9feba4f3342f238365fedd5f204350f4dcb8916f5e6e88256201249c8c733449f76a8fab7648c5aac6ff68a8af7fb6c5390a110;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186058f2b1420eaa150f0b4961e1cdd42be1a9de7fd264817fc1616d5d93d1d61ad05a647dc846e741f95a5894ba7a0e1a4dba88789c8b7babfbd3e8da7a2c2f10ae6d73e147d4a04f89e24969a9407a4542211a0d037c629c83a1c22bc3d831bfc3a55c4be504d1661;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41eb63ab53bf4138a7d7fd736695d7aa4332a23ead769757b065de8bc32ae513a4efecd054fc0ea9a00f8829ddf5bca101ea585f1dda95a417bbb2f923dcfb304657676f490959d2889efdbf3d8fe893b572cf479ec78f5e51a4b9769b20dd1abb4d10daa804b54bbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb0f91a9c29e32e546845b0ac9796a59caa49ead381fa0a2d067a891de02df5f71f220bb4a82700468e5c5b3b12c625eb8efe6c2a9a0a8aa32e2f46bee85832e72edb45c36e08b7d2842e89add367980993f43bf180a539968ed67d912672d4ef8c0b2545a17290f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46c3bba6fa955bfd9d51d7fb1076862053814f753dafc2f91db80c4442b9b9ab33958cfb3e4048e1ae37316b5325560c3a0772809b06405ed17aa491ac62c24e6c5a4f56bf13e5121de4b7708e7a2cd4e799fe0cbbaed2273f09c3198b3930a498dfad66ef2aff4660;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198b4b565dcf21324e93c76473fb8050510dfcaa1cd8f2f7377cc7c0670113efd3dc202710fc7d8dc736e5bca81cc6a7dd41cd07bf5844c4a779f0bcbb302d5bb6b82a89eaeecb495b7a7ad8f7dda82c956954a6e16664be9c1721c75a6228b669fc1f69c7f4cf46dbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83ee361bcc8157a11f5d9f4d2ef633845acc56902d297700caea214572177e45eec222ecf9882bc4fefdbe1a26b47873c8f1e6b7e2843e9dfd70a66d31833216ca4a9afa20eaa74ff62bb6ac13bb5f898972263c7145c0397fe1a0c21b13cc04013799c28a29b1306d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7f991832e527df2edcd8ead4fbd9a2861cd9f8db0e4ea03c2bbdd07f14ccf150eef8f35d116983592e08bb37d289a7953b562a37e10212235b147d6a29a2aa40d095d40bfbb83f6515dea1c17953fa0998cf1252a3c1a4d2efa0819b9af2ed69099884865124c3509;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0a111b7eab84e5251713fccfb1db1fbe1711bfbcd55d2a53532581ca476ee87b8155b23d7fd51da58b0b205c7d8f2faddb46d8c0736af5af82e2984fc89a17bdb97ecddc3d1776db1087a4d306e2f15b644dfdead67ec6a0f046789b09b792d8404cc7f58d284279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10478c8a4bd4d8a0070bd94db7886be07db884f93f31406719ca44575cdcf4a67409ceef673a97668e9a1747ecb01c89200453d0250f04ad297eb61bfc279a92921a8c9cbf5a81c22377253986247a6d65d8f5414e1eded6dc9f29ccbc8de8c404a39f1e5cebbd4bb18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cde609d91d82bba7707452d1f64883f866e14b2b2e4bf1d4227d893fb2354889907cc7849285247193c63a8b7d47fc5f187c69619159a6b3f11ba77f3a9a42b66b6c6c367f6af59b1db8e8ec63bdd796914aa143f93466698eab058f0f56de8368e0ca58478113234;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57d4e69d93aa4fd925faa5eb49169ab43657455d95cb7731519edd1a9c76e6fd4963a1632bb06119574725b56bba7a46f6f46a2c4f9e1ff734285604e8c837942cf265985da43996c227d723dbf60457a9956f5e9fba142ab9646d6152aaad311d9c2c048283d63b6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a0be927c6ef1e877c9d9b60f7c5e3cb9b08f6388ed1957fed189bb48237ddffaa5b5eff03eded66c3ffc5bd89d7b8b62078ae2fbd3018ea89579dfff1539379d0d9ea40582518f0c6a3c3351f4caac9078c38767cb38d21daa06da5b1517284565eab3bd4d3067b3f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b810e04fd96055ad3d326d083de3abf57f61d0177cc5bc45ccb08270a6738b053e7317b2ff56c220832d6c74c572557cf43741bbe51757e09cec84000e9738be2bc8f1ddc8ac014b2ab2b9f54b85c3dc888ac3198cdc546f39ab4a06641a188db38400d1ea22de679;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ccde39d08a72e6eb83b856f882dc2747696fbc92dca219f02d61ee64c16850580d4fade82e78c259082b5b74207b37ae9adbeb26829ac6db1483f31fa6d14ee29ca2391bb30c7415418810860ff019e1fa73c6e515140e1493fbcc6b63ab00d33cd7d4dc47d7450fd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e134348e458f3eefe8700b51aeb4d3c08cda022f8ec1c3c36d428b616210fe2cf1b8fe43575f44f1b7cb652481fab9e8e138dfbadf4c6b2131812c5587dabfc8bd4c6a261a7429f0def239aafc089546a5095a255f2fca22a4f2258862a162b813aca083e2720a304;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa7d6f30e0415b06de3dea248e0e172bdb2e2cfaca3db0c5244354582fe782d3a931f4c81cf7137a8d91c9188a00c5bf46a938cf9a9fb1f9b6f7adcd41eadf84668f0709de8316290ad083a9ae5250a36109e5b92d458ee7ab2dc6724617698ecf11374cee5dd3a59c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f9d41dbd5e2c9649423f2e4f243271f2c3cbdfa497a0b5be36d2472797e68f46954278a414692eb0e3c7719a63536c212aa0cd956bb3e7759677c1220fa8508e6235767631675ff24a23ec8f79a84ec9348a45f69e7dea498ac39fe939947f3dddf8989c95378064e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28ed2c2ab5504a410a8be1d7413bdfe6579a4bb8c4763796e02b2d5e8313e7c936ced233cc53a43d263e874e587962ef946e7dd74d779ddd35f0832160f30e38c7f5d6b15947b79ea22f6faa26610d260a571f083a9d3752458be83c6ee8066106f8a3023b3f07bda1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1413895f8c751238bbfb10fe54cd69e20d64c7dc977e268aee353cab622ae9069a33c59031650f96a648d826ef88913c73400944c1544db238fe49dc99d961a482a1845d5da8dcad95bb0075f1a2e6cf62c40d4525ed0b5f8fadc15d0956f4714417fb93ecb3a78acc8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h37290697af59a1901fdb6300255a4be7a1997d4727f725b1e6b6a80a68932194770290c18f970916e2c0eaa759a4fb8a56a51845bb0a0aa3b71be60164a66c0e232deaa4c89ed47c5a9b41f8bac45e9e8129f7aab750bbbaee8321c93a4933ab04f4dd8824be5a7574;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2a92634ed876fee94e9ee249d9e418ed37e3922afd871d305f3a6d55b11e1038c376427f7ed1dcb1ff6cfb8f2e0f0c69e7238d535852bc77e236f608054f1dc63f1394d2d954d5d5cd596be2db9331ee8f10e95dc0fc2ed1cc55ea6a52bbe81f060c219135d012e9c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0474978b24344085301126b3fbf0cb6d7f0b5252b9a4b25f6361a6e23f763b42e9ba47b700b9e44f79307a37792c8d32d2bb1bd3820e284d83ce1ec8af069e2983e3d8658054a833bf5a569e4060c1f021ef0d6f46a94cc3257c4cb4b75f1b9de98972a48b6b58b80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12134708ac9c998fb332beb9a3b5ddf99a17439df0fed412c5c342a4e92ca78efa50a91c6af3a17ec6db1ca489d36b04a16b04776d864dd8d4d74da3bdf7bbd49a7efc88a7292fa3b4308e771bedf824e0e8e56c25196280d8592c60ab53b2ffd79175cca6779d91bf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebade160b5fcef3fe4f52a68b81fde2f318ea36471236cc635e75eff796d1864fe7cb6e83c05e7c5ecfc64abcb6621df52bb1df6a12013666f7a47db05c92509caf01e8677585f3b5e3aa61b453814c68b36250d146c1b281e7414cc89cd6f1e73da998fca35bcc65b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ac3306a207318844e8669bb2a0e236d22eb9b4164ff04d9a8e6689450cf35b634200ab17b81ef35390e7c35a031894ad80064f0c6e0fd2f3041d05e5ebd9f814d55a13d8ffa3c4774f6316c348ad160c115ca4f32e5181bc1bba155d8b7f579541d85e362fbea2857;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d2c3656953817d0eed85df9e03d9da2847818dc59ce482140eb4b2a8b9f7698e4b6ae0a653f4e1b7ed36f264fa0b96ba39dc7a78c652bae25364a85a00b1dcd78d448369acf185db36366d099899500edd043676273014b6eba4f33c1578b936f4017a998d6df0fb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b1fbfbb89a5c5899e11b77ff858a159a43aad239cb465dcb9628681f490b88782c9f4f1a39d8f8d5ff1e5a247e81197f9fbac9d4fdb0d6ba1b5b5bfdf1618ee41c14c4cea30786f226cf585c721d3dc43b10ef380b5a71df6e663c4109808b21c1eeb0c22a3abc219;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a90bfcde9666ee5eaefaa0397263a33b77422f59695e54ce52546fb0ec732be20542ed0048550c7e9e4582f6aa63f1c9bc9acda6e49460fb5c0af392c27b8bcb7fcace34a273a87678a7557a1e4a4459aa4c87e50daf3a7b90e6fc7b97a1b421c2df7359e13aec5a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1293f23be951eb2d4314934df15015dca7a7d3e891d38749d54e3715f78512d54729a54bccfd35126265e0808308f64bb1ed5be40789e1de141a267ecbf446c987bf4756775cc40840e3b41c35252e279062dfd4e6ca1d457f834d437a0bd85908cc4adb719d2ab60ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aad42ac848e586a18bbfb5f9f275268b1dd374230eeb3a48eaf07b902293621ef3ce5b890b70bf5562bdfa45cf76138be94d185e4379d82d07b1adf3646622f2e655e26ecffcef8c2c6a2646630c5d899a224e4db09584769910de51752f66024e9af921eeb59b9812;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95e7d93daca044587fb62bbe7f42b824348924a041947852d22f435ea95a9cbf18496bb70725f67894c036b6bf2a9ca54d701ec3c8f0399a6c1855ffe6319398bc76664805d37ed92fb677fb9fe107b3404781913ea1c20c2342112c466cb035f7ec3130028206b86f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf7c9ae1acfe6d08664b30765b49546f30c1a36d8797918cc278c7a011cd717c363b5ee991ec44b82f5b8bd80ab34c39c849c915ab67e96dbe24170de6861ad26c9526fe0fb5c337c8262ae736eaed1f78e96ebd8b45b6c784eb6f410cbd080bf13c84a3d07584ebee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdae6a4ef078d69ba771d48ec6643b38f2736ada0abdc61158363c38aceaec7b2a1207bc64df76de821bb2e429a964f1fabd0fd3d0157776f18a7e5fd8ee51f58f2b7c9c43a38e23315ed8d06c261986165e3b65003610c61d2e8fd00153be65233672606c83b22b043;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16aecc4d38c7f60b9be739bab59a33274dcae777c57040cf0b3a4e6b5528b9e65bdc70ce340f4ffec23b3d9f55694fbab212988ba72d1cc33fb1af1d3612bbb4dcb119b60416db8113c773573bd2bf531ab635f47ab05894b4041cfb45c0fa201575a2a6f410178c0b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77c97e90dc6cb9e343229abacda76bcfe630bd0872c9abb0e239c1f40c176bcfe5d684405e83223a02265b90e156842a97e9eacadcadf7dbd71dfaa7504f6e1c7c5537c5452aa4d7340d1fd4ba7469be89c29c317665f62b4933447e7c09b6da862c631f7abc77efab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc3ea9b6a2a776d049ff9ab28f95877aa8c6791afc2d6bb14ec182c7cc86742e7fd2f6335765757317986e7f70ee3e8e507148c752834137997d1c35bd24f3f5ade89e916b97ef8cf1fa84dbfcb9dc43bb6b55df95aa7debae92f264557ba2e42d250210a1884f0ca1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121887730e8a1911e045efe1c4e7ac02e4e929212e91aed3b2cb41be4f4f6e8e7105bfc77f378044127dfa6e8469a0f7756baafc6d0faa3dba001eff2d1efba7b0f489ae54cdb7a646aa3288d7252ff4c85ed8929d3c9cc3cd3cf64f3e72401945723c8f13ea9cb3683;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdad3fb0dc4c6e8b4c56791a83808a2bbc1e9ce96ce91bcc5457e8492cb8310e67d108d52e55e1acfb748df6b02ff7236cd2e077d98759849ec7ec6ca006003f666238a50dbf6f846cb4a3d49760beae757f1bf1a34f323e8be100ce2e9c39b443d5a8326434810510;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da8b0d70f90e5ac189f63a756e1b1615dbef6a1d99689be87f03a3f04f595046f0e3ae367e62ac8048c5f87a4da82a6d49d3f7f0e27f1e1a96bf67b45f6aa18bd13a104eee5f93812dc0008a62706fba48bc1c96f7b2a818070762e89e7e6e52f3fd701c94d1677fc5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec1f1eba8001da0cab7ae191a9cf0365cde9bdce59553aac44c78791902d7cc1938e71945c43da7aa53988a2669825fb639c69024bdefa528765c5ac9f15a707325b4906761c0a6b50bd13e2c4ce4025e53e6550d14a3ada31d324a2fe40a57b50cf0b8dd2cbd37c42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1928a4b0323c0a82d7784fe294e88c4936e87d546f9d8d0418f8e2ebb0b8963ca4600e912c574ad5007661c3e8c46b700dd11aa787eed19749163cdc46c292e4a1ddb44ae9b41e0d46ea4412bfa24a5af7671a06736d59508db86e912ac81fd8ad8f7d7760785fe42c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ff23988b112be7443664c91b8484bae4199da472f59782a02f4c0b4e55a5696ac5d01bac3166cbae534f942bb6d3a2155dd8f76c55f0266544e3ef713411890bb2c236d99a229f4408522e5eb8c5b8aaf478c3b4d8a83a6021f93a35d0d7d9da2f42cd0e8dd9c28b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101c239a1ab9cfd052f65f992264117c3a01488a0a5b289bdf12603486ae4e94b716c7a686ee2d4baa0842d03d23d61d22ff488dde7ab89187291142ecdfab3e3bcb9d6f8be30aeedae4fbc8ffb384e2a68fbcd289aa2ec122d65a44dd0232689fc066f3b109bc902b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cacac7645f0e1e8ad333ec48537a93fbf9a74846f57723302526629dbd9c2c21a13aa3d7735e9e1b3de800ca23e5c83925891c96b64ed4e1145342452e9537dfce8d6e5bbb248f34dd17cb166d11b35ea97b8374421791cef82806fd452c663779fa3efa28efad53d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f5e7c8d3f3a96f49356007497bc7cc3a6a7c651c4ee1c14ca37a88eacaa367392d80f186601e23047e74a5ca6502b0e33a102489f6e6531a1a851c963df9dd0ef216fab8b9ea4b6346c5bea36a91a6efaf7d1c68411c4499720b7d0bd991204d6da04c64c7f2af4c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de95c80af6ce4c656a7b6f9c3d6ed71f205ef990774c932156866b9ef9d3a993a53dcf2810707a686fcc03233efc59f7e4a80da959bc309ef66c8da976fecbf24bcb899974fa2bf22dcfdf2c714c79840f1d1ad956fdd5a8dfb2b35a04cc2a8a8d2b3165810523e0de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d8e5594d6ee908e1303158b10399e7ed481d92da45c40cfd7d89dafdec606f12bd1aa97ce9d96c5c5d8f243a66fcddb3ab5a06d3119eb5a1c8554743c1c2c9e852b8a4a783e7a96492f8d5dd385c07418129ca353d59ceb628da12203bc9e93ce9cfa6e023f86a07a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f02a8a4f227114486a78dc6a607113d79b74f39d64b047087bea3e94a03f4a1be36215f8310809fc66642e252b64f331fbeeaca9b24de7942b2d499299b561887a6d6cd953487f932123c0f01ff3f550b24d2071f475d1d826afa36433d02ad8905e0c29c912d06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8ffb0401b35da90dcee9337a6104c3c0c812796a9fc5aa86d003bee986dba915349b8d73febad0360bec9e43d85bd4bbeb12be473977dbbf9d71f317d1af52c45d0d34a1e2db9d35f99366fb4394b0f3a7ba149357216e867726a124438237aaea447ae17bb3e0070;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13bcae6e63b0543ce055d55854e71f3b60c33c3309a3708a70621c41395da54a8ebf75436d48d587b6e92c374d5da3fe3868bd5e2780bca0c0a877bf8fde3957782c1893a3a135d190878185fe97e09e02d458c4c753cb95ed72c20e9aa0fb54f754ddddcd53111ba26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4bc975313a2e74e16162bfd178e00f77de442c98e5ac0422cd31487904a03275a5a7c563d6f01b04ac8283161e61a17fadbe7baf6e5c42e1c7c4819b7cec1956325cb5bf461b670bde83ed1756c7f5d4e9ede1a3d7b7f42bc93e7aa9317c6e6f22274c58e5a0e884;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152df1c818f3f37109b7048b7eff9b4a248c0cc908c18a0c79d1b5a34e1f531bfdc6cb8cc0d1d6bc3d22bb4320049584de1ee2d2415e662100014130bcd173bb5067e74a286b0413c18683505152d853759a56243b096bd6c63db4b0fe58d5be727f21c551c9b3fa4dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e90480ae4212fe37e772bd6b7d8dd6656e52efff956cd5661e8d0b42535e4ecdbb64152423ea483b67787f0ee7ee6f7c8accd0f1fc4acb48a2a5b72aec6b264dc7a062f6c81be4b9e713261ecced63e068c0f727d7f507b6d133c24657f36a66d8df3a03d56266fa3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6ccdee565cf258ddefea1cac5179aafec14b446a83fbf6baa2ef56d92bcd734507f3460e360986868d00dd3c5e66db68ef943660faecf0d649b6827f521cce0c59be69c415dbae9f235b4d3db836e1ec874133c1d67f7afb9d439df8d08518a96542c535809bfa351;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c265cce42e56b8657427c5e61745dfd29654173128ad8acd2c4dbc2b08c9abb831838bd1ce7f5fb6a096eaa0b5a5b0a42704c20bce78f4d7d517ac00ee08f591e2e0febadb6298d49c83964445f9da3e4281af0270ef57d3bda9cdcc95a1f2080beb431c83001cda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff8f7b2390bc23e3ac4f893a26d1e09613d9511b0e6b3766b1e3974c6b4c3f1ccf24943f6195535f299e8d8cf0bc569a1f0bd5ccc25e1634bbcfd52538f3cb6069059e99f3dc9c14ee167b5aff97b3ea98c20c3fcf06228a5ef6e62e62d40319585b226964e4d18927;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbd932aa5b510a72e20ad00bdba9d528cfeca9f05c52c4b4c3c12fac507e2e65edb224c6633d98c30e725c8d61aa62a6ec2c91d0a4def0080739b19eb876d2b657814d08bb62939210c311efb893ef552c73e55c9c7bd9cea3464b03e0e15217c610c7ba528b4ebef2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8405c3644ea955b3dc309b8d82319a109aa058943dd2d28598f4557868a43a9e12243d47d09974944f4c8dcde62a7a190cde4dd9d08a18d9dcdb93bab52d32551df48bbc4754b8af7bba6a6e0b3e9c7a214e2b25ce6ccda318a02c3f7150571699ce1aed1dc483f8d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7e23778d1c8a4910c91f2e05475a6b77fcb5b880505c68fefa076951affb1c3eeb41d8472769251c3d46d0019d0749a5706741ec58b8037f7b3ba5ed41d8d4b78714b0b8c678763f72a416096218b5d62becadd80c0210a365042a47e43d0760763d20a811137cbef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd07c0a947af28ab8f196d7e720508c0631ec931b0906f27aee5eb75d61da185e65cf1454c7bde57d12b83a60445cf1afa58415078c3d2997ec91154bb324ccb2143591f8d06915f4320c1d8729d21c44970c8e1cc26f90cfbd5ce11f9bf045dc87f20c29085ba86df0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c50acea7477123abf07337c23930cccf02f74f43706c6d26b259f03bbb8d04eb9bf74cb29690b738b83a9ac8ed1e0cd378e977031059b018e16de8825725508e0048dc8fdc09366ec44e5380ecc67e20f02a98d5f27a18d4ba83621e0b9c69671753e933d813bf5f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19077da7571855d4768e92797d3647e05c1c012acc52c91a55dd2396d54b798a9f584b2f8fec924df81e1c9cf654f33d2990acdf1bc41b5386eb733f6fa0fa7991f53c2441c4197409ec5f4fc7c091f5a91882483d13be757846afae9ebc17443fe237f25716bcfe220;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha47fedc3a5cc6d9bd171692d2b404b459c659b90eba982af51631632c8df27fc06e882a93f8958b2807f37e55683c76214892aa1ea480e6e43533daa58c039b6feffb7d7fc9bd23c86fbf02033f24d1b489e1132655698d6ef4f79c540b6a9682fa3f330a07fdebb60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab185efb3267dd5f3c619bf3a4c40bee039b5c202837215e14de332d50379edcdffaaa9d3846d160db77d28a873939acc69a66daad97a0dc8c7a5535876cc0320c846dac96ceb26cbc22b91655fcb6d66154fe72ddab25b3b181118aedaf2cb6e6319bcc0d9c9b6893;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6dcff6cd43572d8c5b8c3ce793b8fad79b38585ad0de11da14a832876c691c471c34a48f2143c1c1f762340c2583e584ce0c328534acf8051508a458ebb061e1a03efb4ae9d7575962a8241a331999c0ec61af7c6f516ca84ce5f7c4b6ac5cb8594d91438a1676c05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d038ed77d7c9d340dad188bbc41ecd4bebc881a54c79c1d7c275e29c284d302eecb34febedff6b59e2d757504f034355c3343a2f5e32d57b7e20d11d9e536f81caa4fbdd5c7176b16eda4440d9a33ffe652a6a0db2b580cdff5108f161a0ec0ba74f4f64fafb73149;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fade8da646a608f3928a451626b21fce2af51f105d9daa9eb654ce2620e0857721c70983c3b428f358f2a8fa79155d18b6ec4ff180f51b0173237b6be990e203389dd0e93d317e044d6343da9b64d2b09b70640cd6a3374c4ee246e1c36664dfbff6856f9c66b4ec2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b287c22dae23bbd3cf5b23a3179e1182c96ab0ec186ef68e162d3a1a9b99ab87f4e047260b12bc4b943a5020070fd24c9d4958923cd4866ba4955b959f100ebd3cbd4faa3bdbfcb5add0c397cb6ce94dfc450a1677375a721b9bfa7c0b8f35f949b44f3f6bbba82d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2f92f81ddb2471b92ba5993cc8b1d0d7a53a55ff48bc6ded7a318617ec6ae9f33f7328295f7fe8a715acc5101fccd5df619af497517aa964e7c4b30c2ebc78c49a2963f894371a770a3e7157d6b2dc8a8232b0c8680b93609bcd8ebb0b97c87779425ca4e1a22673b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1845a9cd732e101707cb3a2e8262349019662dc05878a771ad4af87b57053719db4a50d2299d5aad8435744f3f79e80672905dfb506eb21a6da55537b648e1f7dcf930c0190420af03d476bb9c029086b3fb3e6ac760fb3bb46ba41f14b5fca48423dc4d0c9a9c0aa97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99965d1d851c49a4be646a1a79c0aa705947c644c6bcae4195ddcd1ea1fb1ed056226b331c74d0714ab17ab9537cd748b472e310fa627612f521ed504c8d8db0f2fefafe9f7ce272d9226e1e74a8b713ea62bb57ce7451b4a8198c5e8377cd043186dbf474e647d2de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d3ec7701d910a3480449d27dbe4604291e57ce0396f58b01fa0a8a84c79e66bfd634baae65a04ac4f1969d5bcb4556015534357876212bf42e6cd6bc84d0b98e254531a09cbb4b1fdfe6eeeb932237b51634b7ee2f3a9b0ffcbdc1b87398bc6557e3dca99db5482b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b0d47033dad4e5d4de8a38d4265982391314676e5d6218fbd49c84919cd2c8a510b88708c6e40fa1dab999d24889f998ab4d0e8f167ae546a72961abce7f10da8121b1e6863acbde4b753f4496b8ce32bbe51b609d24da556929f535bd98dac19241f603c74080d72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d24613b6586ee73c98671674f57ef8a8a3aa73b64a0617c3eeffb5c867b536d1c3b282bf25f7abcb6ad64eb3387077ed554e10460bbaa4071e388991e8c069214b2de51e40fad7073d9df46349db14cbfe3d16a6454660b74907f01839fafab1d6c4ff9cc72f00531;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184a95e9461c5eb5ba42b4dae0e7edaba15bad228c4f12b902b54edd145d249b994d9863f6f6cb7c8c77b6113be9f6c2b31ddeb48a3a3d0ba35afa1b95bd074332aa44344e241e4c90b7fb6d7827ee41800ee6a874e57d0787dfd4af51b901c152a9a4548cca1079970;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95e233c65ef0e35a3230e7e82c959ca83795b56f8d1dfa3da9ca044a8e31ab3d91f19651780c10f6e9d899f4425142ac0293e8d6c6139a2cd56b1fff28d0a3cdf8517d349e382692faea7ce70c06c32d0785ef3d4a675f6aec74af29986822e49137f591f7153d18ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc93d96fe99e2e84da7b5ce05daf0983ce9b1e1ad19d9b28a8139feff26fa533bff6797b03cff25bb5bf65e3ff51a2578cc373cb7894bf0b0fcf76b8f76e5172b31350000657a05189464d50c24fe3a8e4bf7af058b9520da4f1fdaa5570653ca6692e7c83e70fae970;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb32b526a7f8798ceae38633586f3ad3871a8b37666ebbbf8cfeda6ea17f75734db64bdd53bf930ecd671aa09d4acd3885423a877ac20afd7dfa117f1f0c457275f9852d4e82831f327cab1bd704810bb9d78eb4897a37cd776da4a5f78d8357cf96aa55fcf8de6fa46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be81738743a01e44d311c9bf469eab1086c196e820361bebaf4b74925906098a09e9f23029b36fb32c78380d0cb084b36cc424e3f6f4ce634ccb2509a43c585f5655ffff702e25b914f0cee5447ea88b570e85c5f2a7bad1e9e3b1ab7b1ef6f766478479b9568d0b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c166845fcec53202960025caabe44d70faf54657f6d0873e2113c843f1396574a376d5825f63b25156415a66252af9e0cbb8c64d0e91143921a758347689cc13b49b80acc6a224d4cbe251da3b3d5c633ed2c56d801b0849e433074e7d2fec9a1e7dc05ae186c4535;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5b530b6aedce91482da05ac013b2e50dbfcf261e24fe91f76f9b6d6a9cdc06760bc5528d98d2606a979370ee05ab0ece8c44d80db633150922455550119e7c3399d43c0a096cf2b5ce04662c79c661ffdc190cc1519ef5620d8ea45d9a52f7f8f253e17d49652c15a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he97a082cfd93d6d91e494ffaae62078afd2301b9ccefbc6862e7098eddb95ac98218c965dcd22f5dd160c05c4d7374ddf5892eea73c882597620f7575ee99dbede6c818f9dd5825b0671592badc640e3a9b6ff680cd0bf84da6a9c58baf7acccf420467fbbdb78a812;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bde43ce00f78e0a5471d450908fd3a38ab0a1ae878ee260d87db549fa807c7ed241206afd531c9fd482d4702cfc77ac1c29d4629634cb9cbb7a4d6a3a843d33344a4fe5bac6a434c830b2f1ce91096c7afff902c2484365a97cd4c436d23c1ecd7303adbcd0468ee7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f4f016ab1997142669baaaba7407abc50edd67e092a24203dc4521f4c14e0bb21436d561740cbad9cc50187f0b718edece0679cd8385c4aef41ac40527e2656a7bd56c6bd389f19fe5f2ddaef40f4a44838295317f23f50dbfcfd6712619e5ff0248e38022e6c109f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175ac21735572c1dba16dbc8cc6d11815cd75c543549c547f16feaea75e60f6a3d44f9e1901e97939da41e91e339e305aaa5454b57ea435e49fba02aeb0cd157b58b867b2e2459c50e1e3fb5c98ca5b3164a7202be867da50ac09b649fc670a45cc49a4bbb56f9b7279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121a467faed3a68e6d048486b4af650bd077905ad63d5ae158cee77843f688dc04a0ee2de5b4cedc7bc6c1d08e2435c99eaff7c4e04b423104470afc24e60e5024603702a3d4802d4ec8ba27f9aaff0669bc9b4fc78a1f5c05e3b099686fc9d72e08fe542fa24b98d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14178fcc32930b779de9964a4ea0061a62fc36f7fa7157b20d87f7fee7f41852f3cc1dbfc196bc97634a7b4f4ee9a4e7c1d433a2c53d89e0825283d63f2add766b5d8ecde801f60f8d116ea84274b3631274cba047b9c9e040e97604870e90ccadfca0cdc79cf0b641b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150e66d23cc6e8dbf1ff3b15d62ba134678c0b642809c3fdc4a22555b3fc86980d83f684b54ca9ef4d014e1366d72d354b8d31db1ae7c06a958c1360f43402ab695c1aa96c2c4217d229ded533bf17d7b73694ef6d742db2eb24f0bbf2872888e630207b79a7cdfd6b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f8b2f887b902b7171d6bf4f254c83b65d1ff8644b1bd6d667d72c198e069717966403d9e8b701a603f3825013ea0ef986d9bf73184d353c9e3e4e3b59c6f49123e43aa128d73a6319449e9ca7876fb8e3452a3f8eeb5f117e073043ed5dae600fcebd22388d1b35bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1170bb68c91f63757450244b946341085006100edf61b97acc730b92526ef32af32dfd68740f6fb2af94fe855549fbc666dceaf7ddbe5be073a464c61a07d3e9b01925a1029bbd90c5dd8d0a774d46d9e0e907a062650c4f01e80d0596c0c8835158ce8d557fdb2dc50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129974ba4b404e6a6824fb9481607629b015aa12e659400552a713b896154beacf157f282f747a2c768540889171da3500257a0fa332e6cd4bc091ea781db11130a7bf35b63b6ea1327f3f3e03f54ba16aeb91365196a376fd24c384728e302ae982471a1ebd13aca58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3860ce0f53bc184c267ca4c6a14cbe4bbd046755f0546738ccffd37be37834f09fb0896065816635ed0861cf1bfaee5e4f74c0f190e959839fff6571b4f6b5e892992bf5d3bd08836ed9220dbcd0b0610fd71a21f04cfafe1b7125845b48524a2acb74bfd6df54ee5d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc2c12420b3dca3a07f4a874fbdf929523024ec336886386b5e5be02aa6fc01a29ed105f9fc197fe9222b1582ee6e3b55a0a7fca8166f38a31a588ea18313f2a0b736ef668925026403ce7efcffbb428f2929de3be7c69df6334ad6eedbf754022782083fd2ba0d9db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c059b630d1aa58c5c0032803a4f02ec67ed96746cd78af8f8bc89c6941f21326d0a45385dcebea8e814e79253aa39f56635d0f98445bad4483dafc77b794fbfdb405c026a61372805dca1df56301622216d8a6a52522fa9342e03e2676c837e1fa1e40b0beb822c28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15003ccc4ef5eac5be5a98f0b3b2a94f9dee6372317988b19118dd4feb098454de78e0a2e2205816e5e9b2a8f7d86cd44a1ed85c517e6e176e4e23cf5248f4bf946d12bc05f4b1c5e5507c4790d05b6da51273d89bee649021145526cfc4b5356e9c20d58e8519d2d87;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155a2b39286223e1915326d1c1a1646d258e741597c2390b63a84f9ed4538476d6b3c808db679e7ec4f6c01c6bbdd68079af537001fffa5f0f7eb174b2b0755325499ed65a506209b7bf1aac7c5b22338610112418a7a3efb868f57d419b5d2fa6de06042744f09e87f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1277e2a51572e9a027eb4446ee451c11eb52f07f15c941633574f9681fb5a0c5f8534f09b07794f7186ca8e54d280dc02193a71f45cce7a0e5d166c847a41de32158400cf84ad7b60b5adc38e174c51d96c9b99548bf29bafb34b61d41912e47131eeb4d77103a0e4ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6c0dd2a3680c87cba010d24563569b3f7f28e890c883280eb89007f998dd2799344fdf08c0d35881289d8a9dc2c785514bc7912c0fd490ae2f8600638d53eb650f803e5ac0619c801535c3521ebeec11a603c88487aac9e43504414f2ca22a4ab16140d9c1c293ab4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf05124fbc5e12c0531fd87030bd5e7d489dd03aba23dc36db52fcb3c39ccc8406f2e2f8a9b6fb9094e0db96e0e680abd302423ee338bda9cba56ad70c0e32e4b243d4562642f4babe1a059c95a66e0aebbd98c3589cc6666edc8c72e027e2bcd1ccf40f9c9a856b9fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h442b8a6680dcb36791580935af6e709b9eab0544dc65eac6cb87f7764f877eba04017ca7ef23e1108e6f6ff5b85d82e04f6db90699c04853a09c202cecb59bde5df23401d2557c6a00f5e4a1131b3c182654e17862e99d10ee2490df4502c23526fc710188e47f0a49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15dfa0e39a547e16b0d9b4c433aa632603877f22d51f13cd194b9bf26fac58ba8d3b0281af2cbe61ba2f11ace264955fbe57b9f18ebd23ff6bd58bf342f972a895f37f0e9394112b5c835f2227beefd21bf7d6e9732ae5a19355b4a469f28898a24c30150483f4979b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f85cfa39da99982c65e9c82a7e48e6d52710937e9225e59fdf1bded8e3cf20b3a27ac9237c89a169f85376c404adac6f5816235b614fb1834077952ca96e70ee5f2d08cf922defe798a3f5316c4975b5b9ffbbeb83fa597a861334e9585dea5046ed1c69eded610996;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69c62c92b7fd855124e330b6962c11e28d426ca2215d21939ca39e8b13206c62e5dc8d6cca6076bef1734726984ce7b52f4bec4b23729080326b8c27157f52422fb1a4490162f07beb55beb371098722ce41d14b2e6976e19ade6800473ae10451e82d5d3b1734a599;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1473ceff13f0c0d8ebf2012a9a4659e1a5b3d52fda224ef96d24f85ecedf6485b9bada13f5606c8f9e0aac36e4890d8d83de8a01b67080f6f301a20f708c6c251e54aaa8a8dd58054d165f98aee923c1cc25e67ca451ccc2302eed6c82f5f9d99c1ca8bc7682cc8fb99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha75315678e7699fba8713d6792dea4c16be80ffd3121a34b824a9b8c09ca1c28fe36b63b581a5a945e8afbf1cbbe9aa540216ca848dc17399b1545654a99b59787f501597c2e835c5a457d7964683141fac3d13874040071203ca5dfaf725b5a8d6d8ed8a53a96a107;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h329644afa6751c97ca9ae96870c0f9d77fcffbf329f7778c1c7f5cfbc267610babdf7fc148c5ebfabe73b667376087b7458eff1290015d35605b711fc03d1dec95134ce7cc9e88d6272e35490479f6051f573b7a528f205f51e2562072d60b65f8517c40921cd065f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1538aa2a5183359455881836c140eadb1cc23dc4563ddfc7af73fe8c3314dbfc75ac18dd0479b1cc0331ce6df14fffacd0ee2c3bb5b3b8095acc547ccba533f6e0792d1ed598c12e6d619cbf1d0c8d116f3678eb12d815c54017f6f5467babc5d6f806bdf1d05faa410;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175d383f9879e48c0ab02db269649a153c72b3446fa4856c5b93935969887d0d312e7dfda898155604c4df451c270cef20cb73169a6e5819cab405af600b71f24b25dc6094131fccfc132cddbc481757ba275d217be7addebc5c2878e42fc7fd6394b993bb2936f5174;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de7a64bf953dbc007c0cdb6e8b718094e01fad634f13b081efbea96ef002b88315c5802e5e396fb98c50362a4f2a290f105b357a3157058af1c9c0998d05e6633edbc6c8293c14bec934c8efc4196fb6e047d1a6b3b038844d644d6903611dce48b4f6b4300b00b10d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d73bacc1624b58359338287f9f3836a79cb82b007040f6f25ddd4933fcfba053eff9d11d78b4fd4ea8c292ef20d92713c8fbbd11230e03a4b0c57395f2c85f1910c54889ab3de7110693f8c0da155a539c56d6c3b28ef1f0939165c19f4d6ba2954ef69bc7c288a38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1551092c37cf5a4f973f005cb07f49a8e57e78901ea559ff1023289ae009d74fc767107135938670a4bd9f5ac6b914c4d5baf47d82c0638b8070d10b157f3734bb7d5e47148e5a3da3e9bb2a06f6f59599c7ea3f0e405107e512799e614a8242252d9c5e20718219e4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127e5bb6fdc13c06d0d422de4b642c6a4bbc5f08ac8bda265e3bf0bc27f5b5f867db6838821aa4b1f1320ec1a18c54507f2a09bbaf872c85b134e30173aab2f54470b1a6aaaa8705deb8c3343f093ee13f734f1aeac5d5a09b0d0619ade0848224bfc7eddd654491bd7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb55c8108e38b6d5e58e677dfb3752abb035885cca9b15a66af4bec1fb18abd48086748705be536cc1202849ce6d20bbffbf4c660a9bc5ddf76b49a9f7ca500674a8f6f3d7b4d687f2b6ba16934a445f9f32b5a923cf83e2f6f023a81a446576be383bcaf68a90a05bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4b65bbe2c7601a36a245ad3720924548915ef6b58cbbf6b5ed935762c865a5cfb6294253e8796ceb9181c5211e41c75cebe4424c2f56ff89f078d74cefbbff3c6601abb88fe8e1a29252025b4572520353930c88628be915c7d18fb1f21248c912d91990f76ca4a11;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9cb097afae545604a5660687473ee678516ecd45ba2e28f6fa95ffb392c4428c2c41511248d80b1360f0096d83ccf0d41632ceef5e6b43e17f52b8368c32eb0a08b7f35284547e24c16055ed8b334291596a2ecfcbf16dd2f2ae6cf5a65c8b2692c651fe1a139735d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbaf40a8ae9bb02bddba6fc47603d2892a592b8dbee6001aeec3f7a1cc8662a9188dc1ebe600d0b4b1907f01f9c85a29cde0a48d5d35a9e65aa5caf00b4e52f72871b18784806a5eb44e6dcc960bc96f7e5db2c0bcdf0c7d5bf6375ac0cb6f8517001211737f025d7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c0d9d0d023c1087b7f0d8d910a129008e0934982e89f6340a747b1356c6c95ce54b186e57114f996295104f6040eb03383e9b4af0ecc4f97a5309572e0a2016d4cfa38d2f4b543b67a14d1cb3c01b790aa54de668c383cea4c1fcd35a90f54ffaa6f344238063c96b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11370040a5ea19812297c2d72cdb62b39497caaa21a41cb51915ff5b19d1c6ac5f17df9426c19965b85389ad58a54854cc9c09e9d8a5a1f9b34296591ee11aad4a8cc0dff46c2b93b381c411fc242f472dcf31a765cb34adfa81b33311c0a7e400d1d9c0b982d24873;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c2429aa9a558f64c656b02b004e1e8afeca494d019b9dc73f2953bbc31a5154f4bc642e308042c8d45b272a395563f27fb28d1ccde2e9e8f26a76498b0c5ccaf5ec1b57809636f5f715a24fe8245110f1bc514a3f33a7e04d12294683aa984d2a0aba7d7ff2cb8324;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h403e5a971a2f309344dd371556a3fd28330006d698c42a97ecae8fb6086d59aaa1784a3be22e25bb80006c21dbe6ad249808ce6a9569c4b71449c700a44887450b5dfd4aa83b325d975b26473aed389a88adb617d3a3b259ac61a9788a0e86650599cc79bb57e52451;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad5ac5322a01695e709437f19d09c86364f714ab55460cf36af5fd63b9936c11f1b8e16bdba86cf0ce3771da3b0dd93f6a60a0289319cef75bd3d33b732c7fa4510a975d62ad6646a4f502a4830a9c1b781c773832ff65a917198061559594f3c3ad13b32efca5151;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had52ce81385e0fd98a81159a57416a55f7f8a9fa183e0289cc3cf0a0bcceeddcf457d93eaa07e559d86cb7fa13b90904b59af8b501f979abb0a56e44ef14c5e1278fc0b4e61990e79861ec85e6b1541e84294b88af6443f968a6716f5f42309fb45a1574342575876;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16054c1f4c0551f9ba8c764ed11b0f36fb892759a54869c0155814378532a33cd661d766b25631cd6e3dfe8813e3e00ec1621604adbc4e3df44a9319d109a0108b59bc03c1555bb45602b57a7f757a9fd0bdcd6707dfef4393e4aa4cde146eb4146a4000b74851d1401;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b12c7e181f3998344919911bd4ecab068c3d197c1c764bd8a35ff4f8556b850e7277f31ebe90419b2c6a8f4a8a1ead4aae36aa5c4128ee534dd4a70bb06e1a62421adb9b0657405a4b1c9d5e570c04cd0167740a945b7e5f9288f7a0536810fd590df5ec723d4150e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7625f83b93cb7cec54068461808bd4091c523b1581ae471f9cb6a40a7663cf93266201c6a5ea05bfc356e0fb7d7ca7bfb9d7271ec0a5898466287749ac04231a538e4399a71aeda7efb358b3c69989efabeabc4d297e695ef920516ac942e4dd2e7d6250520ce4b96d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha827f0fa431a9aae9ca79dad7271252540cccb35d38cef93be0a035c96398fed1c7115dfdf5c3310d0dc50d3440273c42029252477d7e1c9d01a8a404a48a2885e27a8b64f3927100e433a896471403afd1f4db1c2e465073373515744faec10a0f31df5f2c47f75ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h24b1eb9df65e97582ee12c5f0630e788e50fc59edf3988fdf569cc879695bfe4615381b3b60052aa1b00f10e7f38599400b0948c61e2550bb803a7b75fd55183325b1b1012b86a80d491db27476d035b36852f2edb9d2c7399f492cdd219d79ac7fa975dace15705ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3744ba56f6f924bbc3601f2a7d8b4f8e69f0668df7ecfa3b5a8e9a920b2a4936a7ef6657a05b15e3f91d7e572b17a9fdf305405c94285cc40774f58f5a28338e8585f913ab15169adc2767b428809051a39d44ad7b7f7948d137983a96f25ed8a880fdeccbc8c1ec88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ba63dfff75a13702f40763019a85103641575058822134bc7229eef8824e5002efc91cf0f1373854a1b6e81e4ef16379ee7f5181b6bbb72610aaba579703458ad77a4629966c1ca50d10d72c2f2c827e0191821100283a738c92952b2ad15ed9912cb156ae93e2bd3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d6ed0e6660bd9d55383768572a5b8efda5b50204f4b73fe80d343c53662da56ce7d7090fa9d99fb13a9efefa4e8cf98a70ec6eefbcf0b3b0819b2f4c261124f49010a44d838e5a67670c74fcbc2b411684646e097827dac8cea8b7de9ec8d956194580278a4d1dcc9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1077a435c65938957c8e4a32c7a8f34848bd67b91f21094a8c3562fb8da04a68eff4f1e4b1488a7a08a00fc24f3ff3d1277e9b0131a590d5502d02365601f04bf27efcb795aba999bd7a07854915c134fe91711ab9a3550029c1053cb1d490c3aaeee76ac621206e6a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160e4c2f77f4ff97ec63606389863a8db28aac0e67bfe5e693b7d34e800885a0fcc3bbddd10191c163e247edfa77543074d9c2f7a76440614cd35274432900a3699df374abbc4915e57897583f2900335683e4c867321de2bc0e928ed3130b835362e3fbbead5d7bb75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa73b481f92dc79eee83a76fc33b6829e43d4cd3f387eb1f38fe1d5a98a55b8d17056965052aeb0e5f76878274c118c96c69ee671b31704c94909dfb4c02528032bf184ba65e9db72b077c7e6d2f5d3f74bd6676e776c60390eb88202c329b9b6811634f03509197bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8d726c802a68f95a1e411f4235458aff7eef20b2939cbee317dedd5c8074fcc5a88f467ef2e04bf094faa162f51923afa807d54272d6d1be368547d71640e535e733c094aecf38ec3a54e3702b79ee5777d88f7aca52de8e2c1473ee0f0a1d625039fb2e7c57c4a48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h347d12b9d1c168d9ee533d98aabe8e877b66f8f8d0ef8d3777f5b4a220ff5af802f3fe0e70dccb586e8f0fd8c3b69d089038b1a86f2e69263f12c5f2a15c5eeb43819943a55f88f93e7f121c86213d1833fba7e29ff5a3444a4146ed8d011d851c21dc7777fb3fb011;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b8aebf68ade9e4fb79ddb9c60f274d24654119a6231fcf6a44fa9ed83c89bdeb0c1270320c7a8272b228c201b49b2f01c9932b1a9c25a363df3453efcf86947ee99f8dd80f3c15faa709233a5defd9afadde52286bd5eea823071f57c7a2ac3610e13015496cb2be9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdb7731c16922d4eb7f077a318d4f9f35402facc7fbb4d5dda75c2d473c4d4440407fbb56fc3ea498a64fa9a94770d91f1619ed125cf48f6a9efb005471d9074dca4a28959cbd1efc809a7ac6e6dea6d9f40b161e00d11c085b61944c1c3fbf8a5942e2ff763da3639;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he64aadf20380e647ed89d901c5f00e97beaf2a6f129cc25289d32caa7e291e64d1b173338cda4a256fe23f9e88d747dc1e232bc9e6b90437b2d864c9921b61f1fd1fbb7e1f0c90795c5a4be55464fe147af4de93041791fbaabf2697da0a145be6583bf90419f35312;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a791870c3fb08b4cc83f1e723220cebe35cbf803bc33ef5a8d13812e9e531e7704ce8453176258cbcefa564eae2b3d2b4f202c85cd13568ecdf36d7778ef1049abc55aaf7fe30643a17e6cb16fd59f22e26b5322cdaa460f2956bf6371b5ef3088203ff807f63429a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156ff7395245fdbe514b15b22beefe191d817d897441b2b30382d1006aec940c3c904ba6fe68fc8b86b7262dda4d0555f32d540c8d59e06b662186fe34c2963142045d35860fb1c1a09553874b192f96b785f30c47f93f40119592496bbe77dfdb4e311360d1b87bbc2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101f49a9353a3293638b9b0e312904c25498751077d48a9330a60d8f7a02928ad6ed95b57fe386eb0f3b68d9f1796680ac2b01d525dc389cd7c3d1eb3de23f633eef3da16c0c0765e3173471eb57ee4be1cc13753a165009b7cb971fbd0e7a6c945ba1347b14449392a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee4d192acad320e04450cb0b9084076c4b3b44f8a2e92e45e48a1d3a05605ccc7ede9460935c51076c2c49b0b57dac05b22e3f0223f0da525ddd79e1809009fd21480f5c282a14618657c35f4d4aa3ff4793aa3ebacc340e4a35904d37263437c300a170beac843174;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2525962736d72c09afae3d374d0868e68859c8fe4aa2e79959638746cbfc8a54868213c3a39ee02ed48e279ca1d0d28797eacf4845c3ae30f28c38c8bdf6e8b4f2a11b6bee46cc2f4ee5185cdeb444e4297205016c3ad2782ab1fd4e26d1a3e279f0976fd8dd674c94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc01b0a5153f0e695544554a323b6108a1f003a30bbe205da01868d9ce42dba233c04c1db362ca3f4b31650f9824533d0318fa47cb9e8eb6e5e47157bb3537907abb97951deb7bf172f5bc16fa8dd3f79428a59b118985f5ee50caadeb7adbb27d05190e45790f784a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eddc5e0246c31581452977c1fce8ffefd48a1eff0904c52fc9b5cae026409a79e3224d8c57f5f2655cea8db9a084ce865aba25583a75841eb11d55d22e51a93b7fde49ceb110885dc6dc874c68f754e5042a52e1bc7943241f6ed67886810e7f821c35ee55cb43dec9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b02008f123ff8c85986f6e8516750ccbee0d90f10346acf6376f5fdde201e9cd95c1a3137d687debbf51764cac365574a9d5133b908bdfc28194a0c50b6fc20aeaa5824dcdbfdf6b1d2a1da168a4e488cbdae21e75098015c1f4f83ce8f4af456e52a4a062d2ac18d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183353a2dcb32518e6ec6e9ccc8a1e1840eadd5f0504c12bf4f29ede697f48839e4f7f09ff073cbe7fe9a517d6374084d35d5109c7f87593893a71019a113a90e8dd93253ff7d68cda2efdb431c1cea6d600060b078b9b4146889c57bd782c5dac025e7d4ac9f71f33d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f5c51b8f1038b45711e32224567dcb8419389b6267986b87d903bcbe8e907dc1dc1f0ae97568eebd20e8621415efe380cbb0b4006af8476ee6c9250ee62dafbd6aec521db7c9c2e64f08917772ad0cfa3faf0f8de33eb08431223204ef8718b089dd347d0a83ed80f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87f1cc0311d449200cca707a3652fda869245fe17677c337186a1477dce37b58b73d24efc4da37b09d895b0aab748ca0ccaebddc382fb1f6078d671a76d5c0de1362ad3b071816aa4792a5e78b71e96d3b0eedcbd78184232ad942aa787749f86990284c2c912de795;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162f75e347c759865d0168fdb9f2045853dd1b3cfc9fcd7feef2325efc6e13b445cfd385b8ee6cd309db500f5f11975670bd7f9776b9c0532f669a27b961331cbba5ef35b24df1dc75ed0da1d08ba24dd381b8ed60074f12875886cc08e028de9fb3c9a361fceac58da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c30323f5d75269dc24aa3856745f9ef2163540821030a5226de54eea84d6b1b23597ab345d118a0633fafafc9dbfa1c015b0d65262241da1f2a036410704b4cc670209b9e2b1e0a0078898826be8d33aa2c8c69b283413d2a2773b520958a16ac8951211d7bbce252;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd54dffbf4790d590cf50a73263362e4f74f85fe4c71c9c394f889eb18709a651a0d092292d27b77d9c1ce69352b4b1fc9fffe8e1fada0466ea3e4d20a235981a29b8db638c3ed98e660b2ddaa04f22d44c22847a3437c47b4ffad8903755b1a7fb1239e147bee337ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf196d9865161f79fc1886f8af8ebf0bcc5c8f28601ca29fcf5ac27542f20132e0555328be9e117d6cac97da4ce8c991cf0efad0856b18daaa8f0d323d8ff33e04c1b80517d83706083944efb89a36f3c53ad0148e78dfa36cce681b1611673274dd212415909368e8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1a24ba25ea8f675ae6b1d5b7b9c09f491aa3748f8722af638c9402018701e9ab385e847778edd7a8c98e943d26eb93895f412c6e499d93dcefd1a9fd26340b50e5bfe720f7e2ac88402845dbbb0ae0c2ee42a7c6aac80d8126f846ce3078a85b7ee6c5cd9e0b3a2c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a29496b13b837d05f3409bbab55ae0d8d86acd38bb27c6d2b52e61464549fad9cceeab657e16baa36723cb91f3fcaf72d20657de0b480705ec740efd2344e10d1d837dd2365318ff5991cf05df5b664be0303e0f2abb0842a566b9875b0902c4fe9e8ece729a2556a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9f8f9a8076c949041b38c707a0abf04138cff4c664175596caf94015906ba819ab44481b339e8e4bf0b70e7e358d945d25d944c5a2be8b0b14af7e39c6eaf56d614b6b15be204897d94244e9caea24a18f3f3f12bcb7c1dfa022c99ffdfb11f70395f51ed78cc91f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d435c1143f914502fe7f718df736b5fa922b67125cd21f51f6b2d689b17430d39404cf3a06181d4c9841b559a70e9c0c625539be4d2898e3feaf30e5cde20007c7a84c5ef466f4c3af9c580c765859d2d152e21fa50f4d3652a1aab90056788f317553786ce06db64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0e238dc91407493a8e6cf3f8dad79af63573ed5b44df86299375491389e77e500fdfb5696e492cdba370d72adb02a938aab078999ac45ab14c64769d33aedff06599fc0396a2af502c3c86e7e9516dfbb328471be089ad94e710a7eaa5ae8a7408a8c269f65be0402;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7d063c67ab6b55f08a6ce71dd9eb40613afb5b721495e73f5e6d2d43d2f7d26e6db44e446e7552ebdb75c3979c27ed6e45e03f97e94836ac57e6ce69fb064eea296ca0f17d94b7b8472e091f9699b8cb4fcfed35550a51b838bda05fdaa181ef477f1fb54a1060da8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ae2cfcdb56049294d01176bfc22d8e703c95e2f82ee626b24c3f535b3c73c61e48d068b206c265848a2833a839b0b57f94b5809c7afdb25df4d253930892ced3a09c5768530782e79c90c36283a269bbc8db277cedd44a6d63e21db07845d93a532aa6547a9582ee7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h790244adad0b8473051ddb59d9c7f0c457dec174ed9343d03f8c2d669c6138fac4015224b6639e497e2a7d44de5e1b2c7a59478801d43145fbea138e25b3463fa55007bf02a32eb26714996697a2fd2a556d5f8691c335c8895279b73e39dd1f683fde538de55b7aba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf15025e5f5e30bb2ccbbcbb0dcf02b89e946dc61a85e13dd96f9bf64cd45a6b23d40f5456b1793576e974de77b581200644b31d1fe473dc463716430f0803c1e8f02d33f9c34684e9ebdc18edf9cba85beb0f40570fb1a1ca38044e27758fed72d7cadb1d9a0f75602;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4cffd1d066f6050ac2d0ab7c945ab968a70197f80136a75096c07c3580b9219654dea39bd47d2285f45dfef42bed6f6d5518899edfea68ffceffece8994ce2142c3812c55da99b4b3fd756cce840789b236fdd569ea80eb890ab94e904fa7d8deddcf9f01f15720a3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h749cee5b67c007c159aa1c50180fdf3fc802f616919476628d8802599be2ca03e87ba450aa53e4f02c5e12f89c773c070a34b7aa1711797f9c11dcd29cfe5777da9a5508885a283b7bb9b51d5b3830ad05b887d86d8c5befdf4aec7fb2d02150c28af16099eebd7bce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9ba883df97f99822cceb6ba8af680140e4dfd310dab0f19923aa72e21b3ee38e8fdcb0d90c55f611a939df57365a3291c964102decfca9cb04ac2809eb5b8fde8a84e1425c0abf2409b5e15a3077c2bcef95914c8c803ec21f5d9c80ea24694ad05ee46fa72b26f09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h643028120f12fddcb500803fafa88cc06a5758ae37b7f9dff322d2bf2f65686948e6f0e33c13f9dd47002093c7d6468a2e7396003f030530ff838454fd77b453cd1598a6594cb57b9ba50667bb0c3ba3450d5ba5345a549f18470ad497ea50eb7b5ce68300430870d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h904d12e24fccc76684dcd81f162adb7f83d6ae4d0688cf806bcb1fda56e4f26e775a59ff919830de913631b7a7c89cfac33a468e561870e8cd0a39d28e88cf16ecd9d0b74184b13b11abd61d0f262a1a9ce72ff8907318e16c72d97f0c68ca5ec7a7613fbedd429c0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89668f4fffdab7ab7b5053d93f3208ebd4fd1ccd5cfec76a3d45c4310eefc559f1c0d44f4b34a82dd2d1d0940c6ea007d594dfa711223432f2b2cf70731153b20c5ee34a22a23f72f8f3c1b139918e8f3f0f65e8e924b5be523b16401fcaa0f0ee2739bfe7f940ab4f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0defb8bb673f62775231d36113378bc5e392415a13d4d49e0210fab1cfc6b3fa280c21f8c29ab52f7b262d36b2d19c6320cd2e323b9388741f894d5a6e1f7f155b1d0e42032ddd1826ab3c8c4f6e0f4eb0a4ffcdc23271fe5fdec10ed6ea2784d5fe545ec81cc15f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112471c2977b4c531b0077f813b708a3622bc22e1c8366a465f4f36b25804e083f878b6bfa6d50e0696b0a126498b15bb787e270bbb3046f44c6f34541d7ae6c3abcb3923f482e203900543a4e85fc5ba7cf12e46621a38f33fd01f94d152fe65a3870b67ee33ff01d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12eb2b6964774e878402259e60750207e3672384ddd9ba0fffea46e599de0bad96b3025e57cd4d73efb14b869799773cebd6321089e3f88383879b93e30a63349996d6a17c915c1e930fc337d06a7ed64a55782d49d627c57885926cc65abfea54228143b693e399959;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d79de144bed02d89f087661ca033e3df52ce57d969a0fa8d8f1660d34a9b8a22731cb7722c8c90dc10c636d7e507d59ab4c3d744037fa04580e3632ee8a7a97332db9116cb6e9106d43ad6d6f358b170fccd86cd789d386b8e9c4f1f7caee172d3fda1da98cad184d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7d43c82e11c7405c669af71d3744ba891a26084d5d8c0cd9bc6884da57915cbaabf715d8aa6466fb24dbf63d3e66b695968dc7e7399a80866c075647d7ab7af9a6a50faa147bdfd0759444f996f9c77dd725ae409199c9aa66bacf11922ec7aa7c9f12ee373b5cada;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfec9c7763eeb877d6f56444e578136725080b2be6bbe24071a3ab0f4c94f6d7f770fc071f78db1e88e4d8e9267d140f702bc8fe3378b6811c56c30f6f990af61326d6c7348f841e115ade7ff896bcf5c57c9cfaa162aa21bb762763390acaa66ab53d1277bccfe5e96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7783aebb24dc22189434db69ecc586004d01a5861ee082aee8c4bcbc710afe1fe5ce7adc3367055a3291ba148be8070d1757409982bd9e58f53835776808a8b626119dd22c0d5e2d70c0e1526d7a720d083fe4a77fb1309890164cc29c3973e1bbc1c3316b164af39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eff94f2a2d284f165cb0c59e92e8e41f40ae15c66c531f71dcc1c76b330c7943ecb502f96ea47cd7ef1b6645f35123a9c203ad4c0a375482a5cba6a224f4ddf9089d0ead47edb43c4d84504418cd0df0af506c6ccbbeedd86680536f1cc848a3d58da7866995c13a27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d479a31dbb64a7aee716c7103f4041155ee04c1cd2b77eabaa368a0a8dd0893f2a5274f6623002fd78e93135046e402fbb3310b8ad1bd8e4830a807cc0c26eb3fb24629fdc7533c604ee059938f47e56fb8b50a9003a8518c1475527c8ac9227e12fd11f05312362c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108b5c47a9c950a4642e4a9fb19030d8b03241fb7a3876ee003055045b2e04893cfd22467b6c994c366e23777772971051b22af86f699defd04107d7e23fbd2a7023ed82c845e5f1c12a7a8330892f860f646b252b6ae6be97a0fdebe68972a484b258c5a47d0bed18f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a5d915dc410ea6450ac9975b48d48753a7f8dc8c732743b06665a7e8a9459681a9d14bcd3cac3e6356c5c8d3dbe730be8588f66144a9e6bf62cbf96dc2b7011e082fd334e5cd34d00fe565c768e5a6b7b6483a23943ccea0c9079029cb75f0440456623f6ef62aac1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86e16c700aab0ec7b7218e057a892154cf4d18661cb68b0472ade138c106f590bbba77e3a16eb47eddef303e26447051388cb8fc4843483c5cd9a31c96dd4a7abec9010dd0f4635bb62b28396d9366aaecc1f8b9e3bee647d6abf88424b3e615f2678d98b913ab241e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ba3976f05382dbccd9315ba737356ecc884a4c5dae624cad9c6c81a9917249f15cb77192ca84940142b6fd91dda63fc8417a6a56be7204299b82a1969d31bc28068a784c874abddd0d6714d90d5042f8d6941d0be56025d20f57c1f3bf53c56e8348397f6a72857da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4773534f78d8812103a1c95a57e05c7a9520452582745078ac83fbe845e39dc8bf3b965baced660f5765ae9f2b9dea5ee66fd3f670994f8dbe409bd7747ce6d7e53040d168a4b90237c179819408e0633b55ca9f1c1c1c18b4e4e5fe35c2a744bc1d4c72e769ba784;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had7589db7ce6931d3af802b4b9f12395fdb3d52f7b114c514974245369b38c2d4a159c24db6b35d9464f6e3701722d24528f788d16077ac93f4817410006fec042dfd33009090d02b754fb85d9424816a3fce101077b223eeb83532f9c899f670068287a0dd3346aae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf68a0ac843512b98cfb86e45368d017ded25714cc80f561c899a28ee20c9b20c2a27c74f8ebf0e11034909fba616d35c22aa71cf28837a38ba2bd03725095e27c7b2ab416e51fe2d57e9429087859634c76c462384410897fac3c5788005c125de3d884e4d681339bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112efaef2e566391fef8cea7157a640c6ae91312dd28d0b56cdfdc2411d06baaf78d600ba3739b367918e817d8cd119e6d31e76c065a1c9baadd7ccd087522ca4a7dba5f7f0b6479362d237ee32b2f87ea5480f0695abf7bf6c01ebad8337606a07704360141a44585d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95318c04c10b99e769c4ae2da41ba1f360bf2087140854dd7121b8723fdbed4964aeefcf441830611543ab36a7830fdfd8409fff12cedfe89a2fc0b5fedaf41155897c0d43ab7dac5e7cc32d180aba55a1cf6f1c3f645c63e04116533fd45f232b1e8b3e4a869ed730;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5c816f7c4ee3cd20b4b49dfeea39340540f39225b39c8072491be203a05a6510da2a87e6df09591d24a58a27912d02bedb0fd5c76a2a48e17d0617feae458d02889447b25fc0af5a474456a9ad968aebc8c45a5856360d0bb1e33f6dd31593df296b247d4422bee4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1884e43eec8f78351776d560eb69f7118fb3b9f5e28e5e0f7782e2574ce6f8a1660a6b343d6cca30785d1aa25d785e88901ad26622eb511795d8e7e87671ee357701b25ba3459c320b3a78ed8c8d6e397faea9b355f848f103707473fe965c4762f9dcfdcc72590951b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0d9fc4a04bd9f8d0c17fbecd390a91c6cf39bd082c85031673ca8d95f63e497399da02d185170a859619c73aa1892197dfe3c3e983e48a5976021105ca5de9ccb30b3fefc08abd6b35ca069868ecaa44053008181a58d84ac1a2f9da586397e04d8537438c074f0fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d644622ad1d2a1ac6f1d42da72f8535f29852717653fc776a19c40107f7bad628a4061d14b5f6a98cc410f0582c28f9913514b2a8277d80ceccb9ec1fff040be110c4256d08b63385206b9b3577e66c69aaf235afcc8604ab60e558d5fd415e48e093a312b0a6deeb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfef643918fa6afa871dab1137cf91724252f9251106ca0d89168e926133878ecc13e18af0db0ab8a4cd22749accac62290f9aaf5ba58c98ea09c0e80094ff75f4ff8077f212c1d5aa6f7a991c5ebc8656ab9dbcd7812a81ba1bae094216d873a2f9888ea676dbb6d06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h955431cb62ae0fc9dd482b91da9fd56a59e55741ddb02b55749b177cfb733b2616b1775ab46cfb306a1bcbf4285dce2d4cd23d087f0f9525377692726b589feacae8718b1ac71faec6232320069b94311c9f45555ee5114117d245b4e63ae16124202a9a025948181f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1685e7b408c41d1870b551cffb12b4212b3044bc4b87b3f66f2669ed4486a0381096afe9a8a40780303a4f9581497986bc67b5455a939b41d155d28d3db59e8d0bf9a22b54df338f76e1c4b4cf015a605405adafe24c7b0c76ae0eb736c4ce7c5aa0ffa16e5e179d9b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127b47250ddd9a4bc25dfb709b4d351fdcc08012f3367cac8471df83bc49045cdcb8605521c8207890605d1550790660bc07f73340ef92d74edbb4a0d0099094511a2a53e29781f2f7ad76296d3e81c718f788721db398ec6ea353551b07cab0ccaa6c0464174501c8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1861227f9de75bb3b4d0000d264ba533d341dcd7ae3eb9816165eb0fef0cfc2bdae7eed6369ecda7b9e04a1d59d4669da5474cd3fd57de20f38113c683d9c2ab45d4ae6c7c51e22265256c33955e4744dcfe5f038fa9fd223090d11472bafbfa6ef96e9dee1794e228d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a09ecea66aa41c1f02a725b7fbeff1014241e111211e14a319e2fe99cbae43cf9616ae78c47119e2ff85ab4cf98d8dfd6f1fda8909ceb1af18f684ddcecf8c3d8812dccff6b0b2c00e43d05d5d418d5f37ce108fd2531712279f3be4bf59502a701a0ef4daca49b9b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17eb4db8a1650b422a8a3f85cc15396f6f9cdf279b33cd9730562672dde04232b380df28c2128cd312c0e3ef6da5efec87d979e9cf4263ae389b1750f0fc9579f74094f9860600c6553f5b085077d8c727439080bf7b41e072ee2e886703fa14bbbb49b3ef41648de88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfec48fbe4d91f390f9e0ba62bbcd9517313a82d61335809a0b9672b826a135227fec400331c99350b2409f4b1f9e0ae980f0168b817e07387e37dfa0635cb78ff0f90df2ea38c113f92534edec2a5f1d8d552d7f780a632efdecc09c4d4778994e1d3bf3878933d3d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9cc4efab6d5ccd30de42f5214fa2f26a74917a931d09d5c709fd632f67c5e31baa39ffb565d98a33b6cf55a7d85992aefd732d8e567a5f7a2da7259b4c0473f9b1b1e9ce9e7b3f32c99437e7330deff476587d1a043f70283ac01ad2ac5b601b9b2053a872eae8b80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3da52249c87a71935469641892eda6a93fad191e552f6799527d180f24c3d0de464b3df2c5fadfe902f844b1999eb5c139f8e4a9b1956e267ee80481d519b5c69356312cd39e1a266314a910e491babcb1d8ffe0e078182e9e326041f62cce32919537db52386e50ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ab797cc11a0a6a9826e7e4b554bbf1fad1b6065f26f06b662d7c9921b07420e5c8c43db4279a008f81fdaa307133ba069ecdd048eca62d3f9390c63afc4134928d11608f5d7426cd1dfde7d62cece5dd8d5945d4187c3b37a347846f2a3090442d6b61741c05d01be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1278ed5b74eb652be33aa5c004b9b1188a68c9f400a079441996c192a138bbf196bb1c41de00049bec1e98397cba9f433a1ec4aebc48465dc973162770540380c6ac25b1014c07d3a33af0918aabe477ab5d2d232fe8d3a29bcb2866819e6d5d231918cc96a881cab84;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e5904d24e5eab7f88fa77f9a159e2bf4e58f3f881d6548100ebf8fc2eb105a60c38e293fc1861124b03b4ee2ceaad131eba26065abad54c1f388528fc8ce7ee202098ad78829539516fa02c52c72e4867d22aa3ad1eaeb9d20d0ae9113feba666bd5ea0dc6246c89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he21b48237658e2c4e73f01c47227ef72573ef878c91f2684905a83c1d7733a41a670926bac2baab098ccb92bdd1b0b42eb8f9c78b5b3bfc24692de02726ba777860e5743e41b389f2b8956f7979193a9e5c810aaa0fbc19e28cf358474cd2ed6383f00d9b9990334bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144a11a6f561b21dcd30a369d0fca98ab311b16ac653108eb97de1f7d5fc1441035e832e22a6cfb5fdfd4fbf922d8c385b6ed571469f452ab1862f8dd1f1f56dff6ed0e7eb516b1d6224a1d3d310db76d4652725d86880909d65db1cb1f8e1940c5448ec7269564b2fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bbf2c2a01a39d88fbd874455d91ccaf560108a566c0a7f7f758829394cf735660975496a75dd8f0a9376cee942ae0efb4d8959ea1acc833433c525fad3c194dbac7a43a64cad63fea758ae9dfea82276b4bbe816a25f80dcc9314c63072566089d0cadba4f0cdb12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b08e5f79abf5d6443d3d1f03a2842aa96413ac6a578b872e2e5e24bf61035005abc927370dd05f9f28f26176986c17f5ed79f442255617c6c66c7396a7297aaad9962ccb14958e9dc7716cda0c74885baac802d1a9fd22fa649015ef38696cd153f58893d999a75b08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2529b860f923b9fd3a1f259d7957261496b3ea2f97f0fc7391fae29d4b53722622c3f038f9ac2d2ec2afd7dab3e3e644377a15c81b1a235b2777da2281c26fd1453a07ba58d08ecac8c310372448810aea594aac05432bb4cb9bebd998a15a29fbfead7e7fd40a896;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fac85dd3467f099385e72ffe28ecbb5fc6305fa3b376b291b422dd4e706a0b853c6538c5e309e94b6737e1abdea5a250f441c1c38060a05eebd79afc471ef73a6404f0df910df3e0c465614ac029c2541d858bda5291dd845f71448eee5c89d616e102a055bc728532;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4539b13ab40fce9e15016865c441fb899e6b1c2b940981cf30350f83e711f651ecdf1e5d676eab87abcf0d9ee1230743db92f18b22e394b7a274f846e6d3bc2997e41991a685cd03311321ea4708464cf761b4f13feadff55242bc2dfa09b79badd584ce01cec394e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1419673317cfe87063d003cfb322fa7bb10c538dc6dbd2aa93abbddd4c0fd063ad1bb32e1a8cd8a363a6b8d0270d57d093bc675de3b8820f0ab56b6443edfacc4be88da27070343eacdead68849ec95d9d1ebdc2197e017aba23e6b30c85e4ad53d5716e010f4a93712;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8cc9533fba3f78f4eee0da47e270d6eb9a62be7dfebc2d6c056fd9bd239add29c8f9975b988d693d4519e53489af55340d2404cb43afb39d8a550b2cb1fd74f8c786b2f411d7195cc298497d9dd4097ee4a6d64859b7f35c6f27a226bf93c10c3e5a7782a0e86dbca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f78419af2893b6f0390d1c3856110c7eee4c978167fb46ef0ed73fe5a8c5186b1764d77860a55c44225d1e4afc72a28743a4f62682f35cfdb9ad85aa95694575c79fc064feb383f4589689b8c55f5ce54957bd0f4dc4662d9f8ea5745c0f1a99938e894cf4969dae5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fa1906c7e99ac39d3c99872ee50e40a5f535cebc86401939f009ec94e47d0f0dd060a36290a10cfd4d1c28ae1436888eafdd8943978dafff658aa4895f3468b8638ddeaceaf4ff9e51b33b6b4931e7cb24efcad910a48c7631adca3f83551c26a45e812f6c08bfc9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48f343aa5f566ed3d851aab8603e5a565d4f5e1edebde31ce55cad39dc508a65fe2fc63ea8c3fc019229374b86f250615d43faf66776a1e9d2ba43820bda40d89153dd34dbacaa482609c7974d6817e85050f1547e97ba9c20512156842e54b3648dbaf3caec8d432c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d947d9142c6195bd4287661e9c8a3a3591df7ce1bb8782604d3b20e4da35741ee13238eab4cdb42a024c7e20b5b0db5c464866057e7584ad613a3d3f2c907deb045efde04d78c3542eb1ad6c3711491a8c73ce15c34b0202cb5a1b16010445c1d21cf848a1f55635a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ebe90bff12efa7bf5bc773eddcc7c5b7427fb4d0d04a8bd78143249584ce901e7ac44d66a3a6915f9507eb76108909e490e4efde1ae9823d5569e2fcccfa0d599acc30c775cc634535a506c9600264052fa314c260e2eb91e402515dc85865de56d9047f352447458;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15fec8431ba148af556568bb202bcbccba31c06e65beeee096ef2c232d5d56dbb665d09031d33bd434357173da884d705823d6cde2603e92eda0707db8b42353f6d3759d48d3d0b10c94d2dad21e37b3ed4e2022bccaf419e1f6f7e09cbda5db4aa8ea983f07b89c563;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153747b9dc4223d6a53baa21451ba8f88023d516fae850fecdad2282fdbeaee6caa2dd4e0974937c8f4f79f7315719c489c7b9dadcc742f9e33615b70fca56fefeb66ffcceb3eaa00ed4a0a2f53b6cca4b3a6481fa408dcc5cc4c39fffd75ddc9afb2c302320a28663d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79de753d54516e79d456fd6fca018d5c71f9aa764bf9e3169a353fa697a0f62cee703d19452075c3be47b52d53aec7ec22989ee76f3d313ee8c8b80efba0b65f94cce8c8a55b5b9d9fcca4d2a1f23ed5164037de72f9cd14624a9d13dd67ce079f64faefbeb605a6a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1448b0cf5ba3e7d9c590582561ef5d3cfa54d75cc1e66a2c3d4eba3eb4a947716b4cac23b992c91f70bc9f46ab022d28274808e19a97fbfb08fc02d1a2d63a72923426ce97969c0072d985f9df0a36300657e74d54b1246a6c281aab3b97df2366520cd767c26694325;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31945b94a8ea86960a92fc71654d89f33ec8af2ffedc6cb7b142ac2edbf883b05c812a180beb7f86142ac83563149dd6b8dfa16a609f0083822440a4ccb22614dcb8a9a91207721060059fc40f34e1ade5252456f89ad2cd0e7ca5a9fdf658f1cc6d405ec628ca3c2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81e1bcebcf536f247c8189542aa14a5b60e75b5251db21caec9060da3622e739e4911ed19730b43d609101e0174285685c207585506fcaee44bcabae4ca10fb98699e9e17f7393b25417111b60ebdc6bb8bdd2f68321928d1c0409c390a024704d99f16d451eb80d19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184a8c20cb73186abe18543d229fe322f44dfc689f8d631c2795e3206ef22bbbb79f53dca37444eb57fb7b9144754c540d7e544d4a256600d11aecebf9302ec81cd778f8e81097bd32ac3000edc36aa003afc3530e2fbc9881e33203790a222f2010077e1c628fe0484;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea4de207947b46c2144534039e23622589d80fbbe425cfe075fbc5998b67a875d0318adbf0446cb274944a3213d4a630a2c809d128bca5c996a725be07c32245650a895df798b58dffc9f7167ebad148b33ff19a1332e9489d55044975f3cf6a58bd637619a92cab04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13214fe51d3c6e7d172effcf0c91969064ff950c5878d60edbd9923c18cf59ad9ea56c8c38d70e6b405e08b211142d885d384824617bd7fa863c4954339a179cecb2c1808d180d3407328b7e8baf7f39cd000d0970e79d37cf69a3e981cb567c2452433f8cae56f0089;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d7612e75fdfe0d78a59ec0b38e615fd8c197eab4273c288c13621022dc2094af4846501ce56cc5bb57bbda700a9fb2ca9729525591c32a0a053c9eae3e32b1b701310110258ffec75481fe6567c2f88f8a8dc4d2deb5042d5ec71eba8c8f464ee8fb4d4958ef67b2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12aee0086e5b7f5c15c6c88a158edd203c609cfb8a6f5ae96381b2b74b8c27b0684f2a3dad044e763aad591c74c0e826537d5528ce8193b64fdcbabb5856f9896297a3cb1e8acb0e256e29a298859b52b20a859982ec663f1c93118b400367dc1610b0c89f67c7c8a48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ab807685239a8cd5ca71086da506bbded9cf5635b1e4feb63ee73249c20a0db6815e2f8ed4a0ebf591939296a09abc630ffb8661c500ee3ff00e6d4b89ea4cdf4cf9ab704aa71d0c421431091a887dada813e50851010d5268f0107d24ba3457b9345fea0264338f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127cf4129d5b133220709f340f12bbb51c96b6c4e685708cab2c1af471c3f7a71a9e972c443938f43d8501b1401e377b9d92b69b45f9805f6e532ea3559836e3848de8028c4fb1677a43f277cff20d6693313e57325050d2f0f1758259c063f6de59a80f68ba55b38f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160a5a5a8fa258b3f811da4931d3348ef37c4e6c9a7c574ad77d74c3c9f9a922ced8383b689088f3b7196e8f74aaf939d20f0f2af2905442fd2cea357f098b29650c5986dc673b281d83108758374d405a546ed138cebe3d02df1cba4bdc5bf9d3030ead7b182222ccf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcfd736f59bec8d23d410208f64c1093be64a7855e78d18e3715685a7c30ad74d330f5e11241af0e3c68b2470ef8200ba88388b3f5d5ad490ef7d4c1e8ed733eb69b927ff2895501c54b8c8e61efd057611170d541909abfd5a9538d97461172ca2048704ff77a09653;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd5f90bd3ac2b7a2ce20eac0861770bb2c19db134c8b10c6e4f4a7d5f19166ff2ebc938ec98e9ff4b5a9348101c8d96ce2719fd00602559dd2b3de32d4b01ca91385d046bcf30a74c5d56fcaec947d1154258ad756508090c608fdebbf7e5901eb75f03c46d6fe08a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100906dfb72d8986d8dfc6ae11d588c471518a1c8ca90f1342f7e117a858f5a9e45569c3f09bbfef52c4cf7f3b55cb875c58897b8e8430ce9821e2b99b6f6bc09fec270cc7b1e42d4c1a92b3385df5b52354d2d6c0e291d941aaebe73e4119f1ce1f91b4f682007f278;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d280b56e47edacca1fe883851020006602ba4d7096790844f6350c6bb6f29d1874630ff06a0d4b116a50fffae625818af3a961addd84912fd57f53538d4558751a83e855213229fa3b7bfc13ff080b86f15d3247b181cba5b52bdcef17386efd0ae705fc41f47fef7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h706837de96d6ee2eae48efb5090c8e955a79dc436c72b6c921053fb44f1e239b021fc7032fc9e6a264b462efea4793f262bb01bf7482dc6caf9bc8e462f3e9cf152a32a6a05aab8b12b1a1c50e86ae1300f3f94fe295a769734aabba8d76339e7862af41e857cd9794;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h767ea2d1c362aa4215a0684b3146831980812f0db02e8acfa75b990b3038262e0e6646d16b787afbb9849e5b936d1f2056f369b9bf97e4ee66edb76c41f21ca6b3197984dc6da92651184ea9721897ac82405d851ffc64f5d83dc396e62a96b8524476ba872a4b5c7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4a550bb361858efcafaca9bd59c18cda5484c408125afd9c69642aed39fa7da9e5f114e7fb2f1863b84b1b0c010b4811278b35a5fa29bf431b488a7d50ea2c0cbfd96c3ce7c857c96e0a5c167fd35da9c3c47a7476c8037487aa071f4b6e5ed44f078f0f62b5cdf25;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf51212cf1927a03d168b2247f9826b9c38e1669c1d65e1335bf4aae64dd0758465133dd63d68ac5ac5d5bcf2675c26e4f9c86c0de1d0914e24f9a4e825b128aa87b6e435f6ec24d4ed03851358f6a07c760d3532d2f9e1c833a3914f99bf2e3732fe85e00b142ea614;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4464e57f6b3c4509b7211221a9bf6ab9579bfb8faaefb68756d24a1f3f291165b48e9d5bee815b26019a31746a3e7884be06e9e59fb1668dbc6654b5a660f31e86860e4953a1eea0f7b0eb98d2819a3c0fbd934a6ee11b5d691b859176cc8c64c03bcc54de6b539765;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19480393a541b11aebe4782e1fafa6506855a3d2f173a7957637bed2e1d750706a8bc9125e9a62e242965537d5468485ee4f11e66060657868b92ae683a9bff9339212c6dbabfc61cb48574c158ece9207474e3883353823cb76be0c5ebc263d3074f803070e53fde2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10cc7318f12911cbdf4e2aab9de5388112286379f03c6a614e3409d0f791f92cffd3109ea7aa0674535712198dcbca12ccc6c060b23c388ccf4eb7d23f5bd6ded93bd8358e2e2699f24d043fbe0e4e5d133b109dc1ec9a21582b7361d1e34ec1adf65e0d7cf01324c05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdf8d3aa67aba2e35464990e7ac9b0ea444c41564879c004f8f8f53ba7fef195c343959e7a583dc16d1542e44c7117e4d3b805699896b5aaabaef8eb319710d719c47a4898fdc6a16ab6cfffd10aed10a32185edac384d430709815053048cebd74249787a9cca1277;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h373ed39180734c999a258e87d68a9bcd5feac4dbf63be63774081d9f7c116ff70adc1360a9e9c95bc059b06b68406845c2ff56a68244dde3c0d67a003209a9ce0bf86161bb3423a80b1ba553ff54c0a533021f71039d643195e4609d2c73994aab6f3a3f6e6cf38f53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e353b371ceaa0320cffddbcc76aa965eb65ca6698c8c4d656af57ea11f54c82d7abc4837cff030df01b42e60de5559b48a2cc78878ea285a5b8fd018a6f26bf32560b0956ae51829e31a4b0db409f182996bd095b68d87f410b2df31a27fb4c62b239f677b4ee42ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17aac524ee5988ea45da1d461df1ceb220d0087e9eb9b18fc2f78983dd0ffb72e0075c993ebf9a47c11be8a9106f09edb6ed26a4aad003d65988a8aaf7a9ad9a8259205e225cca3bb0e4ad4ba06b0125e006a9159f9ffbd73160908c17d69052aab2c8ca70cdbcec9f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf352e56f303e1a89e939ea549fb19a0deb231628c1576fbcdb74e866e9c647c893543cda99f5e6dfbc98051e3bc9154b30657b650c2e3a1e0e7216ea061203b9b4079908f1cc49bf2648e6ad506cc12696fc8e204096c6e1c0d9cf4da66e53f13e5eb4decf115a8b4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64243048cb71aae8cfeea8ba458f96f1f15fe86be03f101a66f9d88280701de91170c83536dd3c7f5d4787e7a2d6e1cfcf1dbc59d7e613e7aef12f7e2c1c2119399604d25c129bc51adf6c647abc1473a2de0cdb50e982011761a8adf553692ae9f9bff7f26d20df1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff67e613ccb2ad728ed47dce6218ed3538f7539d86cb03a1bacee9b0147f4e18557ba3ad62e3f4cefa9861ae800477544ce6aa19d10d901a11ecc2d9b8d8d13da8dfb1e1b13e83e92567716f7f790dc478c77cfd998d809340a3b9e7d418066d406c6a0313faeb43db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6995514601ac5c28918323755d45af5007c54263308846cab4871f895aec708b369892f22d75a8f6b95c617109bd42b246023f6af7b0228a7c12cd1f726586fc05ec7427d431866fd264439c75671b3831c34131edc25c40a1d2e32fbef541e208221b3808fa7cddd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67e8c1b35e1b05fe2dbde884bea8b3e48fe3627c0b2b3f95609938ba10259f615601416ce1400dc6e1f6d21373e328f7d95867de7731171a843968c2524d0b7fc9c538d1e06e55a8ce1c96ba5ef05986afebf9eecdd1ea4d9573b870fde575ac8e5f75aa9f2e148190;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2fc7564fb218b5b2425a20dab5fda6a8061452696dd892927e0f7d136af14078e41903b424ec9ccba8a2fcd3528d8f3e7ae739c2a035fc62f63111481ef86343a2d2de4c85dd6b3fa488572a27d642991fbf6336928e0bf58dcc0718022c8f56379007b9fa8a59d96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b4e54711dbd1feeb05a414910a3a5ed5adda775ce63aa24cfc4df7cef0714e48f47f208e1701afd4526dfe992a0054165c6a2a00b883a444e6e89df9916981ba400ff2a369e215459cec022fb31485b19519e9dabb009c339531bd8f697bdcdbdc52b585ac459f6e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f819788cd322c5941759ba5784c8f4aaddd39e44c459ea503b9245f2d6c30d5a9422fcd0ebda72c2d7910a166b960c543d68da18b56f9ca8e93c109d691c88890deaf89a149f4201f0fa4750c327b0ddb442ec4f47ad6888f4501988781f5292e00f3e7c45331ae2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b4e75253ef2ae13a9c566bf76d5fa2f24c2dce9d80243bcefd2a17922bffcb6472cd6910683f8ab5d14435c1a80008ec4562c91849df9f319a86fe651bcb1ce608dd7f6b10efa31888df2a9d0a708227570985da46f54930f03b83847e8464838fbc4cd1f826721a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd75993a1924060fea34f4e820a354dc9d3188e5f4b8bdfc1a51cca73adfe3e44aa6e7ffb6cfbae7b1d2de665bc96e27a1d8727f03379d041649ec2dce513ae6d85d145f658bf727176f6b4b8025860fab3774c7ad96cdba18fd77eef6f680324f093ebbfb310fa368;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b2abcecaeb764c1b03e972c4fcdd8c5ceeae5b7c223afef226ae0f1d2daa6cd278128f5c7f3413ddf814e038c508c8d03e64984cebf29bf0712460fe1c9de777c87903931cce89be14f5448939d636becf1ad9e1face098e31a1f46e554d803e8c574e7ee2e5c2a76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85dad2c083dbe6d9afd839512d98d1bf89fbe89285afec8c1a159994218040ed02d81ccb87ca8ee5838dca206b1abffb6d9731be4858d5a155091322ab2368e147564cc43e6607b609294725e77846d01928cdb9045b7a679e8137f4bfeb9bf768cf9a4a08beeffe33;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d3311d073d81f74c2409d28fc0db355a2cd15fe3d9be837c5af1ce725d8a1a5e3875f4378f0061aad2440a11cc03cf6fe847e5577a34c17dca0be72767e0ac07b1ed09fd9a8c49e5c1e9ac2bb1e8bd7534e60e438feb6999c67f30a1935db5e3dac419677cdc3c6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5278782a241671051fa35fe644def7831e9e313179b223ee9ebff31c06de903b54d70e7de5b63ec3ecc44d3df24a060691c5756720ca1fbe81f72ec88cc3135b405ca41567972bbe046fc6eeb56bb106804cebf32203f2ed95fc6ab7e46e01c13dc07427085f15a38f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fe092d53133e3d855dc3544db13c9a242c9abc939c02a1f96aefb672cfe078072673a014942fa96bfc6f239ab1e2d7e7563b6dd4695aa4da3c7c2d22de09392bd471bcbb7ef373ec9e8fa295a5aa6005c3bb3714663ce6b5996b170bd7c77461b06be652b3b7671f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b1d17309da28c53f738785e1cd16e586c8c1f7b790ead07d9b418dc3ca93c9ddfe3de451280e0b717b53962066adbd514119d44a2b3e61c9eb2f3329b4513badfcb96ead0e9c4cfa21c305e181b2130599d6e144f6f7632e4a90bc93a6478a8e7bf62a5c1be7b5ff8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc1e9187b33037dd5bda839ce087299da20af2f10580eb87e44b8fefba8f0b8d4493df76eb6325af0f2718b94103737262cf1968a2487a67f5c5433e1f2f2eb53c1780964684e0d509a53b7bb3b442b9237e19e91f72c0a815b213eb0a898872705b72e3dc1c948a04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a2b39a2bbe21f5a428b0f8443477ea40d614d59994a1aa168de99f42293d45180c8f7c93043727d039164acad6ce0be30407a8cd4bb5a62bfb28df60c4530b00afbebbe239e840a159352709dc730976473d8efd9db2e94e272d00ed3becec78488265fde09287266;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1762c3567d7d7eab3eedd2e277996fce6c6de9b979b79bacc3ddbc3f7c1643d6f4f7395904f73b1be7be4e477d946b83e26de90bd9438590dbe1167d53ab263a81a5e16bf3ada2c85b892b2fc2af32c16a9b0f9e8a71a02d57048f61873522f2410d272184937d0eec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc42f2af0509b338907deb15fd3ad96a330a78446228d6ba4c8765519568adb23928f8da8c7a7a5c2faafecbae760d6def1cb4d35ce050e3de4a20d82edf169f2671ba994d3f8e10b2f70bc2a7c5637f033f26ba44e4f201d77689aae6686d42dec1fccae2effc71148;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79fc9d21322cfae95b4c54034bf2a11d2760240710e1adf318cc9e8e34137a3875298f50d46963a1776bb9f2f8e2a504954b7f35fb007ba813d4c51e79a423103c74c4f2fbbbf1dc4ae86b9beb2da32c983e23869a57d4b5a85468bd68d9b1e2fbc792fa97c8f92908;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f72c90ca135665362a58bb5d0841cb8a93c19ac5cb626b35dbfafca7767f089d93b02d3d12349aceec5de114f1f19341bf64615f544be32f666f818b63f58202918b2c951051e950a0fe4119fe8afd934aee95b9d5f658222a4dceaa56a2de0430025d5798c30dfa4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149e7ee51ccbf97da986550c42cbb0d16deca708bce6472a89fa91962f09149a3872a8447c0629fd6c52159bce2e496dd8b573f5e49efeb143279e6f3557eef1e243a5416649750ee44482cfc3f6860a53c66eee662e099914aaaf6e5cc1e0583dd49331a7814fb1ecf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15aa828b39e68409788c11dc590fe91f312e2d73286e1db88565f206d0c45d5e1a28943d7113b8faef29fb0cbc5da09f0996fddfb25dc683b2f8c5cda39f2b6d8a19573581e83a2d5814788bb66dc310816487c525db8dd4f3b7cec51d9543b1a71160c889e9c27818b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c65ed6bd8b2e45d67559613f630470073806a570532e75f24d16b99c56fe79e2b4844f09ed574e699e1cc6f41a4ac5d18dc38910f87e0e86f68b57022ac9b263dfe9d2b03305bb924905cd90cc566e329d041900a68e21b546eb6c76a3d19151e97656f52e227bd1e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4de4d423c12ca221d60c4df47c37df5d3deeee0c155b2f6be1851631b767918c5280a3793afb849b0c0ba0fd6e6b65785d468af0506dca01aa3f199971435a87dd5df77f2414722c87e02e2f7affd060e86e58f2731c89ab47ffe1b4bc5f2288f7bb16961fffa68f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fc83d3dee49ae6d53f22d7066d1bf96c3a85a28dcda22e5b22093b7ef031df3e6327a7ee71a12a77a9a6638cce24922261b80a590460a86b728483ad9b26e0c0b3a9c5b287ed198223c6bfd7ae0d50b31641cc63d96e2f9ac29473cc3da3cfdacbef2cfb818f02467;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b98a55c823fd50f54cfaf7afc3f58f0eb622c56504d9020cb85354c185ded3fa10df11ed2ccf7342649c1a22a88d23bac04d651eb22490309eb75bc2f8c96e655c700a23034cff2a0048983acf77ae39acc9d9929ce52020db7a81be4b0c0f1be280fc50c5d7a017dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4cbbc125adba5112beb3b358100b3c458f1b788a3dfa487d600706be18e30fdc2fc62862ee09e378fe6963915721742372578b2f9be7413e48468e8c5e1dead1e02e567c66b04d526d043e082e35d2fdc6ca2bdad2e5b8ee14a07068f6c3f217d0856328f5ceaa647;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65044d92f38c8777ace79bfcbdabe3052a734585bc80c28834021b55ad4f0bcce2f5ec3267f8ddcab1f63f1a6bb7dc08b073c776985d6124914c960573bf757709c2cd6a2d346a15b44346057d751a60f68417d05aca01d0f5f0539cb585e3d412f0c01ba7377b2d22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154daa9d6d9feb8d4305f9d8040cbbc02d030037084c1d71a5568e232a19bede4e6893a4fd9b673c32e898d9dcad2c93c07651959b654c071226ee4c60d3a8095309047f8916e0497bffdabb1bed82231b50d266f83e4e61af158649803b5dff1cc39c829306b10423f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaa9a395e9cd0610c32a5ee348df102dd43ebc0d239eed5f40bdb85fde1bde4d3109948a11fc1e58207358aee911316f9aac8d021c020d715a5d46340194ace5f40a141700cbb9e3cbe0a064920e070d30c96b0063f53d62e77ee01e11dc98f511a64662ceedb0aa10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c4064940beb609aa750aaba80ae4302ca7d48814dffb41d00d479be8831ea376b7bf6b6e6acb465552c65bf917d352c44186d832981b05940b804c2743aff5030b87a226c610a8e89b6ca50a8d89da5e4d3bc1541b9390b720166552ff7a49cddae319648ddd0afb6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b713946dee5a7e2f00c87a356566817cb6e517013970220a285e0f70dc08868fd8acb178d9e0106a35ca7dcfb4ce4ca27ae9440094eccc1f2591e133d3762d37dfb198ad62dd0a17c91efa42af0fde1708effc815f51c17a5e869246b21489651af098c259dc53194;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdaac157cdced18e34ae4ba60e64010bf3501b7c0df2a4f1b013a0b39030420171c76e1bfdf8510212de12a24160dbccda1d83cc8b8f6113f5dae257bb561aa5f5b7e8d3a2a0c95a9bd02a806de74dd6e7c13297d0771c3fb34d7c4abd015f791346b156a0c1865c034;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f16eac147528af64699272b00099c246ef817f2b8033c2da8e9b861ab4e446e2a5bfd461a4f943358139f9fa6b954d1ef31c5fb5183ac18b2c0db4f6bf56e49984ce26da798689853538186e8c100822b38846ee5e60060b3e505e45ea96b81985e1dc397fdefb80c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7d34c2aceb6cb77dbda195e9ee1a789bdc9bddc1ce134922a9e4dcdee6679beab3e1e8d112c7c536655b9a4dfd6de513b8875dbdf6c1cc2da4e5d2afff417ed93f197d3b2636fbc13a6fdfdf9fdc60acf041c39b79b14adb89f452ffc225df3edf00834385b1d582a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h334ce9e750cea3843fcfacff9efa69137be6a9a9c5cadf86425ef1e598d7d8ab19055401c1d054ee600312c2c5d84561cc95fbdf8edd63f9a3befa2c3c19dab361488e928a4b4a5acad0e99ecd3de690f9af6b113cf7a97bb8c86c6d2bd3e78adf9a76d8ae1a381069;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b0306a47016e5d61129cc394ff4c04811bdbe32327ab47fbd1024abed44ebef789feebb9399ad2ab59c27cdf52aeb6708fe2c762e3f964b64e55a947c6e032fe06fcef9dbe4e059b3b0219802b298a2ec9d2451b1d69aaed3ea1515c7b878259899f0e15bbbf0b851;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92bb20936efe3aea0ddb52a4e79ee6f45bc7af85182001b8fb7eafb05c0af3316908559b05011d9fae808b76b5c2488866534f9b7ec8a04e3b23de0dfb5d49710e639a604c5ef49a2c46fba51287810e9d44a78c63b21dea75a480881b02b8e95e9ed26e93128741c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc092f93c1cd503b0241a488c007ce375fbb9023616f4ebd3c472d533064ce6b67028d2b6dbdfeb1c7047772bd939854b1768af91d2c24b43cee51549baa8b93d64df384c0d980d32f43dd84a431db38a4ea97a7931749c65bb6635cfe0bd8316775267e5e4249f201;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f84a30291f1c620c2c113de6c6ca398c597be548456f7714531dfba5abb85f1030d9a070c64048d87ef16c95ef892bfd9abaca415442a2aeeb51985574af96c5f7f5309b207bd7930cd4edb35b297cb8aa9f71a75c3802f682125f2e55d91eddbbc14ba005e40370b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1889653d02bf76c2c949e79f3aaf594542fb18b41eca64d888f78395bdb39170e6defa22a44f45c4dde181fcedfc56dcb12cf9a0baa7c7e985676c97996e727e9aa916859b2785036fe449ef3cf2ca1d1e3592464bd8ac79d279b66c2fd51f40146b5402e62757abe90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha75b72dfc5045d59894a42c15ef642e9d0a9ba17f9909f0d7741738f1bdd95ded478132fa3d0aa2d7a24258058a9ed1bf5a8eaeacbec89e4a24154e5b88c6c18d11110452ff4ad0529bbc4bbb89b0bc34da76fb44f62ebeeabc6de2b6a051614976413065722ef91b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca9dba96d1e6f671c5030072ccf93eb56041c27a27b44917a83f41911d6b10205b9c223b07679ea556b12facf96a4f89edae0b376ec2d9180918226b3648fa6aa91573cd96467fe8f2f83b21bde35b523b681cf8d38848061d9eb60fd40dab6f581388282e76e168d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec71e1d46096192486e5da061fee0d59b178b491f5bca8bec8e68edba28bb30211decf5a279a7cdf54e961d27d8feca67854744d9b36665fb449a4a38c9295f689ed7623b90f06571c8cc45013e20f976c827db7bbd046662cc5c3a7ca6955b03aa2b7292bf70a299e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ced33ed1326f5349fbccf78399f17c859234a4bdd28cd8079a259374919da7b40b8ff478042a7f607cd85e3500bf90f22a9b16d555e2dcc93b2f94c023b28518324ed048770a17a5bc1f5940343f0ded64871200efdf63b3335862336449c0b64a3ccbd990c8f07ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee14146ff1b4fc237e6a33e1b29b29c15415b21bfdb4bf3af3313a1106a35e38ad70bd6da949e7a40a030fe2e3f4b9dc4e789b6ab5920304989620f495473d1f703d60325c3192e7a2b0a089a69614fb6631ab027c975d52580173c319aa6a3801bda7e91cb07aa3d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152cf2abd1bc6d0072f2c0e1c3d4aaedb83fcd7f02f9fed4d57f9b3c55625fc46b08cc532a8dd0a218f2db6381eb488672128e6a8dc35504cb96a10caa720805b1c47d37bef103894e88b474256588da157514a39f8dcff023b51f858da5ec570fb924f99817e8e7e99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14899902230c6143bd3832e0908cfe2f695e894c6fbcef9c4fb9b5b243f9d6de796ad9b4cf79671bda835f4e79b1fb0b356631aacbc153686fb72c2a4b1a33a2ec94ec2788a4f47d9457121bc713bccb526aa1552baf199b7d615d891e84976bf9d0bf344a52f137e27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7ac5779e69cae929286a0bb45bb407420ec347d3a827a0caec1e3f6cd1858a47ae11e2859c48a240daf9bd53fff693975312fe8936af5752ea52c16032dab7375c0801338e4cfa0e1b48897626c174c6f6a527ba07fadd6f876f6b410e38b863e5adf9ee95b21c270;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd348a0f5dccf2709d239543e3a8a773c35d74a99b19aca71a38b450e7134acb246d291b1d350172a8aa21d1040834939b393da8bd347ae1760e5d8be5dc8ff6572a869ebceae59a1183008dac9902b51314cd2fd8e5e8a667cef3aff6a4b1199631ea7a3bed24ba69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha34d8f76a21738c9df8a86c457eebb820dd6d9d618d35b17b054e7f653fc3b769dad8381880029fa0d72c906b10cde96eb4a59885f7fe77163304a7a413492ab8bf3f0078fcd9cffedbff0590c3dd5bf7bf598a216f97ea35531654160ab04b5ca6d2353ad8b160580;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133a11b1d56329d4bfa365b1c348da2afa1617875b899236d5d2b9f7101bec5c82d00eeeb6621aad8e41778c40caa723b8ab748c86e011596157fcaf217c276c3d0d0513e39e930a1690c86caa218299fa61dd68b0385f9dec5a10bd740b145d14910b0494ddb462944;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he151dbe713d1d1ec53cf90f7f0e7a95dc7546a53d78cb059ca55f54485542608a27a724869c9aa72b505d85f79975b4670c96ac2d2df89ae653483ba073d6db24583e634d629e4e5ee6801c025b7da47db13b99254ba38e02fe743407c0c320e0aca7e198aef84906e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h678cfe88af2e5d0390cd831dbd7f4ebc258bd15e7456ca5ddaae1c1e126af563d3f2a49db6e2cc8164e635be1257da240ae95d380248b5052c00c019e2d695dd841e0495d2b337003dfbd9001f9f42a38d630d83dd0ee8a57f953ae5f88ba6b3fce2cfc34020441887;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc10f9540e17f692712d31adf08f02a3eb2f007891d292847fef8d7b5e374b7829c9221f0a66de9ffe3dd477a7775b13d098ddc717b5dc9ead32187e091733f155d6981d258bb70d79c17508be78664a38077612ffe1c9a67d65bd2e0e22d85ac790f10731e86a77df4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4d4c1760b53e11fdd62e4f68a8c035123c5c4c1f0f7e25702743f733b69dc5065c084ec65b506a3e554a2d847aed899cf7d03f3fa70309079b3294de59a043ad89cc6457c89c57fd17f3a18dcd8f5d89c4171a52e26a41801be25a0f3e608cfe900d7cb330de5de16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d7d66081a020b2e9152431ab0942a7f327a70e57f2625d9272344571ccd4713baa379ffb3c232905a19e9294558cd15003e519558b86ffc38bb3c46ec0191a3646432b6bcf3ad5e5937bf6f1b06cd189ab75bbe4557baf4d97e715a9914678cee62ab200518f89637;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c8616e5864cc5bdf293b52ce0c24ba2c3e14e037621355e02920b708edf6e886f973ba1a6fc471920dc5b4d373e930d862bfe954d413a05b85f1db37a31fb946ae7f56d14c3cd33f35ce02eeb10ae2b4c589b8baad2050a4576faa80858ce489c3a6e0bfed350469;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112fe105585b2aff57d87667d0ec512988b4da6b18e4f07198fd78ab1bc6a415713671cce3a59219b57ba4ad7ccebe4586434a56f56e39b9066025f9399c2d1f25d2d81ba6e4c1a6ad28adb772dc60b5c6b427ed62a1dbd90efb1d14173602a494d5ccecdc8abf23570;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137213f3ce65e58669bed6c6e48f69b88baa733cab354eefcc5917ff630672649ec74cc8581615a365da2bf5f3bc3a14e45737f9aa6c520fb708e3dfbdb2c0ebfb31dbcd0ebf14b9630945e9f28bc3ad2d91bf171c4f5c18060244ba8c4813b8d83019287dc5cff4cbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce83cb128b87e06f412a19630f2e419a0292a1984de8cf5ab1b3fb2eeecd1d96473dde8a98bc8344b122efd33c20f6230cc9276307335989c3f39916e88e4a598d89f5bbb90903e1452de868fc365f80333c57213100590b78684a7f46786e5c99b7d068a9486307e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17160afdb7b7997823e676c1259859de4bc4a2f75b326722aa8a94f390965bcba805741d76db58fae9ce4ddeb35cd2b6d0b14a5dd7695affe3d8c81819973f2006ff4b2ef3ea09191895dc0ea52b51381ebb7702568ac442f0f9ecd1a52b85c19265f6ceb17a505b312;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dafacd093f97f41ab35da02b9803f3e51e71d4daa1d69919c097a0dcd9c595baee655aba1e44b05817ec66a5d5425a4bdffff4c20d915ec1df66441651c0401af9d7bdd503a581097d9389d00e8585eb94230638c8e1e383d83228e649b783c529a17faccfbdfb8de2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fc067c72e3df7fc6f2e627a17b46f29ae23ec52eb40b4c9a53bb8aaf9882ea3c636eec54ebbf9cfa95abcf24d2fc120a2b83437c48430242034f8eb1e4a142c935f419beb1bfcc42aa40022d8184f68b11c7b9f369981a26d6558cd84f85b6505bf34e6fdfd9e56a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d0160e81bcccb6192a61fca0ba751d4da84f59a822e392b258c48a080de2311da371851c507ada64ed46e271e9cf4f1bc1f004efd39897c90381f64b01d12a6a922e8fe91ae11ac228c0e781e8cd008ffa73495b7b182dea8d0cc93a0790b7a0c02e470ce309c1f61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cf04631e0d2dfdb6c40caa88df2a3283b8c51d67072d3aaef271c6be61f1fe4e3e41e19aebb0cd4da8c0a823ff5ffa0fdcbcee89c69b81d76e53a9501bc3b6893d8d1653b5f2df19fc09803d71a3a58d3e04133146cabf53a3295200e7384a97ad3776b355f19d6d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83cff3e48b21ccd47b4587d4ef987444c30920a54de7e5b1b725033c5ebd32bc4149103381c4dde9bb944cb4722dead9d627455ed96bff4c5a475eac333aaf50360da020dcae2d464adbf997cb9be0260ff768418dd6f21c617d020148c196c1b14b12ea24aa986d44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h756c5fb2b20b97bf2cc4290469ee83a15c4a3817c96f2052f70f227113e31ba0d90db8fa920efd5364c63c18e00d827bfc8a599bf6371bc4d5d05edd53908623b54714bc085f7a06a2d75ae059a09f5ec02f414cf59adb752124536372f4a1e4aa1939e4cea5f16184;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f87b0ccc6f3d5a5a64c9b29672cc020697b3ae88c26ba1984718aad7a82e9d8e837020f24326451a485028a3eba9b7d75325a3596420b4c88c93db80ef1044043e70d4779828d690f7302cc13edba6049bd1725c5345770b1b2d036683c0dc2bc719945a042fb3855;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a648606e6bd6c166d204ed63cbe1b2d498def64671a0b2790832e0dc30153131cfd5ab4a914a2fcb8467fac12e21371434d9d23fa14e1c280dd5b877c5957f21d0361c7f7616df14175342ac035a1c50193af0c577acf701c464a2941bf3c4870ac2e6de4a1af9a8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h223d0fae3a5b709b19ba5d73395f3978acd8d94a3a33b91622a6f515bfd39faed817f5d227654514c66990f1a2f997d1f882d4e2e00afc8e7325d13da2b50bde7033c3e6f13019e8fe309ff4067709cff63abc9676f4b4fc8937913f54ff4a58a5dabb6f2ecb168df1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8963a86b8edee7adda414791ad2ad0a20f08aa43082123516d65d214f1bd19eb7842a403178bfe8b6fbf29bcaea11f6784a8712365192d18ee3a3bc54262ae9397101ad65faaa864a82d6d39c6b497321837daacac4fe0bf351a0cc49c1a09fe16bb514a6fcf913e92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d351ba85444f5dd15081419f78f2c10bdea4ebe6e015956559e535b7088d6629a2d2009ce3833a6cb400496f48878544e376b8801f24065d26d0dd5b72fd47ea38979ff5696f6cb0e79bcb69a17026e99bea497732dee713046b1a0315f86e8e5936708f110fc4c636;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62d2cc6b26284e7e6b9177570d34f2b039e5ffc229b15cce61b03bf1a11095603bba80c05c41a317d1278111abfd2e6099a00e926826ac5aa221bbdad31c47d40ea71c0011c7b90206c45e132b44ebc133e4a3b884bb397804c30487e61fafed4a48fb7d474a1fb8da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5ade22d37eaafa07e3c37f271330dc68ac6c945ee307b68007959fe9aaf983a7856263b5a6b1670ccb8864322187e8de0834407f452ac40e9e09cfab92bb1a64288160dd870d62e05b7e1fe40da01b743a123131d6a0599c65af6d1547fd4571f2a04490a0ca36f62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b97d2eefdce91af88efbd53783a94493c5cb8b9704142ae7b7cd20c42b9c9d5a543750c2d6df519bb448be5e509693c36f573ca0d844de30cd4786dc7a4cb2a012920a101e8bb0dfcde09d01b6c3e317001700f19e7d172b8f283e9211fa04ae4571bcccc37c9ae5e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98b4da7ed666d257ff4c618bb0ae179c8bdc936348cf5c7bf503f0e963bc678781ecff12cac7584bd23c77d584311db92d7a562b5b855f670ca60fa3044e15a677e87bca7c0f9a09930bba4c3158ffdd87e92a74923cee514503c85f85bc59188cc1311dcc45a228f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12394f9838b618a70f3e144c6801005a2e61d5d66b2bba9d7dc2480b417bf16f5cec6fe09612b6462654549d1381abca79a03915ce98904a4d083205297b2b513eaabaa4e2fe52b1e02ad9e05e4184ce8d532c12cda3ed6e198fe95e3b78f65f137113995a5746dcad7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2d791f825cce4743bd525628de12ce1c23ed7da405a534976e9fc4d310513647b28f5f2e280b9fe4fcc32e4d2e4c3ac8a099cd0b61e1061d0680c359defabf2c521d1ee26e50fb449924170b81cc9ad361b490fcc9249a03f0b2289f1ee2043793c89e18279c81985;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161f2dae598ef49d0e1ca569302855a1bdeb6697a52ee43f7bfc3e1a5e097e8877baa9c58040fbc71bfa00bc4f7f5cc55691c402c38f8c2f1857d6b0991fd67e81b29c2eabdb0bcdb0d804f8faa1b845ad2b23d55ee38c92855893c5da7e8d0ebf8404f61bf3cccb2f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ee8a26c148050fc676c9ad4ad08aab3f30feff2c6c681b4a6feef9d1cec0ed6f3f9911768e9e7f7e7c404091284940f4054f06a8b99d78338cef4e8426abb0200036b2fe9d2f97cf966e75ded8eedbe5cce696e72790a2eb7074e9caaf578cc1293a87154ec5a2be5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17106c3d8c71096e5c18223c136b26ed42287ec462ba3d0af1f38fd6492947cc1611f90b811ae897dd8e2731afec41394c8702fb3cc25442bc8dc54cd5529e80420eea82c9721082c0d798c3d9e0c91de71b7f2297c36bc0ddac0536f9e02e0ee8e2d9e060d184f4592;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3fa94a3d37f19f46e295fa4cebbb2eddc721ff3ba5ea9419d43ffa0f2469ace2853a91501449c6463e344f4d9ec1c403b502524e764e5751621d4f0ead9222ec175fed199cd03c978dd050191f076b52a9e5b7267fb240ce1b7cee1de346784560e65d2d474d2e7c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38e67469664315d166a8c24dae142fba12fd3e9a533fdd58b52dfbb622d53a556bc216d053e2441a99ef34785f94fdc65ab9901bb66a81e7431b35da6446f6d11815a401ff2f31848a6e7230c74b4785f44cbb21c1a3815f5b51907d9fa5abac3b1a3b1e0f9ce216b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c711a18bc31321f996a6e6ff782f05afc1ea93915cf8faa847e6d31f9ef645f787bdac34b3fe32915bb4580f208722f03dcb9656e04ea5c0acf64046fa92e70ef888cd8a50dbe3f6f4d6c2b5e0023dde03faf63bd9a82a8a2b158b25043c07c855db986ba6e877ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106d222cf2766afb0badf1b646155acba6ea543d4e75b7859b6c4f9b2fbf2f6d73764e7edd19a14847e54e4197b7d1bfa0ae3fef2a1959e5c5e84d49258148738ac7d8de12e2d312708efcc1fe6426797880d90ada31d2b5bbb892a03d29963ae3b4546e4ab2f29c0ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1248ce99b063f39d42c3ad73b1bcb575f6cbe47e19b58484829122e9d2bf030223f5a2beb02907d8a9789a02ec348e3b42574e1d73ab083d54af8412988170e9d50f5570ef85593003ef369e62d6d928daaba28aff5d0424e808eabfc45e0fa97e125ba8a37276544bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c20b598b6098046cd271f0cdc1e28250680dce0ceec25bf57006dc8424ef7c22278e0aef667697e51386a3e86991ac7b921b3d373e463dcb944bb60b3e23e3fd30da332f88d940ebfcdd44c8fd8120511eded752aa8e2de5f6e58e8751ed3ca67d458a57389acd3093;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150188af99ebf30d6efa877e2c9204da669ee7aabbbdbccb100244ca4ec322fdd0066946bdb0c27f572af70d86f055db48b65e8a3beeff26c72db2cf219bd4fc3159d2f5343245510dc354b6d5bf2db746af9af547e59164b21c2abd37498bd4165f32b4d9bfedf7cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5c637db6a48e521aa4bf70937ae809af5feb7bd4e7c5eeb4cac1ceeec34bafe4b772451fe5c2d1f9112f12565143f02bdd012ce28c67049310722f84f6e8ea491f5434f43a4b79601b026cc320f7db4c65abe1ebdaf325efa1a52df771133477bc8f690d33f12d485;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3111aca9b72e0cbb1712f95659bbb05f9373ed4bbc57606c652c35ca1d847ffa6b157bd2f522babcfbd7790af837cc098de04102542d4b876bbd8c2e207ec30ea1fbb710e80dd628c5e43b609b069649e82cd2c2263aba49ed071172753f8c55c010e2b7b61e6ef2d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3bd98f6e3fa2b0cbb713bdee855b4788f55708c57b277a10f50d37b3e48c1113b918644b239da94d6385f8bef4f0cccfea3bf972599924b042d827f4ac689e86a3bc60fbedb30d9031d636e4e1c26e166e59bee70fe4342b0b4fe8931ca42fda7e144dce2890acadc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb7e5dcc47d6fd7997fdd2debc9020570c5a5a7c29a2c0b697d42375601c37dc742ec258af4ddf7eba235b4675f9c321bc713baf01304cf58a32f7a6ad51517944e0862f673cd9f4faed3984a0dec19a7caa615049c9642566b11cf8311945bf722507c5bc19b55f91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8aecd9980c489148db1c54fdaa54a3c24a02e544667508b16a217a333467b24af633f0990aeda809db8632cc2234fa2c55404a33ed80e49686c56102c86935e32d794f40901cff967e3a4395ed94346345089e3db0f8a8a9d00e349f2fd57bbeff4c2a825f50a1c6e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9f2a553210f661e086921e52181a2be8200dbfe180181d469b9e22afb5dc012f3ccd71148a3612da9bc0d1b2b35821ce385571d214519ba079adadc86872cf182da10fcbab3f824b74250b46cf7045974844f15b33b121616eaff0ce36e212f796493d2943fbba607;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f496539be3b9f597a0fee261edf5b5bc4a96b1fb951b2f7c6f8d6829def0d929ab9719c6192130a34a022baa5eff5f5a2506f310c3c8cc78bb066b178162bd08b67f98b2bd3db75cbfc4e6a12e8a1927c4305adc13e0504096df2dd52aab5d5b269c6401fb7bbee4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f9afcdecf8c3219d48fb46d9b63e16edc5de91491ecf43ab38e1e1e6579cc67c9cbcbaa3db85878ca0e99a9f642d624502b2ab114189185c687cdb329325593a11e1c1cc3a97b5700ce7cf106e18a2bc4fd17022c735285d8662f9e0d15f1af2e7891c64f9fb9668d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108a79d2a21b0acd764dcf8a031d80a5cc8fdc411f88b50d4cc22441663bd54e18ba7e7b79e579f81c5f6ead508ad02b8bc2d1813bd91fa6fecb29577d6147dcd9b438f13f80db42e914543051cd188c4cc612c9a4c7380d85fb696ae71faf44f6ce87caf29df3ccad7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4560f7ada63a18e05831d6e6e424a17454856b7bb4a49778230a687478ce6264b0d06444819023dae4dbb2230e70b2d50df524ee4c4b0e269c175071024dce27f38b0f7edbf642a4707e94cca9e05620042719eecfff915cdc251d5940601e519e053a7ba31d44f22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1151d9cbcb7e4f2d964b569bf79ce56260bee23c93995e4f3d9e6691fbd7a23aa09854bc019e6588181b9a54b89cd9d85a5a821b393c94a61346d517b8552ad020ba49c58c3b1b0a97858b28d9a0ead02942d123c9e6a370211e8b46f3859ef72217d74a16b93c9f2f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1100b0cad2aabd9265b4c1ff63ffd1dc211e91b5334fbc75449eefaa69f422decf3154dc6d0d0e69c6d3fba8b2d8c7305c366dab51ec152e99008c3c6d88e1c4f61cef45b595c86c65c77e2b25f6ff02eb8b13f8f0f750a4b8b1e33a50cf09f83b98b21612a48c0bfe8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf432f9b27ff3095bdd579a62abbcabda6dea3f8e1a7b77794d6b3b351da02bd0485cb19e1984e3dfd974bbe169429309c1c743dd8ef10dec1d9cfbb71f2edec516a0a17413fb134f3abb14b80220339ee2cc76562720773ebf59204652c89f67f76172033f7185bf1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c974d503cc30a46ce49d1dbd11e14e1d22bc66c7bfe0774952d1084efbb61d27b38c21dfe847058b55171506f16924cb233e588a0680b69fa87ab1a6d9fbb85c9146186799b0690862c6a6a386f13a014bd50f62301e00d67fb72b515f06b16a2f9f1adc29ea4322f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc590e400334731285a0ca931000fa4f8b686b33c9c8f137d5af23cdce1d1abdf902222a9b5e9adc93cc55fcaaea931bf2ba136cd235163f5e2c95195cb2ac74b9009dde4032f0dfc0f1562134b1c1dbdab963ba385ed34c84145ecb935d6b5aff1735784a92dd35bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2d0c773ef765e1fef1cf0f729a866e86617c13a8f55c125bf0b3e1e7e53ea0341c5890e703c204a098ec7e531550ce1afd4b6a1c0565e16206dd0d89749f19e1b962704649d66e85676a48bbaba2a7b9ef6aa27036dac7200cb233a17b7bf8050408a7bb3dd815300;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8624096070c40c6deee591d1ac78ce95432acea0627cd6ca61b87fd69f0c845afb831006e592f51b56558ad5179e6b093e4aa3d1a16bcab9658197483abc028513225f3d56fbc91f984680fbc7b98c3bb3c3c390d13ec376772dc08a553ee052ed4e06a27f50dfd04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112f28904151799bc311cf283ca9e23349d2e17e58e2cbe959544fb3a2a67ca8749f93ce5ffc558c0aab7b5d31d215c4a8b4f46b35838f171926329ced386d521227c657b53b8c290685983e7e7f2ba67544b5fc79577c31c78a53e3c9d0e3b8ae32f3ab3aa93ed5017;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h326b42b0ee86bbf70c83983ced2496d1218b21ed6a68b5f8f9d81268bd8314ae6465ef5ed3ed5541da896ee7ad0abd96a24885c34c71c136f6b589430293fa34ec89ea89830b43a0492595b7697506af24ac469a8eb799fa3b568ccd32e14446f76fed2fa48a2f4f44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151624f05bc29f88ac112be372388c3181e208b5f552d6814d6d76ac45f3ba79c4475f56b71a44ff2d2b0bf9ebbab4c9c8cfefc89ad4a0f696442d51a36bff9f8cab9f6ee14776fe85f81ea412c57d478ea667e5b34d27a49ec0fa9727e721aa66bbeaa67bb8218e704;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2a56a229ef738f371365f9a404a8767a11531f2671ab009b70acbab59c174caf2ee98f240b6e77646dd435b142a083d91a07ed717fa87e10fd7822cfabc5a524de135e884bbdca5ddb2802580d423ad1098338b34a5cd04dddf7107587cc499e98020ae447b57b5be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a39b3a46aff9bddf73d36fa0949a24c0f014e8c0581702228ff120c7a7b09b5713e62309902a6742d732f924de45b3c9a9f183eb6ff2e8686dbf7ec1101d4f17e3eff32b42e93b836610f8c868670a8db3cac0b9f4f63a910ceb76c0a57fc43b6058562586624b9172;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe2a0ea896f304f8749872809b3a14c3ba9ebfdf959e3b5698ddd787bf430210108ee776ada0b79f793886ed33cdecf08b01a1a104f1cd665fcd711945238a566408a0119d916feb251ec1b7b8ad295280e749abd4314abd0093a146261fb6951d6ac739aa0841d7bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h306777e6365558f27a123a58c72cfe64dae71746e226ca28d2de2f18ce42e1414c7698ba825ab2bbdbfe371d8b337c4fbc3f1ba140a414ef4299eafbced0f5ba2093af74eb8a6285f17453d124d1f988abf8725eb7e1a8df21faf690417735c0dc63fc623f41dca29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bd481b132e2344bc1d48d57bbbb214779492cd083bc35d4aa55b0833bea9555fb211a5df67f4758e714645d9264c2bdadcb6fcfa1722b21d73f07a8950de14d818d0e90dc285e92cb2f1fbf0c162cb9676ec2a9c018d936f302d9385450df669ec1e065073b1ab8b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec98fcdae293793f04de2c03d68a182ef0911a80dc035a49c45d64ab68fe5612e29f36a3d3ff7f70c2fab920ee49ee25982fd08a4eeb131faafc3b09338701f1bf3f26c9b98b692681526e878ff338dfe03136b0a9d98e5f2c25154972e7db6cd41b0c57a70a490d91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195da26467500600d114739c9ae8421562ed11f70a3998a16482b1660ea72f412afc35a92bc601fa0e20efb6fea44d7b381d74d61d4cd95832e0a5f063fd5e64270a335cc4b2b3ee8e096421aa594c855e15d025bf861ec575f3969be2fc48633dd3c4fb028d2218a22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ec74102fcc2635c76a40989d67c4deb22559eaefcb1027e52480c803874baa136703e1a521193e7731e486573e68e24a5fd1b2fc187b4cc1c40955aece470994d1a947e5be59cb89bd40547f2c45a90ed66add47ad6e6f932fe94284e5ecdf864e3cd6df35761ced0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17711b97400bf157741ea49bdcde8dd00d0b3d6c9b9a62a1b630d2db7066af440bf6de7149e8a74f7d9a6d594407b0661b7cb07f7c997923bff9cd4dd337584c6dcff1a92eebd518bfa1a3f9ae3b0fcf38b92f1932287b68b7d4fd72e91da958e84b2ec98e0370bca6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a7717d38415f07adaf11969b0e94549ca9577b01e31d4c4b1b69a036baad38a4ac8f1125df31973eb0df2430bb4376e4f9e80735e30c009f6b0283ecf0fd41eb860f7db67115bfddb820c6da991ed43f25ec7c0628144183ab9e4cf764c95258ab2d5163334ea7938;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e9ede63b0f8e1e7106efe73cf7d60828711d7bed023384202d61db12a43dee388ba1b12659cbcfa6063d4066041d5b1aa6177c13809a8725aec3a7bcfe71f6e11c7949b109643543b3e21e089fd47e17e74171fdc45743423baa03ffcc07cf43bc2f9e6513e1b671f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h794569e9e6236ac68d3fac342469141d4899b715353ab842a761288627efc12936534bfe6fcb0398a6204f2b35b42ab47858a4ca0da2ca922a857ea26d27f170496dcbf26f30faabea5073b4a12f27702caa41bf23e5c2a03a36d3f89da0261b7c0199e5f006be4dfa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h839d28c6906b46ee65d9a9c277a4e408a23f2df3bfff16a25618f5e4079ec8f3e1e407cbab336c8c45c135b70ea12ad2f0fc527d9a583f7bdc065975004ec47f063d7c0e1b329a1afc505ecca7096f98fa105f6731a6142265136a1b2cd902c8db317000d0286a4d54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134678220eea9ecc0cdf8225ab01c92b8baea5a94e246c11ada354edb4ed077f40d0a508ac4b2a24d58d8c0b675d3e9ba2f55a39b820080633885c1cbe60752de24fed3a270b80ccf3ce6f636bf2664d1212c87e91608927fb0e48acc3dcb3ff3b83b6070cd309017e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d81e90b63ce30ece17ce5436f2bd069272593552af469fda85436f3a49a0729b3f33acd929578e8a9abb80df7905bf0fa3847b1f273d9123b1c317e00614549002c791c1a7eb024b7de11861b4bf02d82cac8080d3a04de55c8de0c4e7965d69c0bdaeb68325ca062;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h581201a9c9beea8b64418e25a939aed7248b1ccaf23062de93083484ed3e929439f5e5cf2fe93b4d57c5e7f0163b2a5a6504a14ca490a66cb08e1d514a69ab451bcb486dfdc1ed07cc518325f33df166e35536c36fbed18a8abc66d7609e83c2b365577fb992ce120c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122f0f39447ae739c889672b51fa4a894fe38a932abe1aae0616c2506424667cb95190e63ccef8a1c710f2d4997347b8dbf398c40cab0676d31245490143de358054af00a0354fb30b6c98ad2f0305c1a407ac9d5a87d9ddb8ee058fc1b18a188a2742e997ae07459ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e968778a4f6ed9720ccf630d7fd68380f06dd947393c65cef6f53f72efdb612d567d4b99e6896eda1482d0f8f46da321ed73953b93c25002576869d8ff0c88b3c350a5185412981cec170c717a57f9e26e49dc5a3da75b5f41d859ae607771b9eb0062e82692fda0c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23915472c8b6e84872e1edca83f063cefe9edaaba81bfcb42ff785a226dc0cc84633c57895b6fd0abc846b4692cc77b8071abefb9e6331d48fb2de7a6c2b7f9c914f22838d8661d83850cd220584b7b342d108794b8a4270b5bdb8a04d7235fc770d6184e916a29d2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a92f7e300f0205efd3017450a516acd564f2d4008d035f0b70f623ae4b9b84375cf1a3cb01b389e39de9ca5485051317b0dff6f641d33fe9ff8455ba7636ab61e994fdad38f003e723cfb0f6ebb8afce6dff36de3737f98dd1ba0ea5978365047f6b368f6e4e1ab3ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d64cd5bab2678364fae6a98d41a03a17437ff3e3761198b555f8bf4b2e1fd8a18036b58b167d5f68d3a7632a6f2c7f8ad6f383affe2676c2bdefc58c00da866094fa58472b1cf589e6be7ae65fe272f7ae761ce53aac33caef726e8f6a3b03dd44257324973f7143a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fdbbb76951a5222333f07d7a71127ed2c04b89e9705c924c624e92c89d25715af42ed8563f6121e6fedc98ecbef6931d76d59667fb534343ec870f83f26c7616653be25f6e188b701cfb5ec51a8b012a0ee7210bd0012e602d39f8e250d135ee21e0c319d6582b511f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148006281c46e86c17b36987323af78307b96407d827fcaa187b5a6257afb57d3e637a9a1f9a2a35a65d6ae4535508e9931b78f5478fd0f443651ea4bbdf9cf4080d47ebefcf53292de82f413f23e944e644e1e91d974e56aa1271db49f7038d4d18df3c6f6b00c3fc6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4985e2c599b1c65620cfbf92063324c21333c1da41cf1102fe1c16455db8c93ef7d11bf6b382170fd0240e4614a94bcb3e2b054c822184ee1ecd6f0e41aef46f31ed08307ed3ebf322b347ce56442e297308686fb988e6931c41d98585f44f27fcb60089683a81e08a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c8f411bf35dcef532d5fb49d2b17d4bafc61301e264302b9298b024c767f6e33355e0ea196a63b65cb04a124b9d833b2f3e2b3a1e6d06ab1731bfaf0eed0ae8b58f437b70f838177717f46a481dfe92f133625be65385c66be31491693e14352e23248bfce75b7264;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31eca86dd23a4135aa467546ec15e35579adb9cd6e4afdbc5e371cd09f6e6da9a8996f3a60cc979e3caad95bfe583297a024f67dff8b48d762a60631b931197aff40e718d51047c75eaddbbe036d140e1c31a81b4753ef93beeab5e1af87a048076784f7ddc74c16b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e80b6bb548c95c1db65ce24a1eb7f543748f564512cb044ead6a36e388eb5e35b4d5eb91c7485fc4f7dcff824ca374885dba1c44bfd6dc255808178fe47f1830be34fc4df60ace3d197b3c98909df91f77e458f410cef6fb635114e16583287c6d53a9b39191d7c56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c62170edf55d0823d1c451e398a9da3643004a73106fa58b045acd76e3548f208f8c140b30b4f14da970c80e5a7151f62a130ea60b039010ae410fb488c6078f82b9a915301a5fb1d8f16063a0ae49eb0688b748517a81dacae987ae99a64b6e73bdd63d3a354f2e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e32495981cd8ca2c5eb58b67a6e3719be3ae8fcfcab9f7f5ac046e2c35278051f4c7d4e53be9e3a5f8e82db8da5039adf986fbed3cf2d2b246112100e21ac259fd9adb0ebb0a9f7119b8bc628cfc2e88f467b9ba0929a7b5ac9b18c089de662d6651763a32d00726e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fca6589688d153d7e26ae18a51c057f21ea3708df360381191b98b4275c33f52bbb69790b84411e91a022749012a41f923087e3c965001b5a26cee57f6c46f303d7e7c09bccf8125af8186d385dfc52ff1b919a490aaf346bed58b71b1717e3098d66a628b568d734;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1549278faee9a648fb4479b3647c9bb2eae6e1e42e95a88d8f272627b5c17b648f2c2c2fbddafe8d0d97166bed73f8cc019e23a25701bd16b725b7154b1f658ef800f799c07917441723851ad5e5e0ddf0fe43d51ce5047da1a392d005f6c5989d6d5d0bdb163ca1271;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12321c7625f8f071cc7e15b42f7ea56e776b432455b3e16bc3cb9d990bd54f7d60d455cdd4626269bc26fce0cd8bd5217551472992089414f1309f580c40252db83b5ce8e26f35a739c9bb48b6303580beeac1881868bd5df59d04e0540576ec5adb069160587e00896;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91cd21dfbea795b51b06f67e0da59a7479818dccb732716632780d4ce5eab630d3fc7c49d6414a38638a45f7d7a7d27d44bffbc1ba2a5019dc44c6a89a4c52509b5f0ada007eb5d680d0808f241b1f539dbdc4224b02d0b85e8a0f03b3a27a7355713b91ed06812ba6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70352da80478d320b61df0924689efcf6d7c8fbffeaf53e4c7ed239586a571513cd17b903afccfd336233ab02bdc916ce9e5281f176b3c3dc803feaa3f17b1a52cf540136c4cb303268713a8b0f4cbe1bb78fbd50a320190ef4812c98a6c3dc29a2b7d555cc0d24a3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f6c8c65de464cc8ffe51d1d5c814138437cf734156302bf9775f3694d3e846d82446b76cff8a34cb85f1153305815376f135c0676a228ef9b91d34075fe0b1bdb2bcf71297141922a1c43c3b201c9b7f3af36f90ed31c43b417a967d320fbd1406f008488d705eabc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5c80b5e8efc4513df5900f614ffd692e85a607951ca5e89fe2df6203e2db42ebf1f0808112bb8637a897819cf7cd4c2ecd47f6aad316c3a014d063a49435136cf7d46e423070d660712fb376e12ee40ee6e3cf4dc31b47ffe5fa3a9206d953c80b6331721936649fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15312e9c7632f05112b9266f8c1e850ec54534acc0baa2d85df5cdfd558c8db9e4bf9c512f343e6eab484aac61037d5d8a31a61caf810470eb7eb47bd099c3e9909aaa26d808692dae8d3a364bb9977e45af7b306bd8aab7da0a370a5f35b93a609b7c7376d80ece0c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f27173bab4442b58573abbea4f7a750620caaf39260e3d7c60a1c21e6fa856c049799224f443a43645c49ede3925f7f6e47a999ee1e113af2593b681379106e5a8b2ea2a461d777996df3bc7dc431d51a1d2276fe632f9914bd4abc9e946820092fa2b622eda14c45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149cfdc77ac2bca95f074d4d29a88212a8f3133b3b678bf46905a315cb6d3bca29a5f07b7f547afdc50a5e7400cbe0bd2515817593781dc3f81ab68521b919d7e0191112faf39318fa49b8310b4206bc61052b6bddd428bbcd47f4399a1bb22bfd21c1dcfe3f3f4f965;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120e8b034ea670e6bc32204a25961a239d1d5a6c98d96b621cab3cf1e0091a2b423a91d9887833b00e2c7411da5ad6ca47e7d2237d33009af5cad567004a7ffc131d5149793f0e0d434a2bda38019e888f9b3abfe5b49f995809cc2d4c4152af9452bd418ec4d2ea9e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a345c8f3b47e26f61f675f2de763cb00bd459517ff7206bd1f04145d35cb3b6ae2a5e9fc7744bfa11d642a28f150af12d9148101457ee2ca1e0c675726bb608631aebfd1fb711777cd80fde50c80aee35262125a8092cb090f9d4464c0e1910e91c6cd1661f0ae93f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142257b87af06d269332cfae9cdc89a5fd655879f1adda01478eaeb990763589f72a1b2f3b36674feacb358d671956101d4fa362e0464bb33c0904a7c7c19c7935405ee482171c10e33df3c6424358c250d33e159f156d362761c2eee077660e643be6aaa7107b47188;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h728165992974f3348b03e39c6b5ad86cf3be1c8a535d43a153ecac4a9170034397a4be540c167a066d9fcff5525a7ff282d14811f012223e5df38cd467c6c96899675d713ecc663a925322bb6298a698dab6d972c98dcc02fee432ee022f33c33de5a8ea1932f59fa2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ed0e0a8e83308e07d710bece06038a01a070b2517caac314ea3068f5878228328cb527e47d09e23b7199a1a78ec5291f543fafcac130171acaf1a90049a19104c4d28040e3919cb9cac7f099d3937334238fb73bf71ae1fcc469639425ee3b5ec91749157bd929fb2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f58729e80d4e478d5657942de4074658e06f002b86658b999e113d2fb3aadb84baac42be541d3e921143951fb17188dca1a3d99cf122e385d883b33b865fe09cb72b664e3ad112eb8ada37eb1fff013f7b391891173980133a78c58db0c3b665c2e945d41dee0a5db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b6fdd11485fc547685f00af44da525a22fee651083a91d6898eb4ec6c35376ec0671a94759756ba0f1149f34409a8fcd85e308481d390c40e87bed8be30762e5f92925108ba869344978be3c5dbe86ed3ff677c8ef2757ac552b34a41e4d17f117fd766b68c8712c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9588af3ecd4cacef36cf11c506ef1b8c69b23cf46fd5978e850dac120e78bc130c5bcfc380bc58ced56be0c195046611cccfe53b815c32c0adbb99ea212041c8f8779c2f023f46d97217ca1ee500448b128ed19bb935dea028ee250140c451940f68f511b0addd5ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfa88e14de612b7ea17ccbd28b09b37197cbb3dce24ef198895cac1d026623bea0ed7f6a5c01a49bdb83a8af6ae7e6b3a82067b1f6ec97943b47f178af52ff9fe7e269d01e8eb164e2e45f16b5e42778c2db5f6f74d4db7cb435c0e4d2d5ec44373c9cc849c8283df3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7bd51ce8679f5537e5e94f78ce791d05857a200fca4d24275027123902d156809ec91f1a50349a595d246033b1bcbd6484742e9b98b7bbb340ea484b4373091536594a01a67a0befa85e319ee5708ec5b89d2742384f99f5a6fb7fa498471450e44818b12dda9c855;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h270e0ca23faf13e0cf89162351491e8a82fb6804929c3627c42f0901d28701e577e5dbaa6b45c70def42d4b10bb4a270d0b85a9783ae3b831fd614a3a0fc6d0c8f7dcb8413296fbb1485048eafe12910ae9f32c59b12adce0cfa13f328555ae620ca9f6dbb2eab9199;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81bb5d359ea43d96795e677ee30702e6c6d83c8ded797b455bf99ad4589baa42d9d716ab337b5c20e68fa2b3e5c3fd9ff329e8cf8766ce98da4f811789d5837f25bbce402a9ff410ee0ef2563feff3290fcf7daf5b31a73387184f8d26cb72a27f47ba6f20f959af97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77862c4da5a375bbde7bb7a381874e7dfdda3b7430c912d0666d673e83ecc301d1210ab7cd6d22bc77ec87bc13b3ef7b88f742b1bc1452e1942c67a5962fec9eaea7b15208a45990281f10714319322dcf1afc7d828dad8881498213270facf2a3b4b79e850c9da558;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36cd213faffe58e8d9ea4202b2ae4b3642853ec1037d6f01654d0661318a442748290af57e7fd51ca77669fff399fdb6d7c2f61a68c6c0c081c797dce31d572a3633af30918a2270281c2dfb8f516f9c508462cc631ceaa4b5940c56671f0519f7b6c524dfe5f872d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he55c867d85a67e39f6eedb027a43abfdd5be07884aab298e9818c728d1a492b2b55b74272e022f82e58ce321c6b864259a626c4d5e8fb8337c6d84546d4fb16dc096ce9d7981f82f0da32f8219dfa5826a6be72bcd62e731e03f15013c04da7c99c7a66304cb4c4847;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54bdcb388e2a0b8587c5f349e80b5d5336b1ec2fe96e735f97196ddc2e14ec4f60e9045c218cf40cff1e1c306d3ae1297ac98c9777bee8f2a61670e4702b7ae56a8beaf273ce092077b7eee62b94977681745bc79113502d30636bddb66f450b5dd61fcd0871579d94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha02eb4c2961cc77dfea8cb3c8f873acd0a0eee505a1753e53ba5ced02d0126cbbcb70fa99f58e3dc2ea8e4c35999b26daff8594977d86120b1a2b0e48b4a0fff90f341b6016d9207d810dcde0f5214b20a2d99aa803dccb3e2b0b6bcf696566315513c7b6572a61658;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef57047bfedded26778472eb3a5c1d79a8de347b174cb04fd72bd07b5456b97c77312478ba085af998fc9d651af5653cdbb9728d88ba310aad0e16710d57552bc11a5058171cb7a82098a27a1345e2579c0ce47b0a4ae51208d25e1fcd9c20931bec8456ecc0af19f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc67296d4eff1086028b121e2a0434d1ed75f887cfc038138b8f71b521700cea21f150f2f2ec1ebabb577c4ef0bc1824a87f9aac9eb2690cb81a021bf218b8ce400346ec47058f50cda59bb82eb286d35286fe7ad60ea193c50fc93b0fa40815dce82d8666cc3b69373;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f08b991338edd71d0a8b6129adc0988d2cf95ada9330064da9ae26cbea691b2f3ec02d6bea78c8c87c9d0ad777aa04c5fb9e845fa1cb2a5d5ccceea67e8581d9d6d359e70f2e6bb7688860ec1fd47bd406a15c323b66dab061fa2ae9796b0bbefeedbb0702e192095c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19520f4b36f3e9648f359e7558bb780f5beed02850434e1219056f259b3df4c64b26fc8ceef02291a582724154b74beadc171a3543e70c59a30779653d3e20982c42e69ba4975d220f5d578d6b89c3c053635fa4c7f01eb9a486da29798afd13be0c5a8d6ff45a8070;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc40887e84aaf52423c0a9c6350da21e6edc85afdb4e2e6f72ee9b16272383c83aaa6f911abe68c2d29cf64ebc437e02835a9016fe3be354f35bbe596d148742a079cfd7665be6e543651d90f9e55d2c035a6a31f34d31938486d61cd3486a503060490f029510b903;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5e40680bad41eb0f3a7e003e244208702f8a384c7aef31759e4740ac0c2af43098604815224dc95e21a126cc254b8f78259c20f33e1dd06156ba6126262226915af7a969a5422ad0115e6dfa1114606d8547c525157a11878149b58947d6074e76081a66ca131595d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10786b067c4a6a9f14b71005500cdf429a3e36b99b7c493133d0421d6d603ea7169dc9969404daa183214868ade85b657361b6f6112e47d0812e8a6d9cf871c97b7898cccffec0d2cf01721d1895bb36ea8404d9464435c06adce0f0ed7ab9c738872bfd01c9ec0bc03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1daf2c4da407ebebee421074d396c78c8c097fbf01846b64dced27c4a112e2d9adc0fcb941d3a729e226d3a487ecf03a0c3a28c92729a557bc0349493c7f64d8f52a0f946b33514b446ca6a51e818bc8cdb6bfbab1b81e7499dfc33f53a1a41696884e857462b50e051;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e7370baf5e18e4032fe1cd9538c387852f69ebfee7fe66f221a6d8ffabce3df5ad05e5a6f92f9fa0942e8f9c1e4535f0db38d99df9179b5ace510de2f917e6d5b75fe8750838f38147c798e7d6c835d5150db4f9a08f42a974e15653ea0855dcab0b168a358d2bbd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c69c568afaa30011297e1323930d580018e49dd6b6c50ba60de7a7888b071ba61d7b60cbaf14ccacc3b66e25f3bed45cb246dbe1392fc89dc120eedd6aa3069d7bc32fa1a528f02d8dc76a4102fcae713a1593f28f28edbd5aac914b2b6631bd127e11493ee4854581;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b6c36ca4efc226c6b2ab6b8a9fd190eaa98b172c1e31f5842ad9ac1cb3d9dab62e1710de9926f73eee4b7d12838e8298f427f9f807ea63f5b59809f581c1f7b0aa8842a2dcce399434ad5f6ac61da519eb8ba3ba6410b326be5e86a0de32967b3b6adf226f3798e9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd605bef4e5281add12df7d825d2bd4a8d43036afc42270de2563f303091c0ff541b667cc4bef6ee99412cd217615c74557654835d9acf60203626c784c6fa3690a975abb6bbd6bd60710cd9b4c8261d8da0ef9b28ec13d64d38c471fe50fcb8d0a90f7deb59253a3ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1358ec1dc207f6eced4b22173102625709f1f8de5f2d50c6e2beafaa5040c13a978b7fd275570394daabbcb63fc51a4b146e97599a83345e0a73102c94401e07cd517c4c6042d30fa8378e259d83069ddc8f4d0a29b60f9e7ddd19b14c5a28740f3029316df1063e727;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cbc3a27541a851261e4eb44fd56e8df0025109f7d2deef4f01b062543d9007dab90456b68549f0517569383bed0154e27d70e6433c04f7007f172423fe2510253cd0ffc7c7b9171a37b32e91ab36652ccf4792c0f1e47e7fce4ff2a6ad6d3d046fd606c763b69d561;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0f9d45cadcfd947b27491fbe54bb9f65ae6012e5a79a2a61d46b200f5bb6f94dccc3f3dfad758b573bfc181930a0f4abccf62e8be6f8fbac28cdeaa10efe41323ef96279cc54c192efd1fe6ac17db037377238db0d44c589907092d7eef33cdc6c698951d7015b482;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f87ef16f46a9785792b4c5ac771d243cb46939b1a2c7a1d3c0befd9664532b52df7fdd1f125da321f3edcc0a6b66596c47b5e304c368ace95bf636cee41a97c7c127ab0c548788cd842da5bd1c8c73d4119faad3d34d3e740beafd1311350dde8bdbbcb6fc41566be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3909fc20607da2a0759df4afda7786a2ffdaabc88751818c08c04f7d0ed40662782093f54efb79672cb6394e6b5198bb648434e6582d7d19359f035be6265f48864ed5142d05827ee9781db925429b015f8bd8dd8c6f1b6e2f29748360a24478b1b4e10686aaca4fee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc12b18d10dc21c8cd1004be9f0a23836e8739b6d070891645bb01120b94bf661cefe7d8efc18f9cd8b5bd7c0752ad0e0277fd6273dffca2be472a8955f7a70f29d4eaa3a27b903991d4f905ae728e71ed3d699df845b42f93409ea52a6b3c30cbd10dd9bc92addbf11;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e03df037d329d85574c0ce0cfbbf40f877a2f0ccc5d74af7b5b9f8abcdf63cd0a3db62503bddf94b207123fec45459bc62429ded4153d68b0095c5151fa3880787934e5b14ba70dd54235e69f45e82b94b8710e3b9510add45ac2a7924c5c7966fbfcf5d4c9505028;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1564663d2260dc865a2c526426b55386c6fcf4ea1fe08f659ac30c8f352d7fe1f8bada08bdafe4de9cf247443a4b902f0bf5a4a80da097fb49cb10fd3e3bcdd8cf50038944d8fbb4ec122518c608d7145aaff1e7dd1cb8f2dfe4ca8d7a67b68a8653e716f01e6919896;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162ab4f339ea0cbfaaf2e26d768ab7abea4c982f14e0e262d0d7928cc12661e9aa64124821ab744eece726fbe88bc6dc6e1f14a6c8167b600d3d7c9db0fab8a7ca8ba89fd0c60ae3e0abc68bc9ad0bba140d1a938690822bb498c297669a4d4248ce5fc13fce13c3a30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1131c0656597caca28ddf054516474bf7092c4b6722bceb819a2ad6aa939d7f93ed6a5a1248a2ba9acf5b69d5f04e722499c8100ca101157cafa5ab0dfb08b80d4e79e5300a577ba98bf2e5172bd0c028deef35816e4753ab3a46b40e242a6ecbb2e657e6e47140c718;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e5e3aa41e349210f608893befde8d10a9b8b986e95f3b4eb1230c8d1417616ca8c7e628b3343a6d1ac8b900292e473706ebf662b4e9a006bc80ef505e0d60a7aaa0f601d7d2e59d7c10fcf420f7ec02422d1666182fb0134f7fd25a651d17d04171f2c6f13eb49770;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74264fdc9fcb1314e3a638d0cdf83065a21fee460233d02eebe60d1a0fed5fb370f7628afe54ab9a2095dc156590381ca697b9a55dbda381e98c195cd7167bed4ba4c5fce65e20cd8f8998767c6106c0d35a2e3a3041f88b21345cd08fb09da79a76888d24b91b0a55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108f02ae82f9d5613e3f5f66bb3dec5725af8ea98ff063606741154f77327d7be3c22c52ee77df52c018d11ad99a25c5a87e26d01a8e84410c4891dcb73a6bc27ab48b985618cd690619e5f76ee8925c746bf6a149119ea6ebb6549f28711c7b39f82b3c952aed7e385;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4f7610a934da71eb61a3d848096b4b232de822e0356b5217dc75c17c1daf6422c631705b5c4664dbeaa984a70b96cb32653f6180643e08b3c70f1a3af26b417d584a10341495b04016ac594b7f3092b106412bd6c7da1d1d461fca496e7efbfd10c9d191488749510;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f3f87d2bd86c8c99a2b491dad0a87e8e23da976122f7496c3f7dca2f2a13489168b04028d6796af10e1a2cef63c03f176f456f52b49259428eb39bbe0394b1bc105f025c433f956bb10571b01f9c5daa71df0bdac2a9ba8567a4d15fa3cd6cc198931e062725f91d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127c1f470af04d794ba49b1e4028628cb8a808dc4b600413ed9aedce41e50a9168e8695f42ac0ff54dcba67ab03b28aae3dfc870441e4de41ff53e1a30bfac09426cc4418bd874ee4db339fe3fa8353057757f476609881fde8735737ef78f550836f7a6ec64002d252;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dde740b6b7a1c0b49efc3bd9391bfcee59c61503a6bc8803a0c7e2c22d5fdb2385bec9e27875390068608934bf85a534e80adb564af00f5f4c40ac32c20238a19a6e54d3a45f7294f8b06f8a9f94ec586a45409efc1cd3b0327dce592205d2e9fc9416eeb1e371a53e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e2baba0c7ca60a2c8260b43112f7c16ea71254aea7b1bbe6fe7622fbc54dcf7e7beaaaecfd47b926e8a7d4d93bd2522ee89abd30fea4eae0fbf6032b13875691fbe6d15cf60a387afa33bf4a6461a8292fb51ff71e0cea05283ee3649aae36280d5fc2f0051af6aa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha03391b2197f5ce06659281b38faf5df1b4e8860732746adc738b79eb7adaac19bd267e46dfc18a9ec1eb7411ae4aaa00a4be972e93e3c58b8987ca668988207f74a776502f18ed579b5b631cd83e56f53cedc0ee3839aab98ac9428c077c8f4afc4c60e89c09c1e2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he66707b346633cb720dc3baad6e23bc37bb3d8b868e5416ee86e84d2ee6899f24c185572f178fc4f1ed5f7acc8993fcea92d209725c85db66bd32214adcab70b21d10e126d82fbb3431328e9ff3fcab19422e18c4a78ae3205310356fa12a4efa1149148082687283f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165999fa6154390afed17765b33fb1135590ac44584377eec49a6cddbf98946fe729d94bdc5b87fc195fe14788dc9bc125cd59fa6217b674a5541e75d1e55a2e5a5e5986a973c383afe951a4d03b0672a3e1f0bf9c918987c1ad9b6f498e2db475b793d6015f7cd2a39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e5d63bc71bcda21246596a54143106efe6784feecd0dc0df1f14ef686a1cf0dbaf4cd0fdcaf328b728446b1c9a96f070fcf946f4d783b2b64e4bb41385905d5aa083fecf0234eeeb9b36faa5ed64b1db8ca87e5ca37a3812792fb310baa2d5742da2f169cab483693;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163a8d1797872cb44020aa14ce99276d3f4eb03c4dc0c4d35c1e9840e1865d3b16600e22a5028cb3c799ba45c770d4ae68c7495f7f1b60eb343d479a97ff81188143bca88ceddad39c92745e9f2d1b8374e71fb7807b151d331151d9eb7814bfb157434c3d0838e2bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d1bd3393af184cbc13a7c282ae73820c3fdf46da456e2670505397c93f2b2f3598b34a2f697313f47d1201cfd47f34b94fc43355df24582f6e930f8b3b8eec118963dcd8904567bc648913701bca5c2d898494c80895aed2a6b24f39ca53ae1b3d300bfd41f23e67b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d56545cf1d843e77a8ef3a5ab7e73a7fa620e8037c6de1b9ad3dbb3bb8f554132af3e4b1586c6ad2e367440a72c88bdeeef62ecb71b9eb4b607c01369697f213899fab47e70c936b2069423ba95b75d519c9738e7f630cb2a4b9650f81119b8fa5300477043014b641;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18558945b2cc857cc47e16b6b3e60ef14137268b228392e84ba5fd4edc3289b25ef47e577eaf985515bc9f43ec9f51b1a91581f4149f03814a7bf6b14b403116571d7037caa7a38021734cf999834aaa3d6a911db0f188c630a7ff1a0b495c8a6ff1019c94d64949848;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bf968760535a90450b43eeb625df9dffe52189ec029a4ba12254b0cecaa952a2bd3e83a7e60199d07f6c30e2b232bd212f1bf3949389c4b956c7cc278dc227d3bc2376d2b0ec79ef5c8f43772ab4b7bd7ee42196c6c318eee824a84d28f66caa22c2599ab4d235f3c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12561e93efb495326c538c6067d130c1520e542282e41986bfce74fd46b52dffd3522a196b817130281c33e1be1c4e52f62a45259ae3b2a39da3ef9ae6e93247e9a827043fc43c87923b4dfb9f48f370fc52e1b710df64700cf55f4119f9029d59c1f5beac40f725e14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18490e39a59618024d9804fae0984ba0c2d907498c6ec2b4117f8c6c0269d4d6ea9fc2f591614d24f1122bbc777fc0cfed1560c8b0cc4660919b13b3c97d528abf1393ab26173bb37f85531bd604f2c1497afa2c5cfaa03df7b02e265a6db80f803789496ff5a26344a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5868a8f1a1bbb145bc4485c7b45cfde7c2bd89edd1f38a7edbb31c4bb56b2425407d917b8a7ccacc946389ffac23d068f574bf2d00130106195911d5d37a56eb6edd7116a6457235c0507909e8b835d0838849f78b86ac8592a350850c5012f9039126251df977470a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fad665aba0a2c551d457a3bd034038c93de310a912313a140f209125280f449f330e23ebdfe08508b84bb0a98b56ace9b0d904db3167147e443e78a99cbe35932e8900a644a25925de8d65d202c6ffb1db3198f96b88aaf36329daf1d5fa45dfeadeea6f80d3fb43c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a2bd897f30641aa74515f184731c63ee98bbb621250d65da78e3a7f0053ce3fa7841df82e2d96d2cfb86542e980db84d7740541aca4201ee28b70aa574eb8b28de7e0d7fc7ecce0a128b9686fef4048452bdfcacce6c7a665c606fa5305b64ead9662e8aae464e7b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd109c3b4dde0ac5c086c49b2124f058cbeb5e31f5a77b1252b864079ade29e7e8ad37b5cbc5d9839ea994a6c64d2306a6fdc80e27c7439af68ff367697ed4eed72507752f0d6cc796edc3d0d60a2d7f8dc8870f491e0541391029694aaed2e4c39fbab5f7f46c2b354;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h330b5ca985273054258b58c86a534a3612e06af3063728c3c33a0b938a331c49fdf7150f18a32a48671a81c3b6b09eb245add7bacd1f2ccc87528d4d3e67958ab63f818f63a85ae6526ea3b90be26b03574a389e2c5bc8a24bf78499dd0db7e0cab4ba4c49bbfa028b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b25896fd199783d729d0956ef832dc00b4b1f2944c364aaabd1cab7c67692a87fe307c296fa0da258aa997d31a8394f2d0c8fd8edf52e5159ec6098621245bdc7c6cbf8e480e492a8a62df54050db3a79293bd05d928a192b971975c31fb1215bfcddaac7ad4fc3db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb517d69520a782d2418bf884e431365e6ece5583a7515301280cf74f6952bedad575584945f20be41879bc1fcbafb051e396dd8cb5e521063313e5dd944da7b25b51e0d1b21180a9819adda3c97fd2e7b39cf18277af73ce2f3b956240e70f119dd4eb3551c0d0587c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9351759abca2576cb1db891d58a16808193769688d89fc99c550f1a41e29b7605e38c98643da1508bbc755934518dc2e41200351f7aba4c052b5a37c49a86c7fe938731737d3178752880f152cc7ac1a2b9576eeac6a7761509a458a77c8195cf5379f1b89bd20ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123a2785b1b491519b08515af4fc30699ebe6ea5ba4ab02ef1128b0003351b9522a99e4de166e273a86f8d9225d5409235fedfd296027cffd74f3ba9bca9077dbb3ef019a5a4e783305d3686f206d26a9b68049447f155cfbefa834009a8d064ea74061e4e7b336d8ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116aa0fa9c9d26eb4c37ded8e951746c2668b60794750fba5543832bfc02055c6b20a586d1594caf70b52853caf8bee6fcf8ace3e033eac5de221898ef30f3f8cc9ece577bb8e09ae9d6c940011d3148135e82ba4443333723aa1a3d8d8da8b63a3af1bc6200e61919b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc045604057676045ad303b1876e54d226e3b1202ae41d55546a740d37d277fc4b34eba8406af743d71461161e47b8c441eed2456f81c1e2863e60d1410519ccfe7fbefc3ce7f4163cd919206f6d7f7dc654e9f2238928cef891563cebdc9afeb8a04dac8e6605673f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h938dfebda02dd7ce71db62e27a859432b371ee07e33df2ff76320cd7fe239b2222ce4b0ade19a9e01de5dad0229c68c88ebd2a07d5730e79c7a34bf598dbafd61980823893120b1d4f8ad03fa14dc1df48bf437f0435887bcffe5ddfa81bf1e8688a187fa4575a4c92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccd38d1b42bc8f3d65d48d298662b583e952abe9cb5a6614bb9e8ec6d3ff0ef835698d8cefb07112bc73771d94f68e64b472cdf79db9aed94cb39f9b83284dcbaff187e142bceb5b056ea9704e5fcba47fb60877b654c746b7aafbcad3649f8b99ec547cc5a74bcc60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0ebe4280622fd42ff96fb875ac4cad20fea92605a4e715f5cf9bb096adee0b14620556838e142664da55e5892d23d34522486468914ae39f6e180a4720bd6e7befe8478d6e87f8f1d882e6cf6fb6c658a4de0cec6b35a30dfc678311f59e7a82d62a4341152e58d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7e7e98463914660bd70ca174c1de3bcf9171e7fb82640de51eb776d160f30b08d0c0bc9ebd185270dbddb8b4e407f5817d5d80f75e4c636950c864d07b7d153f6cd46d8fbc42eda57b19c0627a3030698842e770331281e31ff58c4269b8096139e83ea3dfaf41df9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff261c92e0c98ee48a8ee95982a847b819b8b1b8a474c3138255a7cffcc6fe0eb59b9a32dcacf30bb11190a246b8cc6ba038b8033119ee70b77500a2f8283b3fab76f913939158bb1a78963dfdabe019c1a478acb6ada7299a3155815a1eaf753fae0b044806cb712d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a2d6ae9279e0d7fd912ded5c118832e72cd751127ab9df4f145974074ff846ade9a3aede7e00f85f6ce3b99705cf8bd9287de1eaca550fe83f66e4e337379338ab4d890367024da527acb2ad4e5280099cef32a6917d4c8e6780211dd78a748ef1a53c44fa520d3c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bdca4ddf4b4450ad2d7275c88189bfb99f864fccafbb374812825036a85451718fc756e372e6debaf25484f5282c2f9e9bf397bc2435a5a84a0127e3b291fe44988a41b84f5103d1731ef8c7330dc31a363f4a7408628b938628d7d9e0352d02602add08709e33d7a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb40309b0e1edf1a509da5ebcb647693fa55ecd7cd6279ea012b58358a5a7af48f31f7c10daa74dc6b923500283b2cacec7d344d0de08e65d145c2a823dd3efcc33f15214ae6f62c28e6521db14101f0511da1ec643390e364c89934df12edcfddb59854473873af91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ce1b896c91f3317a5def6f4f01a69632d7e5a26ad4c0438b55ccf552ecde9e4632546791bcd952a40e90314f12584c7ec51559e541b642520f6a77a9225127ecf5e5ec9e109f013f28fe25b8bc89e2ac09809a01bc1142444220f1844775364903b58ed94c11edaaa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41c1212d8a1cf22fb9ed6be3866f39a8671a5ffa4913dff7b3460bf5fa0d0e295798d370e3652de646e7ecb6aaafd963f93e193ae32a499098dee1c9f4f2b7ab07831913857fb6f937cb8d2dd15bebbb635902beb18f8f973314825d81f8b80f5fb57a202623ccf1f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10500b8927c45bf75e9b5c6d82cbee0f378286e4ae4a2963f90302f909a58cd9dbe1e790646060e7d5d58af3d9284d48ad7f825b3aee304574c097cf4ef685b693bef7027eea59772f640aba60395acfbcc8646deb0d3a2b30ee3eee0a0e9b88b62d7b35b6a3a649e14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2147bf64e6639404619c9becc044c016c3ce8170b74b695c462f9b431396503a46d171c1285ddd5098014e89410a86132de8abb11817c95a568f5c325c0baad6478efa577ec8dccb46e68a38210afa1d469dc828d36580ca1b37e10144d9575486a188eac8291be4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c3bd802fb2af204bc836c6183c9b1166a7518da737c57e7c36de0255f17a119197c331996206502eb03251606ac20d5d1f965e849e7e61bbb2cc383d9009b9270a344a1ed90d9d1994ad716f3aeab83afdb5a34ed63303bedc3757a7fd532df9ae248e7911868ee94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4d0ed88d96e235001b37880f49d6880903602060fdcade54a29848efb0869ae675c978966dc818e6534d90fd93cb332b30070d785e2bd9d37581482810c93641c50125f3ce39f8d0267bd1899f8225aa1666662a05ef2ab52ae61ef04ab53a80c557734fe60e51b91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da212e4e3cfdf983a68a53796b62114a8034a4616995ff1bad16e6ede78ebee4a3f1f8019d49f9415af83e013074b561d58c5c585093fa387891c161cc8e438209b6b23e17466ac5b591743a18b2efdb07ce5d5db4dc3370c94f60396e6584f34b31886d4eb3575421;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4345f8bf3a7db5301568e7017959d4180c7b75837da2ef879f932da6991732b677d0dc4486bc6874695d295d3cb1352ba76449773cd524f4e57d8a3508f591d21a938dc498c50b40d767b5cb503f6321f21e9c8b75625a373e4f054e1568189ff193292860e894a11b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102f36f50c5c58a60776a96a3370bfc3f99e0a11dff736280af288623e217a5fe7e6557a0b8631bc5aa5e3460411869b459108cf41d48f9081794872f6e21778645854b80f7c5481246ca781b900ac0580914bdfaa97820bce02bdfa09670fd307eb0518955be7c22c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b7cd78e3406a8083694153b19415661a9d715e60fc5fc29b31d728a288e906e851c0d2c598fc5bbce2a663b45c79cc76ed462e6b8c1b7d7cc152492f9df90e6b223a30c81b20f19f631a75fd4073e926f53341de26a1422258bf459169b493412d21a48948b4e9cb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa6596461f1afdb96c2208c454ec3c7613f3d9d92fbbe27459753dbe8143f4bdaef19c2fc47098bc2cbb2c9f916d231c97ff9035384f662855cce78937805556940d1e64716384ca8a054471ab343f469bfa1633fbed79b2c140562545fed3975baf8b13259fcef7f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc40bbb00f49e68526e11f3007fefb7227da2444bcbef2edccf91a2dc39b32c402a3c42618c538c605feb1af10cedcd0e19f31c53997ed8d5c50f3b96d5bb049ba134a979384770902668935bf5ad4ae2a8ac26b28ec98a6dafe6a0698b683c0491da436721508af270;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5510e632e281b6bed230053b8337cd580f67bbd949fd44eac1c504315864b1cb73f14e7b79264879617b9e999218673647d6967faf7b4485e1275bdea97f656f085f1c4b55c4de1da5ae17dacd942a71be3d19242d4356868d7820b329248c54bc99e3153626616f40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf739daf7112a8f522a35e2022fdd6d13782f9ec5f0acc6abde500fd59a754745032e5894e3cd9bc271dada544ceddae35202fb452689be8eabefb88713e458d2cd981efec3e817cdcdc0d5870b988374a42524fc150626aac85a48727dac575f511b4609283a1f4a92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff3a16a8bfd709ac9dfd58df491c94a18951618143e377189af4f69dd2a79735afefcceac0928f97b8ee6888449cfac68626307d57a12bcc26fb4be74b4c1b9112374a8ecc37a9083ad3fb00305614b5e3d30d985f7aeba53c623e297dc1aa5d81ddc4078435e15acb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122aebd353b0c3215b8e2e66ab178351d07365a11a0f2cd951e8173a22c6c6e9fbe70ef36484160dc208798f7ebbcd1c7d5d46fcdcc40084c2fddf4f8af2cda19ca3d058d0029548f92c022784b7d01e0e277ec3f6ca5df86ba4af1bc2a15b641ea73df10b001f05279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121870713c061f08acb8bb1d4de631b7b44479b53818ba0e52ec85dcafc30e57519c392b0e9d4113caf1e9f5b82321ef2b5f32c32a86e3b575b7a5deacb12dca41c35a4ab978c51d81dab5f34637cf280ce4cca126542c57560ce0f37ee39c25427bba4d2e1ab9431d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9bf071093e868f392ec68f00c5bd3e3d37883cefd2eaa4766890fe28a48b7ec03ad6b83be5ee9134b1b4659112fd28fcd876fbf5f9e90ebc0404d66727d2dde387e74f9995f13fda506eb7750c8bf81222de1b3c8a567d1668c447595da9e8f1081b965e66641a69e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72f87c104500cafeea16fc814fa7d23e970bc941ead8a31e468e16544068e4b6112705009b5c139ac6f1af39f593c3d89d9c77d7b9c778a122548ab28c3b7cc1d60d48f3f6fa890963acaca877beba103d74d2228e366f4389a50b7f5afbf02c3d8497650286ca3196;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159964e67ce6835176e01c8a1d28714d8856727657458f3fe9c778c91084a5024a52522434256aa0cdb428a81951ee4e92cbbb12e02b5b4d48f722aa864bb90d68ea3bbdc81f30b72f35e00d6584b2ce7212518b89c173f21f2cee98c66380d77202f0deadf6b0f0692;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe19a49489a64cbfe00a44d5cee0ee3dc6d392eb2a1b07d5e1759ff64482c9d76d8efefaa5563b236df12d48377f5e6b20ec02290529d0dc3bfea953eb2c401fdedc785018b2a69f02a9a44218b28cf31cbc51554a9b5b9239204d5218969c0fa8097c12e5407a3d9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h940351a2b7e4b294f70ce7cf2135f666f6f03a58224af8f536d33340ad077b199a159b4c218e6e032c16a189edc244cc835582cd260b855ddb9b5e4f8bf447c217351c9025196b219d537284935fecf1ffbd7606e7b78935757f687baa9b41566cf7137ea96532b138;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1321dfa71e06fa778ca20d53817d8ddfcdfff3d61ba9302bba2f45cc6e2a1c6b05eab266e6de594662ed58662d29c0f41d9e73165c3fa06f7f140a3d275b8632f098161fb9426f834afe2a19ee9b6ebeccdcc0b86eaeb3ecf6381430f591bbbbef272594e368f494c0f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef3f31571e76bb8d2be20c5aaf86766c7d6b2ea5f1aec96628b9bbc6f1929530430db607af8bec179704492f24afb27572e5e50871b5febe5df729af0765962b104300f8d9f7b444c98630c3eb43275ac7b8491db90535bffc13612131b6664af8efabf9845cbec6c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec9ba1f4f2b649222afc89898b14f862aa6e4e159024be9debfb8ba7792abd6b10f70930755f1f669b778ff5b8b0e449d1e101de83a30212cc4cd2b189afa1920c3c173541966b61fa3092360ea37ea74704b0e032d0a9594cf430cb4186dd510461fb7d46723bc4f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff87b6e01510d7e2ebb926a5f2a29e660434f8a8a3771c7ea2367cd73d0016ee468862ee92fd55efaf1be73599530f5ca842f73ed634237e858fcd114c8d0084a4e7c9d8c750cde4e32e48e82452575afeb2f8b66c25d5909633362310b16e661c55c9e5d23c6ef548;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h592055a24d28ac6b7238d68a169ffae8223bd718b785be805fa596c83d2804c22d79a1cf2b471f669ebf0dbd2f9d5a985194e4fcf076997b76fddfe7ef275f88856771b985968fa8579e7c651c20db9db112e1de4aaf371bf50afa36ed23c7508551e672618f68a9af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121f4169402041f3407b06df283a42f7cec52eac27a33601051a95be77d60c5e30a1ee3cae48727b4b270f19d7c9754665fb7e270fed0127bb6eca651715fefcd1ae470d8f8961160f54bc4aa4ea378487a8fad423117a624497a5445f4634616818563a0837ebf9ff4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d722a22a2abe0448b8732b9c77a013212ed77916757a754872cdb7ed4808e86246aab7ae7334175a7f446df1e05bedf77a4972cbc5ad721702bc66253d8a0ea21ac36a406603473db21c9c55f0b191717529ec4219543d6729589379c44fbe45cdd3018487d60463d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1377d62b8dfdcb7a3a2c206d7e64e4dd1ddd09f1584db0f6fcfe566ab0a76f5260396ec067041e5d20296b89c70c6540a0c8af1f557a9707e135a272d3e81b03bd1d658fa374aa597005f247b5eddcfb58973e4a6b92b9fc1a3d071aaa78c37bec56c92cd55b41ac903;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0ae30f4ebb058bb9462357d3639a32c77b84de54b3849e3aa966a26312879729504981ea216a2a41abf50c49cbd3c33ccb5ffdd6f8a13b49bd7dfe9d25b3c8bd7315091f2e5de5c0a70355a9e209ada25241a296e70682b8f48563a256c000da94b825f6554b03ceb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5e53a5428cf2299f6ce3361e9f7e991dcb9c80cf29335abee360f411ee5e41101b5c9b6cfefbc9cabc4b96ffcc1fb4952fb72cea62a84a7eaf8a8e0097288f9fc79c5cb274efb7b20172e2864397fe37535e907eb3a5ba19a596992626f6d21c36d8350ead0936ec7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2c799e87369f0b8924cf47c64405b386582366c090c66519a7fa34f222d61af1d5ba463711ab8c667a43a4aa0587abef1640fe565fc4a5760be6108e50789337d806267d7b1b8e556cee806a5883d525f2e405adb052ad57a524c6cce092f383fd170376adc14ea4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1374e894af97a04e6ac6d821f05c9232c15d10589e3cad71f8d4d73a83afdb5269b2dadbe71946657d591b39c3eb774e81cad6b3cd4e5279004549c754fdf2b23b7f695ac0b6d2f12bf69048a9befc43f20523b17a0e2ea6df14e62009bc16ee94bf74c12fc923d0f05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78bb43177952430835c26de9034a342e6cb72492b69d15cfbfc52a2d8b9bf9ef925c370d502ce7eeead21ced28f1b861a8aeee0b7caf76dd4087043b4c3760bb143fc99d22fe77b0b14422a27c8c50eff9db3205dd16ab45f7d706bd03a107f88a1df6b7322df515cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed7de5bd7bb30d290c94d95748b1a3e9fbed88733348c9cff0ad6018b45392a5001be03754c7d32b544481b3bdb89678fb993ad62ef1493162f16f4a323442739a81958f59bfe53c849c8ca8f7ddb0444ac478c91448f25fea2c10a7aecd53e37772d298db132395cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90839420dfaca68c940077a051ac6276cd825138a8a083202151fdbed51a8d946a6f359e2a7657ca2b00e3453a41536dc9c802bd480a36a26a7e9c268b7f20bc8eaa86ad9a2ce97107e6b04fd65b3f602522318f0e6a26ef60c32e7f5c932fd19452c9fb9277393efc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17650125b1e223eea5700423dff5b8817458a3cd247a22e1f43b93b27871dc4e843de3ff7d1062cf6ce806c09fb8e927e12aba167bf93fdfcc0e2f38c3bba5a52a7f6b9f9492f4fb5afb72e524d336f87e3bfca2b87473f513c582e89e8bd26964deba60e6e7be237b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ebd3e54b4565ebf3ba728b330cb38bb98b61d425cfb41840083ccf79957f2cd4da214983884123abbb1fa1bef77d1ace6d8548536b3bb8a2a3a0b8aa7c72ecb4486e521128e645a72a4f03591b06ddf53cd2bed3dc415a4b8e143505ec7015b2b0cfa987d0352f8b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ca4be30ba8641ccc668c171bae48cc4f0a8c8aed7e674efd2c343aaa80de2475f2d201b60667e8644eed414427bc2f575707a84d83942dec48bfc94af17daa724aaf8ef707586f5332049cbeb3ef3b3fe129ddfc4e48daa0a0b4f82490b273a2cad4cc28b82140dc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18bbd0a67446ddd69ab2d3cffbd409f1d06a35f8a0c354fa036f43e585d29141f1eb3e1d9e2f12b1a81dc064defef354c366a885fcd804d427d7ae1249e6acc855fb4249f1eb0fccc0ff4ca9f2a5130add15962b95378e4e5b31cd77230458db36d29b740c141a6ab10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133ba23199f630bffa2d3c28c856a771c88d717a7a546673b164650d3902fbea23e7350f506d2f3eca723c3740952f1ce5ff6f1f0728d22d267cd71c9868f094e696f9427151c78ece8c1fd323cfd7c65c411c79f87d3387bdd839bad490ca971c21491847e0325eba3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h317dde612671177bfef17b8fe958f512650de4b3a9567d9daeb3737dece73411b0d7c3a5c3ad06dfea569871953431936781fd671a62982de76166f86433e06dc23626b18da09db28e403b1b4d83d9afd46b2eb309e7f7780acf086f2eee6afcbbb3eeb1ef6fe33f07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd70fc7fa735e47102ffcbc47561062f69f1f8c4244f15d0ea4d27dadab148391ca5f01a7f9df3e1bb160c9f698ec1277ecc7d322523ac12fbf3081602b2f632a91340f74dfe98233b89fc41253f5767dfc237f865e7e4f713ba825c28daaea6ebc2d122792fedc81a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9cff9028d8ddfdce97ca01e8a37f1404cdadf88f7c798528b7704f792335e676345adca941034be3d23d88e89e87bba160cb073b015d47fb648031c0ef267e2990dcc59d6d30e4dd61266385ff4ac04a6af7f52551a9179dda8f9035f77a90f981604f3dd60affad6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1366ab755a231cfded686ab36c266b6d21d576c7308ceab8f84f913296d2deafec70bf7d411bd402aefafc9970e1b28554214da7dc6f8dd7ab1c03e3a7568a785b61b86d3826de767274381e71838d58df4e494f30687daebd14d741de3557d7458ef9dd178eb6c0452;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h386f4d4432fdd19d37a81f19945d32e3b5adf71d64717edd90b1ce9ee6bb1f58c6e42898bb98c2aabd51d6fb310bd81fc20d7fb2fb5a842f5d7b9003efec9aa1a9bd997ef4f71ef47ee63fe9280979d002cc6849e8cf957c5a756fcc523388c83fe5385f32a610754;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f68735d9a692ee202273fb007025a4db27f8725af415236a0de96195db77ec38428bad6f8087beb8381b3a3d0a55cc2b70e237581fe6555395b995ccdd1a79a62da035b4563abad3494cfdaf74450f7ef5df500bf6ff9c3467f0a002c602208200c597b03d161e143;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd36e8ad0227ace5d6842dbe8b384df5295c079c7ab49e958c039649af969de1a9ccb00df9248bc6ccdc5cc8aa592b287edc9dab5b17305dae34c7b8168fe38350b53d05ac8dadd6501c0c069f765d832de4e6171ff7d1f2959156e765ad8b0b7f67d6d2696ee215c43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9e8a8aeb8a42e3a0700babc7fb80a76e129e35f0ff8552453b0eb465f0cff8ffa634b583c3d30e1321eb00a65ed9655c1a820dbf4510bda901f80d486e80839c4dc6b37301e96ed4abcd7009e30081f5742b187d23599779c6c8f007a75cac1c27bf5639162079688;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd4b59ed59e1a535cae94ad1ecca4adcf94e9c95304b4da632af780533d9214fd3da66e72ac1ebdc3699c53c24a9d07c29cef0a34b53a06cdede41189fb641980e130e9c4793f78b12a219de5e3c8e2c010edbcacfe7e1ea97cfddb237ab4800a1e2ddd038f300cca7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8dab632c11f048ca0c75dd9b3273f0450992ff6ec9916fe1069558f517e60bb1071f68dc5807773c22e3b67a4f513a8282fa8683f130ea03a79d44ef461f08d825f070e04073f701a62479e236a39eb1393c5dcc78bfdccc0f0ac095044c24e473445a6328df5c67d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4973b45b19160e47c021dad7762370a1fe8a6b27a3aee2f47623766ae897ba3dea786139318bc766a093e352ab2f3116e385547efe921a2d1992cbd9f1024e1f226fb33101b85654e165da11bda6950b844b18b4762c91a59db4d5eddbeb908a8d4b87264a0033d24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1002df678e98284515bebed0c4cecca6dc82f69fd33116a84960b368124f9037513a32d623bfae5cc73c79ee9340e88226ab7597d1454c2a70dba773e6635597600b13dda96dc2beec6d9216de17420b7de17f7eb778ce97c82254e8cd87ee87d5f5feea1a6c698b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b03792f28e0c98aab16e5a7031817e8722dba3979eee612ed278b07d4a284759ffb9fe622d0d354bf5c6eb713c744952109d4839b35c6d949c920360a296fd76acb8fc967119abdd15a2e7d16d1fb05ea221feea3da07132cfbd8de5164a0da3c13f63b73372be61b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb603a4289dbfe153bceecb506b9186e95fc81ce610069095f27221082bdae4345aa4a0a64acacfdfc8fe1719bde83c22d55e971b1c8bcc66d01928c758fc6dfbf3be062aa49c4fa27f7988fcd0b10c01d495659a77b8d50f6d34474dd2afebbe5f571d3e7c81b999ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0980d867f39501c629b70c02f36a1172565142b64b66e81b4242bd3d647203045f6dd57b9795ad15bdc20a6e27843ac5fb0d53b934fe6670df32d74dc52c6ca12a8e2768653be640a5e1adf651dc4137dc0a8b105bf4c33dc527551255f2ef78bd77c40457dfa251;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h390e1b66b092d505570fff785804bfd5e3334000b5b4683978e85c387416f3e8205823e314df6fd34c450042f06287d5ec475616b3d001fcab6033e5698a9c2dc4f88e40b6b5aedbd27d126f0636049fd940156f3a5968b82a7bb49e355cc6fc1183f4e785b09fb977;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb35dd3658068abd89d2403c0c1337b8d85886299b6c16fb32c95a3a3803dd83886bfab29c4b7c5a646b4f0879afdda43d95b5de9b2fdf31e5fe28a2327587fa1698b7737a1ba8d233cfb2d0c625c45ac02b23871faf0b5eb0edbce26acc8cd2e5b5a3fe2e1dd7fa86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c53fa9d6024df3aa7ca7932a6d5b85b80aa72590b224fe2ac2fce8b0c2fb87c4bbce24a76cd7829e4a7a7d31324b58b2132bf74cfd59ddb12e5ae73ac7c58d48e7f9aa5c59a5baed781c2cde81a1d53b6ea99cf2f21948b1670bdf9fae24a324ab1dd33949460dfbd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b08503ccc952c07ed4730d4f0cd24c3068ba82f0c2ac2d70a8cdc8292f95513934feeebc8edd24705092c45cc9f45b9250e5a8e523cfed0c1bb4d0956ec148c3da4e6f633382b1d2a8ece5c7a10d6658ba8b30652920a2dd04bdc505fbb2b9d3e0e2015ec47135cb6c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d9f5821b6370987283b0a0e974fed6209f7ad3e14a64ce3d64d486fb909b17e51c3b097f3bd1c739137058f998fe0bcb0199b21ac50d1480dc30243853c0058ccded5c0b3d9f3cb4269669ed74457479d4ec7a8260aefdd8f3cd218dba1c016f0d27506c04eb7e56e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99e39b4737ea5b880d73021b3720520379d2c5a0fb631014b1d190944ecec4bbe5541dc57bcc27a8f88b2f98cf927d721f0a921add3b5346a61d24612e5ff1678450357330c2cb6a240b171c5593cb287f85d99e199720cba67830bbb70779a49d2e8c2023b805a7e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he05d4e0b3d0b22bdb64ee789003fcd84a9f453bf0ad9b63ae9d12232ef5ef6e27c4aa5314b48077751b6a9baed4e1cc03c93cf12ec2589e255c79d0ead4230fb0c24f5ccb8d53b0f787d4a5a1ee5386f137024bc9b54bd820e83a3ea9d80827a6a480cbb27912401c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5bef512a6e868fd22601a36def491c8ac70099f550d33287930ce95b908d2214deab5801f9e6f5a0fdc0a82455061948d0f319a1ffbc62a97e1de0676cc3f0d0898bdcb171800543fb30d341489cefdd5b7b40c0c95f945035dba0b449b07e4dac81c839e1b556a94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf166cebb4afa8f126d5c307636ce5a1f9aa4974bf942c8b14bd8ba5eb877e2a379bfbf63913df532e4170b306546797d9a443d285fab9efe830755f681dd6f0a98f05691147a40f4d59612e77fdf5f05f151dd075d831c6d07519a458b6d047fc1c8648fc5ea4c339e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc9a1d1625ab9dfecb9da4f034279a91112bc81ea4d5191bb21a9558f233b9dd39e6ede8e624ba9ad74d921f63b026881e0c9b53319d67514f9b558f0bf9786a9c9b4a466538478a7e92a9e0f7f3d0d04529e3dc22b8cbd6b2b0413c2e257ea7b101f75e5f14abdc3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebe06d36198cd7c9f561c5580b20a85c50f7a5b0580803633d34f07bdf27f31017122ddbc1e8a61179d70fb085932f60f2f74baa0bd6476c11cb3f5bff1992554005fd18bd76681923dc73bdf9e9db5a8adb82cd3fbc7ad90b1956dd5c948a9848bd33cca106f65c9a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175ef66747ad094402138404d7cbc7ee3c0ceadc77db1fcf31b48f49206a6baab42203bfaa8bc9f0a25903b05dd213e322f0fd1b1e56255b17a2d9415a12ba44556a6d42dbb33297b23f0db548c53c00741f2fcb22a76abe2b514e6249030e78d7967c350bb3630bf07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc20792adbf060a748c066d79c4ce5d9be46ab744b9792a6cf8a9a7c81584a9ce7a5652144a90018c01eac4f197d8b76015070cc0529bacac798b97a9971658857b89c4ea11b18b287e94fe2b7d7ed0a3a9a61777f6736d8929c7826695cb3e3cb757c90723aad11cdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h37391827fd85221777cc226ff7e9e62ac2aa5f809e8bce7f528f1e2e3a2f25dc218d30d2903cc540fc3560a7c2f628ab5235f8822c18124e3d426539948e54e819561a0c9b348faaeba380a6ae487902a18a3c79fd37e224583ecc3d694f6a52bf916ec328e27d859a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dcc4605f22b898de03c4262609499656dddb1fb9d63cacfe792565ce4cfa70256069f50e14e40f5e01eb579100d44686a62d30f9d60b6004b8b0f3fa2075175645b21c8059ab4f10a730a900ac7ec0433d4c3dda98d2b8610afedbaa3732b8def0b6a96c6f82718459;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118e4cd3f0d1eee804df91b4a1416364bc9004c1427ba50e58e1314fa3726e1a75bb4e9f623ab1a6c2d2eaca01db757806d5ce3b9085151fa529499b875b7894ebdd7ae7e68cc51418a0cf4d61122e48a4906c29db0f18142e7de39802726b854537c4aebd5495ee138;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166634f33e62f5df0e1276b4a129a292b200dd656a4d5f8879c9847012db254da7066ca880a114cef4e500743d98084b33d7e62de306ac2d49985c6192c5e7412de3fe3e575c2664aab0730dd2400dce9497b0cdeb7523c455ff117019b658c2c79f8c93e5abfd03390;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183b8846f32566f8172544927656ee3e4be1eb0d0e8dded9a6d8bbe2524f10f97d820c9c88ef8c783a2028e727ac904d7f47c1fcd1b8bf7f05564b2fe3029526c913806fd772c6a174180d81bd63e5eeb3381561aaae3a513195c7017e7ea1e76c2943390477c2a5797;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2fd89a090ce60d897a894f879391f0c36254cd95d8fdbb50e2c93fbc2c02397cfeb5e3a635e222dff77194139fde4820d16540b09dbe5f78262c6bd19a268e01c8314371eaf6d7ff60c3d8bdeed9acfc1e5339c00761a3a2dbd93e63342d877153ae7047a13d7f1c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac952ac8c6f915656086f528310c6cee7d52b707388f59de225d74d81716ab4ddd0963579e542357df99674381eea41691d1fc399be4d2098468f1b56e05eb8a18a82da8f88e6492a0422a3f4b8a9a89e32b0bbed6be02d040626260a5c97c58c41ece55c5a2c5e55c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6a037987d15bd8b4a0424ae02aec0eb371d5efb18ca1eb5f62d6a80b1c837e06674bf0a7b6faecbdc5275082d2fa2f0ccf766e2ca1205ba2ab2275f3823d2821b1db34db05655417955e92998dbc7f5cb92cce35b5ba0cd76091ee03995d6d8bfbc2a73431e7656c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ccdbeb203cd743f2a8911abe22ab94746117ad8dfa6a3b290a7502127830973c47ba8dc04405f9f975842c0fb7b3327888dfd6007e48a543ec8f028b3e3b0f3ab025b9792abaf84a4ea6c1344a675c9aaaf55f7b00287be2c59378816e4f0a963a38f301b89ffe666;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1970d5250459d1b625b7a3e93a7e7ba3578d31aa97a74d1dc32d26cb9f6bd44e07dfe875aa7e5ec7d07e9883a101554105d89be763644e0bb28c3e4f9656a3c33a609c1417c1ce1faa721751de01c0b463e2e6907c283104e8957ce3a71c0c7d93cc9a0c8b5c6a31028;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16738de0eda076cb76dc02c0d9ec0ed32adf8925dbcc5adc7582c72f97dc4a41ebc7916777fea64ae19d244e02afe694a1d48f57400b375740f11a94638e64cba41ba51123a1c96d616f0781a350147a9b759ccb08198d84c297004e56d4da5087dbe8d07fd991daaae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82b2cf06d74dc72749bbca7f0e7469dc0f31bc928cd7cb990d03bbd513c8d44110daac447133854bdabfc3c3b2a04b2ee4b663a72cb8537ee41f6b43097aafe343e23d47622f19791c80c744222aaf8bef2c907d37d64c00920c6b9f63f42ccb69e1e4b46560cf1533;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a62ccfe2ca569a04cd1ecce295542107890e635b09ba41931d33f1818a9fb10036d8097e60672170a1015a3475b9b0519591e08faba1266138b0207ffae683882d767a80cea96abb24f0eeb7b42671be110b684f5e62814cc2cb25c5b0756dad185d95edcb6e73353;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8ad83b9b03e6ee635e346d9ab753c6669134578c666a087419cae19ab7da3b76b9fa977f3f740a12d35169c3eaa00d1773040dc0b84721dc78a6d5aef31c2abe5b6189d10d923842bb5832fc6bc61cb431c6fb65a63ea7fec99ecc06bc64c900d90cb5811cf14365a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac729d881c4a152252fa0e493dfe3d13b2d3be9375720026bb4fe4b82cdfebcc241e8423bf87d72de9d95b75934b5e01bba809843fe9b59dc3b04b3ec5033c4e76bc2bd2ee20e616cdb955c354ab727014431a61549152e6ccc8deb8f04c6f98f505a128d189d275c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had8fc847a2cb2228f811bb3ab476f1de1f2bea156b5754643660816f715e447c9f381f9dd107bbec0cce40a83248818d7f068e81a2b013803ecf900a772e5e8d7cfb923d0f5d9e7c013cee341aefc9113b4c68d71a7e779ead97fc9b53a77c67637e75295064db3fa7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd271c2a126f401c0d655ae8faf345c0925a1ac788ac75563b1685bd784d773f6d16b6e29f85c1cf84a91ffd2214d61b2aca26449f415cf6bff4155bef79bd8ec0b2e13d73f91a16d286b09053eb945848e21a8051d923f2e8753d07fe3ca9241f61962a9529deb5bdc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h573c87556a7db0bbc3e9e8ac29b1033a042b4981b6d0ab908c3dc7f83bf115a85431198065c16319c1edf57748540d26472c01e5aec99c233ca06da28dd19322f4eb2884e122263b5310e9a13211be30b5b21bb8f7b06d4bc253eb41fe34840ddf949b805259deca50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abcbe29cec75b950027d8f6140f2c305ee015a1131ef171fbcaf5fb5b383fe06cdb3a876118997446b5fdafa7687995bb2e8c5b7f84d2eb7f8119989ea60a7f838a4bf9f190e3ce37e7d923f29ca623b3df7b765e17f2af2a1d4b1629d529b7785d8b8574133ffac78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cba61c51f9a1ddec1980327998cb840b198b0a88a02b3abe9993a25a6beffa2c04f874c5854d6f086662e4a76ca21b4bf01dbfdfb82fac8a2698b8fb00c3b43aa226d3c75a4789946024c088003dc3030df7d601ab04eb88726eccc845ca42597ada7d5e951c6ef704;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6e3dea6e051772407d0b34b772b0dd4800b550cfcdafd6097ac24956da8cbfdb3ded8a590929ea83d621857aa67a6ea2a969729dc9c20961fd6c5b65df477c8e47c0055c3383ac32ac8b0ac322d7292571e77219aa1fc5d50649dcd160415212ce27a382c9651c6cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bccb7ab31fe79d782f58b7c3e0dcb9383f36bd6abda4e3248c53c7296fc1f9dcc1e747161541c217baa3e5a2ba967794518870e8464321c1ca3d8af0e0c543a4f8144b89506c6c731fb36ede2edc6673438fadce88fbb79a8e4311978886eb5dcf5e7ba2e3a8a029e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4edc6079663b0af59d0854509a58db228744c14c090c371ebbefa134466d1454b5e7bb2ceec4e6c4f6256b1fc1588668d2d404535f3c6809562ed3efe30ac54fe396e19e40db59292ba970ea52e35bebc8b2c53ace70ca497299969bf87ca9f9eb844dfb3a89fbb12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cecab2e7f114644e2306d6cd9b2ba751c94863c0b898382ccb50e02ce2093f3f14bb3ccac5be5f1df04062bb1f78a8d3110ded471e69919ea16daef97b04ffc4b7eeb00659f22be8fefbc73eb76bf90bd75814c082a22272aeca1f20e472bca6884434b70a4b1e8d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28338dbc9546a06d29d1321389a83b5612541c1c30750df0331fc9c54ff3ab897d7289f08cd2af01a3fa690424013f3d1ccc42e4a9ef1349bc849312be45b4cc32bc4224ee4dd3ee83d1e55cdbaac07285ba2d56a7093cfd1ae14e98821657c121b6103eb7910de6da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea09d3987627ed707650d6db7a097d5d0c9559105991f81e5125ced5f4956ff7553323e1813f16c6e91dafc2ee2813d35f8f63e90896868e68a7a071757830f36d7945cddfa8e5a1b88200f64351748e417e0faca5a064392f5667c865561174b923c743736c8eef2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59ccd343e1629eaf80b7bc7efc219bba57f582c8331ba5110cfd35e5e69cd43a2585f99d9e7bcebd0bbfcfa08290899f0dac4a42d91a45f8762bc76e5c52905fd0a80311f75051185775c4cde550a9689ea5a6d7a89e49fafb57c366a659fe47dead4c878e79a52d75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b7d2444cdcb612ad4d8f01400471aa0cd33fdd9a52ca63b423f6219be72b1c938e765c89060b9f3eeda777d4a8b61ae6ddb6790d0f24f67fe5a15fc8c22f5e702e0784baf75c094a2222241837489cdce4a254d20a1aa4fb2f971becc05d0a2fd37d5e42efb9c74e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fdcc542934ffc789f3b572b7d659c75c8bfb98b1ef1232fcc9b1292d6c517168d8e48b8d60839a77ea45d7001fed69b3c2e6dac8833b033541aa8970571cfc8254e5fd09a816671e167ca7556c72aa42bc9c9f8dba73d5cf1d39d610e5a62860793f6a140e3d856818;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f95934f5a8a842983ce25a6bbc51a7cc993c1488a85219184ab0ecd5766ae1674150c455e33d43aea1e2fb010fd23a2460ceed2d9c6811e59fb1929c1031de780965000d33eafacf31517cdbe8766c406393842c368fad4950c2fc357e8cde98e47ad36c9db8adda80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88de07a1dca644ea928abb8e5ec5f1850d2eed7be22d75a82e845e7a839c87a54c39adfbef4c1307db15a1ba66af9e454876391e432d1659582d3cdb1820214c51ddc39eabee65dc1d85edd2df004f93db650fc88bfa6ca1ea2db80a0bd89791a0e1d365aed0a2c904;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16dc5cefdc26323135ebd773f2182feafe50b338594f0fba3279145cc47f29972440622b77cb324d05b59117210837aaaf75344e5eb97b837b0cff1c5d571be2615eb4cfcb6293130e34f57b2f08927435d2a880a00f3b1602656c0b3b23e13ea76bd9dd11caba361d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eef553675505fd0ee438546a18f64e6f2013cbdacb1dc446fd239e33aa02c302617fc996c4a34aceea5fa479ee2655d1106a3c1296ddd78a2dfdf9681bc730133d97337e64623f9e387d673b68169c39bfae8c6adc1c50c0df4c28dbf3266684ecf052428892ebc8b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0829b86145d6347aafe0108fbadbb5d69beb4bca07a64f616751b7816481f14489916e24af50046c4fc27f0e8a66a5d423cef5b84e52d08c853689706914554683a4ef928e61cbea2ba1c2a73baae6052a7e71e0509a507afb72160cfe7301ec12ef6fed5d02b28bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7838696e8f874e1b7e4eefe30b6869bb15dc86291af6b90e18aa59a236b67f95b9262e64e44bd43996b6fb39d47c38fd2d5ee4b186ada45c1c152363cf6d5be2dd4fdac9c0abbb33b59acb88d4dbbb9e4b16d2dbe5b926649e9ea4a7a2679d92b6e3d5af006c4c741;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd6fd1b3f0e9b073f185ff5b47dd4c16e817dffcdad3383a6b7d80f405864cb12a50ee496ed53ca61e926041333433137dd0a894625822ed59a17ecf4f0cc0ac562d6e9ffb4aa5091f4dd91e2367c8a48372ec87551dcfcf54e95e1eb601f247c11a9bacae982ffb4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185fbf61309620f5e0641ae541d20f4607ff1b4a72d7e4058f23c564207f85ce72084899191f2f26589b57d9cea175afa8a12c13c0bff8cdbba5ecd9b9b3b743fe630aa41f2ab63d68dfe8bafb0dd11c56093d494d0f183cff7273e66e59c882ca77bb8c631d32a1e3d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13208951ce6e955046f7fc4d1da249d2350ad662b0e5bbcf2af0a47996d65b0d8d0970eb6119c6c6a57e093e4639da7d64f9a217e24463179965356080a4faeab84182b2f36f87aa4c521fc7afd7e6c992e33d3fc848739fcaa51fdf67c85e4a45759191f54bcc17098;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1adbdde127280a59fc32c7456a0ed3515a0a9cf9a3cd59fba282450ccba71c5e74393374b98ac09527d4b9e5a53c926c36e9b43ce31430c06ac86f52601b2410fc1a804f6049dbbdcd189f9bdb7cb9f9c9d8a2fd3d02cea9236ce353a91440fdc2b185adb81de575750;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h859c598d3b32f57c8d7029edcd524144e60f0274096a286c961dab48b5096356fc7b1b732f3e9f70f7127dbf22cb9f78425b9e1460383e56f19a6c186a16dc4e84693b248e126250a54fbfc26eae8dcb188af46479b866a78cb69aa73f0b95a4c6d3a3f7ff4dbd0dbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c85993442a605f7426af6728839032f11b16380e0cecf5354602baad4056f0ee60735b8a737775626b5b60e5cdfa781c4abeca9dc4a3389761f05ad1bf5428440d22e0c5d4107e038a5671ecc22dbcfbc178d507502f29c9b8f10c785e839486831a5284e5ab7ad4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b630ea99226b0422da80cd5b5e70a5b98c97b7bba2c05bdcc17692c327428354104f120a39c436f7dfa7802ae5164eaf5ab3c7cb51e97da43044604cb570e598a67ec8ddd1909b54d7a05a76f134ef274382313807b120296b3fea21027ccec90910619ee6fdb69e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d51bcaa252fb8ab0e42196da123f85ba6db201b4bbc662eee018ae6f7ec8994de718f6bd45208b0111367722d966c33c90794a9a4f74cca5cc3036aeed084ea9d8f0f73c95ca7d52f55ea65a5c50af538eea0abbc38ce54c5722a4f381ad65e5c920b837dc77c147e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fb67cfc077e5007eab090380881501a991eaffd10aa8be1bc1689304bef7e542eef8a1fdf4635f9448dfff45ed1059c4c3ff2289eb74685c1205d942fd22d3387b5587f3a6c4dcc537ba2cdeb075ac86f4c7fc05d88ec53ad202a10904b3f5eb01b519b21e5750f54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95fd0c431c80ced9400d46807756b61e55a772a069f7c4154f3f09dd352f7e7b11aa3ca0bdc79620a3268e790cab42de5dd225f9e20061b54cceb83be174a35d6ebac2a4ef222f93b60b9621107b8b9e8790c7fc56d164e7018d228f37bd2040db80b9e773da347638;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2450a117071a94014b502a02dc250a595d010b7811ffcb78327d4b5ae9614fbbe26f9b3280b8ac854b17addadd76ff5e80752d2b040580af0e9a15ef8de3aa6a659650686e6ead06c65bc0a3b58df5bc789fc368bddd77a56d367f5ec9c2f0734b217571a6516ef24b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123c8e1032d7a24b4f2d277944651ab372adad760a9a484bf369f279b08d383d04383832cf027a83292b81905d2177490734bb311c84bc7e4a2e0495ed34aef3fd2c2d2291734b5c022be502897df2f156aa5f09761e1f272b7d2330b5508764948fc6280f669d302fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1feef3ac221bd963b85a5bd9d6f686d47c98a843a68c9962e2c00366dd81a048c1b1d93b9e77ada3525daa5f5b0a9be084237491da1c66bef4b52de23023d72cf41d67e2a6017fa59584c21b612c3f3b8e5853c25ad455149828983f299e014bd669c3fb934e79e1ffd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d6f07800a64f2caaee871bb912a2957dd7a908ebf4f6e1ff43c8a86aa076371d0aa0767faa94819743f4aaf7e46ae57025a28822c19c9570c92d2bf8363ae75130ab864250ace3c6118427853333f40717494ad742bd201a477e434a4baa684ad78ae0480c131e8a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148055ea23cb063b128f6153714d1f7c1d148797971227f47f8f61958ed30bd8718b64f7e6918d028bc1fedefad6e299311509d1a568c7450f0ef6cc47e320310c94c6121137df9279cd46a1ad746a2778c10f472274a8da8b6c5f05cd1fadc0b633ec889a3d08d3116;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h426f9988f4396ac96062ed4b504abce948a2995f19ef13e9bd9c47dfd42d8db17a8820888d9c4334d0b73d7a9f01038ed7f25e87e6a0cbf78ad9858c14c1060e36b87ceca1b1f414d2e0c1fe7d32a5864dd22ae605eeb21af88d2ed8094479c9a6166ba8df03434bc4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hedaeb2c1b0a8c77c8ca5b1eca67014eb03ff174a2c0248ce3a090d24d308868985edcc34e88028161c63598a6527874b488fe0633776c2f85b344944626fc650f4bf4bfb0d1ddc0299d11da50328020072122e197b47e917dc5ea2945d6d51257a852462e795dff5d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f141f5cba4f312149e17fe119ec40212b93b8302123cadbcf2cd29747da1dc0b996ffaf8f380d9701857d43c7c9fcbcdb94aa8f923f6da8bd923b15ed05b19d6b11200ca4569e640542161c51cf17d140e83cd5755986f11294570e34c241c3592aadeeb7d024b676;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f08d50ad3e3bfc560d7818d954f2bad12804ea505a9bc4f3f33aab492449495d9817dcca1f9d685b90cb6f4eb576b026eb194822f66638382aa92ca6297d0f1277dc1bc8a733528fb063a632f88943337200ccfb0e2d296f5362c5b9bf4f075ff1f7e21c7dd27ee6ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee289e0280c2a7883b9838fb7a6bcab579a88f6b0c1844c26f70903e356b7a31c64ae149f675f3bbac528cb44a730e173c2afb710ada560bab903f19440bba1b289705a0b689a5b5bc4f2e78072785cc8d1910e9d35c167ec3135baf41c475cdbbf196e4a531c72289;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h747e55cb2341114ce00e5d330645a553d5f2ff73de2ef80b93063e8d47a30be8ca87366a9303b2a7bae01f27c7e152587244d0086754bc5f33ed7acb09775ee2cc2e0bc7b24fca12997fb2fb6841e0972e14dfdf139109be762b55cac7f28be1249c89e5fb7048bd62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab088ab27ea05470622de0398b37ffa7cb1ea6b779ca7e503fbb5089a2923171dc603756d9d1bf52014db166a7446f7f3e25513de64637b8203673dd787b34c172c463435b0e54a74701d6fbbc528142a3b2f9d884b75655340d3e3b0d14de5931d04402f8b89d4abb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4649aa143f11e9551acea2ebfb75e8dbf86104b4a8588bb4d0c4a2eadcdb782339748e5d81575f21764bf0491f3695a8718f6168dacb6f9479c07f2918e3f571bb582a1ab47c7affc38c473f2bb811e48ca07699552fd2af9e6c58b323e2d411e1912a907c60edc43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a088d82da2b96cc03c38e58337532f26877559f01270ff9001e98cd33288cb9b07aeff8b44f5aeb6b77c46647bfdf61338902aff437a2803758b4af1a1cb628a3d5d6a60e60d0ab961839ed9905a635e1cc3cbef29fad9cb8c9e1ce9210aac4efcf624db1abd9d19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98fb103f02e43a6db557db4ca2ab49ebeb234cb75c7202e94cee8c36bed87938db665d41049dd3a0fa47cc3e3e9b691e1de6cec26a4b79bd348978f54e5bdccf389b19922f5c9e0d0cbc0246b950b063e08c658ca856f58879d320a8000395b3ebd50b9f3ea770c09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22bcdbf9933c160d4d28603ebc5c3dc6d21c63ea65145b8986e44a3217c7240326ba3bda75e9bf7bb70a66f52a9dd1d600ad72e21d971e4ca448c6996f12a8b616b88cd182dbb5939aeba629a8b56adeceb03040c54551b2df2f629a848f72abc4bc3d97eab3e41b81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7545ba935d6c3ca0045d9902ff97893534d1c7d7bcbe33a820ac0ebf771f11f9f066e3f85ff2cd8002c286e2597b03a546103495e2e875abb1091ac1714115eeb95e647b4af6609102d03b7e49d39d68e706ac273eee720dd5968eb399be3b758607f235d3eac089f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4d46629d9b75fbb9ff396340f1628b1d380c71ab4819f2ff09b71a6c80f9cc3b7673db6c5f381fdb95fc09e126172250cc1d44194c7fa3c9fe2ddbf6e2a0d042d7d74505a1f4ec96b99c9602e11178a428bbfd3287eb805a9fa26a8929e02d4bc65be8c797c17d3d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126f17d76d796b4fb566a8b0c514c5e374485192d2fe456787d2ef707117cf6d9e3b73ccf9a0ba5e8766a18e654760b3d0e7e9d939a99ecddb6e4879e1f17833006d6998d4815153492fe0803038b8fdb648abece792710f1c8ea38d491a3a9bd2133984f58fe1c8cbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1f9f8d129f3404b9f172eae5fe51f0afce9f0529f66db203555c1400b721ddf72402039ebdd8165801a98e670aa5b1fd218f2f9c843512907c7e6f8ec9c91f58276bdb5e8e7a4c7e296c97bcd67aef07738b9d077851a5765bedfeaf526f8773eb84b002ccc3dd0b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c53c83c6333954ab878fdeadcc094675ed03a78efb1bf4c8e671df1b309426558fb5d68a06869a810aa720aaaacd27accfd80253846e8342b81ac4586c4c4064d57da98e366c71379df9fe9778659896765909f5d26549bc2c594016bbe1bb39c07682c1f8d73c5a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac9b912c25fd0f1c7aa5dd4c2a245e7ce1cb729580f78f33a1475e0a040fd3e1408a28ff01dbba68e443f3269fa28dc5ecd1a8265154ab9bcb85f95b06f7ffe45a651917af5ccc68f8b9f68fe1ff7d2a1fb243d9fe25c02aa2c68f27150a94cf21a4e4a12927e6b187;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2a61e64896b2453da9ab2953dab6ff7af6799224f6244010c1b155ed81cdf98a359681ee01c50dc4f5f60c9dc2cc7d527dc0185c0985efb3ad0f2f8b4db8fef85025af4b7b8efb70b69f398870a67353960a24e85bed478e3804157557ae42eb702d2c0365c713db7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfccb71df7c4484b8da67a2ada8de42a9197d5fca8b0c78b2b1e5f265ae65cff598d4b7510f9b949c39e66495479821f8cc19ba242005ec633b9cee620b8bc649ff1b39fe62d57753eec1b88cc6d16d9b0072da9ac02fc8229caaa4d8e8a1cb80d485071eb27186a0b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150ae1e82de20a127572d976e23b8b3f5fa3ea48eeb2589d79abc8d094c18af15b2290c7ea69a0d66052cda94e4550bc752cf24935470eb8b0c7c34700914f98d9838224a2a569254a033365871b4417fd1e57eaae3232479c3f0cfbd895c0fb59ff056771aee33e5e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a9ba18b643b11a77f972a719eb4f1d8a3fc005fc40049e38dbce4ec768e1e0a27c4dbb9c1ff03fe687fe11cb47896392540696f6646a8d33d7fc2fee06016eb828dd3d1215e9d9d44a760ec864b1359186e1830813a225ab8c76b4e7471ccc53159af36caeef0394f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbb3798c5b92353be7242946bd79958682e3ca59c2657a20bb387ca608f4b94f797c7cbd36beb3d967e922f8aaff9d8a3bde7a1bddeb5d9d074d5b3091a60d694025959d1220cbee699523e549619eb06a99d3f0f5e8d3d72eb24b9070847dd4b7039787f7976feedf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b50f3c0dbf27d7656ba3f6e0d56ce498d0d1544000dcab8ee3b241ba961fb5559c56c0023e34e328bb2fafc981f061f0f494388dccd184137a241b83b4287bd9102c2e1170b1c571ebc076ffd5e188ebe771aee88375b54476d9753038db62e0ced5c1a84e2c184ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha76f7fbd7f27021a396d459b5e7b941936a5e88ad3b73c2c82eb09d0c1d00a7aeecc4b143edab76cf58d6e6cacafaad8d96db9dfe14fa2a46681028b5f2135fa6d31537f91ac818159b6f6028b3919320380735f5513548154694962f098223b78de16d03c29328a79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1910615790582d153b20b918fb8c0e1946408612f5e383f87e353667640e7fbff87076b5a444f4312023a26f1e8a57f68c404c19f6cc5318449de864d23296be6a7f35a7dc35b065a28128f79b4ebc02dab8a009f41b9cebb62e3a371d2100e08743f5de98cc1ffb1a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10cafbc7c463de70be06e06510fd8886eb12b6f3dba028bf8759d01d9081b2209c9239a5e21c4317ad290822e41f5e8c675d2f55e17ed666cbb37546045cbd00b4bf689a8382a46fc6c4ff5396ea6fc566e78eb9fab435a844ac6a34f713f6d05567e08f5be61cf5f91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de46fe479d2b1e42032828fb0805643cc3dc14a5d969693ef516ddf0dfc8180684c91cc5a076e55cc5f4c9e64856349699cbd06f3b5465519db4c0d7704355b986c0621b3be268ce62b69bf39b3e0f722fd144f309b6c9d76585b5860988d5bf1a00bd25eabb8194a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf99dad7852259c7bd76a7322a204455ec5159a3748f15cf5a911e75abe062a497a5d74bc31210dc8a94fd1339d50c094d96115347e23c1cf413212f2253bba325380dacba32487f1b45a9dafbe2926fc4233f3640f811251e961500f3e7671624030bac4a56061af48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146949d85b4a0f5a0b38601ae1e7cc4b9df352a56cb62a044b6fb3099e0fd3c5ca5c9dbd6e39c53254fcf4610089e9925e6e4dce2a8b6fad877c6f286db785737d1ab959d657a05b28b5a31ff2d2cc97bcf4a6def5af97eb15dae1631eeaff941b8e34483d3acc1dea5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e58aad5d3a7d238666c208037db8541ffa0990c7b6340d7af456c225a6e8970adce879f465f487670523d46bda98f9ae8e7e1f00bea88c881141f60d1e62af49871f2d4fb4ddcccc499991de898c0003875d82c198bbd3f9dddcc886b1ece34b07244aa025a1d73e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10db4c65b526458057e1e0959fe47e9c348f24dec1d60f4ffe5afe5f1ebc54c408898abf9a367c5f0cc759744115264de6274e17af995a550c565326e19edb76cdc863e4c67e320e309242e331135c376484d6ba97490483a9b0f9eae4679b06af5e141563939b38316;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d803dc688ebf5e3ed9e1770ba67513dca93559424a0eec222be1324edd72cd37c0e77124eea77518781d588c097b089aabd09b6c213ab8eacae4a3e201a4dcae67f0121d764694d7997fdfb31f1d9c72f0c86d187f97ea5800d25f0534b6e3737572c60a615663b6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1e397dac120d5402fc95665072cc0dcbb64c98baebf3cfcbe6729996b17b6ca82062ce754f53711c6ac17d3a1d035b133ab7c3ae64171aa372eef04a9bc5849480ed5d2dd495d375a81618a0ad94df28e722c593c6b262f8f998c3d5178bb34962a31f74a5a7aef0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h925a8857d8dccffb79b607ae60feee72c383c88c4f5a24489014699d80e903625318fcd50164c47362a52c6e9b4fa0ddfdcfbd2a504365338aaaa03fa661dfe3a4ca1424995027936a9b4969e269ee0edd9207829d4fdbe270801d202dc4f429d1a6d9b8d69d5d9e6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b6be8529a4d7787c636d86791d110477deddfdd138ca87a1f0b8e147846e490766233ded70d7e20fcf66ab23f516ffa593c85deb60f7cccdaaf560b16b3937386236b21b746cb1526b7649e1527ea1b19297fa45812f5e5d99f156f722e77290560211619d656123b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7799008e64d25896251ad6830631de6448eed7cc1e2be1ab0bf37c7e25389e1a538fadc96d7609d3db8f42636f99d4dde1668b2c9198093727fa8fa94edd3e2da9412554fc055dc1971d0762a4309a5eceaf92bd02cfb1268ba99df649cff9d1eb0556d70b0b0ca0ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f17e15870577fef7679f7c6abff88bd70d372b427cc5bf55b497d5d690d64aa5f6efa8a3f1526b72a9df61f03d99f1958126f71b94f173cf377aaa35c8575607f9032fae59556bae3a0ab163304f03087a229688eb4dd4abe61b9b89bbf4660c59cb6f656edd90d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c5c448405e317a1bfb2450f06fb5c6ed7649371d32d8f6cd642673dae4b7c27b4b51f5aa63fc2a7f1bb0e46b41d9f5395f5b50debcb52f718f64e21159b317c68e9b5a263b7af6dd31d40a2b28a410a23ac5b19ba6f74f02469118e921ef93b4d118dfa3c2bbac06b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h387455cda385cc12d5c06d8ddbb80acc9788c216de257cc22da1709ca4ed48802cf8564e12a65c51c7b38320a95193df67524c2bf7194bb4455f5d021d7ce42bbd2c0ca5b39e482b57506b6b020b42ce4641d2c87f8cafb7c257468fd8b02208023452212d035d6f86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1268563ce6959375f296dde071d884019fe5e9351b2ca1fa0e2d384d268ba0261cb2ccf77158d5ffaa14c085cd4214fd700a3da5a2c6f9a6126c40eb5650b87045a8346bccd7adecfa4438c4efa0096226ff7248cf983830ed2e2e938cf712b375046e100cbe4e7a50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142f2a329db34e1d9bd6641dec13febfbded5503b476af683c5433636613effc62237bf585021ab6848eebe9e27c1c8f105089e7f30d8ed845fe8f94e1770ab0bfb0854106e14e83ec3eef44b370325a4397886b9dd15a0dbacc8191b01ac5712c9ddbbad9ec378edec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bc8ac8f58ef491c86a97afc58db031cdb50a6ee8afd7ca4964a98cf60545a849a99237350f7469a7391feeb365ba3a44dee58c442c77c0cbf9224c32e9a9fa81d0c97e8db6293c8041b493b958fca2da878d5a554493603b38e6d1fa29d21e4d75aeb2d7527f83584;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h770f9937799ade7538b1be32f7639ff0c4b459442909a773fb8b490e035304214e88d7d789dfe482cd1c53a467a909e8229a2917d081628d5831a47d3ced55c4e1c594f016a3a2479beecbca132e70e0f4aebd25cee06a8d44fe052ec7770553836757cd9cbb217cd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fec6d373691d809ca729c05f9295c0c4226cc095e31a9ff562b642dbb5ca21c8d84bbfdb353d8c15fd3cef9c5e15c914015bdc285d7a9b70cde7f38b29b8b92e5218e2be6924379d0f01f1343099c8ed15104f527920502c766b3b4f6addd18295f8094165fbebea6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8075fb718de0eea7b9c3da5c1d31045e1948f03f65af5e5c51b4784f15f0b8b13bd85baf98e06c0e3df4e7a9e71202131407a3503b78c6954e4ece712ebea900b8a2a68523afc55414983daa2b3a7728f368b2d9c3c44872928a82b15f75fb5722a0387a01e06156d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bfa656405d2d604725847b4916623c074eee4b19e60bfaee703d10087f23a4e2afbb25a0e9825737f35732368c82dd2d39e2ea1d8cfbfd9817ea74072bf51a95eda341d5553fb0308fa4ab5bcd66c140d53e4fa72580f6e112277946675f772f785f64bfa21f256a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40066ede5f36fdf1d0665e5a000ef416a4854e11d80ae3f5e8bd50de2a1840c37f22ade5fc0fd6c5d2328838747c7e10181255f3bd58729e3e52baeb1924ac3f172614bea5d158480ed0ba7a937ed16ee8b9b809ff4ce77fa3bb29d873ebec681f5f393d1eeeafcbc4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e73627d85b59e82c77ee1bcf21145ae55d4d1b7475e2da6a2cb4cb875fbf1b5e16710936ebc8b9f0f27de9386d16013f26a5aa71560f8cdfb4c54543df309861b095edfccc8496043c1a171543b7edd6dbd48af0e8db1a91b20f037f51f057bafc35576b6be6626406;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5de8b259e69029e8ce5fa51f42e11fa4e122fa710bccfcb71bcc0003b5c2efd824f4f73ef0cfa18a06bae73cf189e7294ca8dbea93c2cbb5f6fc7becfe6833c6f26b181ce5056be9b2fe812df225b6c1a0393ef4fe55a10fcc2b00e222679b136ea732027ece59f6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153acae52434ac7ee5e0054b16502b3543b0dacb8653f73accd416ff6fb74f142b2d34997e5e31b9407b029404ef49144b6c3e6147403cfc35dc4fd61e89d5634785b4191bb13e8b8ab847c9bfaee20f0930cbea6e3fe80a819e3ab1f1887303c45ab7f0b104a16dcb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107562993500db4f9454e1ca374e6d5e1c47670853d44c71285a70480eb713f03894848319f4c565b33209a6606a2381cc03c02e039215ce5338809385ac63b7a79364435d5e59a51be7d4633773674dc6a348a4b9081d013f216d9382889bb6316e226fe2cab275db0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f333745127104d7f361f3c29d1eeb3fcd16bcfb80f6a4ab3fe71550c7d5548d10dfe11efbbe58206974bc29d5438473eea34a7c8318e3d0cf4b20d865fa43b2ad2b44a2a9acfc1c7ab96c6c79094fc6d5149f2270436ba27b20886c8f49141d2c0c05005e8cdaaba41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9c19dd9767dd6b8360072cf03e8140825bea27f8ee4bca1662ee737aeffa10fedcf051eb1240401072a8866b970b21dc1b92e9a528eb03efb3317552e8916721c20a243f0714799e59721cbf190cf63159a48f05f6feb26ba708d97c868b9eac802aafcc99f71b72e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e230b0d5555251c3a2f49ceebe8a00db5eada78842a2a9e1ac29e37fe7b78061e12b4eacbe856eea5b06edb03e20721c6ef51f2ae6f79b61eb823acc5d9d6d20764f68a680afcaa386e4853cbddcd4c33d89882a434674cbf5f23a7c5c44b8c33877c74f43b0e22a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1089990619d3266c021f8db83cdfcb8a40bc19a407ce4e8248a668acf7c03a2df94a228d904cd34e10a1f86fb58dc2d2b23052b43091d5de2feae70f0de65d16b54edbd54957fdd9af21e2a114bd7b88b64ea4be351dbea76e64266776f438422bdd07157d7849b72dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae0eb06593ae0135d9987298d164dfabcd95bb3ccb7cfd1b1ae983c2d5f4ff39d657b274e9423aa24519dbd76cfb568cbec050680f717f47c4cc77f945e9fc95f5e619aec9bc76c44ffca43045ee668a94bb39603309c04a3ffc95878aad47b50fced16cf52d2e67fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdf3f24831fc45635b89534442248ba44ab490bd12dd100bb6e4f10c6a217919f35f5c6929d52961ea9584538e44e45ab0ac19d6828a4543449fd75b5aee3c0022568c4cb86a6a41203c167526f808c3049c07c8888dd37c3c59bcce76f8202f2f1435a7301e003abb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff4deeade42fbf5885975cacd34e011eaaf774a86f538affe91bc5f85c02a6b241982031e3c397f15183996bab21618187b4c755ddab312916e32241dd3ecc6d94f65fe18486704b093608be98e037e9a18b43554a0a8ea476a96c5c97b546034694084b3bf576ff98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13008f7b292ca48e847ba68fe01684d39198e5483ba07eb5155907e22c0d3239022a56194dcec3b5ec9b06677848b56e5af96a4321d58f9fc43a55baa34d666d8da6309ba6ff4a77eebbfc456676db99b973b475b310495b83b8bff93bf4a61c2799b9d017264ec5c10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147e1f1d7c788e6209fff83d059ccf9e5b1d1907f7b2a037cdbe1ecf5230de4149fd5197d87b838431e233fbc849bcf1aeefb4f9448e55a09d67a3aec6eb5eb74f82b662264a0e994d994532701a38011c7de7a1aede61ea36aaa7f46108231a64a6f6c945418356a29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e509d9f87bd52db125faf252dccf8c3a197a4b19ca63e2aba3f2329e0751b21df6afedb88760191c834cd7af9f53c9c3a4ffd05a7ab4a95daf9cded6d899413f4a03e8f7987cea40c4ad57fcf2dc7805273ab94073c3510c7915555216e6ac003ecc740624857cb838;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c8fe4223bfada109523f644a86a7b4e519cd210af30a2c526d8466ab7cbc11e22855c81de7c92147122753910eedc76e74265160ad3e5890c49765bab480681f5571d9791333cda4f83c6ce06a3fe93e21a2b645ce2de9352615fe4358354c7f38a06fec83cf120575;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158fba23cab1df1b0a691ac89e887a79f2fa73802a46473cf203884ca206747de240381dfbf196f2ba41ca05011c23e99d6d77b10ef7a496035ebb68f16f84aad889950141e8872553de7fb0ab249d38182987b07d178dbd5bb641a771dddae37858d1753bfdbf4690d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4202a7fc48d308163f21fd2e4c8909d0dec2f10f61caa6b86f1f77d94b32e7e06e3b198a87dedbb4dcbba4bf566f00b69fe9b36c6becdaf14f0ede31860583867ee7dc4d3fbec7c0b8c505316d72bd044c7007316a2d8a2f296dbcd78ca53ddc87e3b52e1bce7bd6c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he31b633c8e11ab14b022aac4628150409b8cf04ebe28af0fc2125ed8ee29aa9b130cdd6552680316eeb4a84d70dc3cc364c6239fb69be608ad98236896ed6a417fb2fa5a94c79b917a156914af5805650ff9feb2d51de8bc09653cd26cb0649b9459b50a4becce1d12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ad4dca2bf4bd72087997d08ca8d5ea8af8bc7446be68aad425569e4b29017bd77af5b872b30b56b35ccda15f03eac94e3aab46a964a19ba51752aba8770ae8f52fb6165cb9adcacda38463067aae2513953739ad5b4df24437b99bd19e168d3fa894de2420384aca2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142758970b8816072cb87734011d28a926c3b8ba6014bcb9efc2ba76d631a2f6fd08bdef3a5df394df0b183104f23ba7bd6ab9ef7f2725ecfdf77496d800e5e989c501ab229c4262e6f69b0f392cbc44254444eb383b17982ed6a3bb49e47c535ff1f877db4114ab70f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea97142439d63e8f4cfd63772b6457cec148233b899c65ca79533e63df78363a25c33cef61a6a240a2c02d023339783ff5db7c406ea44565b4319e310ff399877a5356f2582065e83ef12dbe58a09d5d1608f0c12864bdba5029b502a22abb147a9c1ffc428a66ac75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a4ed90afc818bae6b034c8eb4c686ddedb9e22dfe4c5ecf7e3bf85683a54bb0cb75cf8ee251314ee930b1b0692f45652a5af9075cb675fb72f5e8fa1528a5ee9868640099f6485a5da8872c8b7b012f18de694418f82d3ec6f3812db618758f7c00d8b63f139fc5c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140a9d0335c2634a688ac1383916d337158804dc037407258a0e9eed75f55a3444801c6fdc0aec66608d0f6bcf4716f83203acd34571608dde5d12c166cfa06aa811fc5b644f07732766f1c932d4a6fed9b67565ffd30ecb1c13282c46c3d27c308186ebb540d0f6076;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae7573efbfce7cabcde90cee9a3a85009ec4641d8ce7ffb481d9c24c385e7d5eb3e356df710851e1ecf59460c28bea9ca6e9ac228243eee6f32b1158c49659ea5bd7991edeeebe1fd9a8ab36d4adccb0e24c9f3163056052b3452126a3802bda37d46c5f287222eafa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17447e1befb67a48040b0ab5b35d918649dfbf3c7f3a6a8b741e6b4fdcb5493858844dba31ed89c2a4e8b032bd851391895ad624f921a560269bf498da5ca8a231eded2e4018438e9feb524c74c582511782a5c364c729dc1e48a949844d25e07b2c98aa606293c87ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fce44005125c60ac751e3d15e3bd52e8747c51b983d5aff352f179a792f6a2bcc9c3f4f756eef5e9dfd0d5235f3ec091fbe38671b66fbfd8e359d8957dfa0457b7b284f3e1a9a58860d3813d1abd90d43c574e9e92450cc59c2177d5118d30d566cc2c9a03e01331fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffaf05bd80b962d22b1850fbda09313ea0d05df89d589009f77f1dd20bd7bee621329698dee2ebc4a72519944e194a927c32f49425f7706930234c05ff451334d84e50aec77b3cb86dae468349ae95140e45d60adf491ffc7c4e21eb72a57e3860d8147e2096d209eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1532a1fd59d66247a0221fa7cb743cbea0d7ac454b88931df7c071f6aa693ab790386a503ab9b37dd66d82081c60dfb584256e7b5893f9b9d30863332fa410acdb162f3ffb29945b910f48135068756c58945a5addaafb888bb094a48cd4262ebfab3709162a36ffd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e11a09ab9bec4a7cec151a365ec0b3e4cd33ea58786a8b76fd112378a57620851b8b90bbc22bffc99091c06900040ae135b422753a3fe5c2e4f558277854b1538bf9fdfbfe4bfdcfdee90dd705e6dc01ecaed921154d650d2dc4089105bcd393e64f75fd6958b5f15;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41e3387eb942d84b8b99e0f4ba6ae850590fe62eb3baa82019ab22d11f20587b8b887b1a285794f02924601a9d3524be652a7aaaacc9d7a4bcd77000ff946cb0e2503645f4069f4a2d637aee886aac6ae72355e552d3dba804cb9d788cbbbbdb387092c74252e22315;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1619b776cb418c3e1206a391004afa06862d0ee3aea6e137d4fe7f9f5c4ee6c8d68c60cae7c7b8be5c28cbe1ed772cd7c1e1592dcb1cb691400e84187846fb3c9923110934ee264f2f9ea517ff86ef854c2c89dcdcf7ad3fb42badc9419d0b30d17e5fbf4cfc4bdb6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50c43b38aefca40d98ff467af72fe00089de9ba7454937e71d90f2d22ed0a59b8a9adeec8cdcfffdbc6131c54d3f1b8e7495dad95fd492fb0c4e1341a80f955d327b9a81d87b2606e1b3eba47c9acbc1c79279ee551dac5e76a4596cb0eca6c409c2376206475c58ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83601e9f51787fce7bbceb52a7893d09168c4ea50b20440bbc910d541a51ea80cd2f8186807655961e4ee7e24eadef8ece4b6e23efc33cdd62d19059b9da1aee8fb5d4ec04c5b740c43ecd513c1e88dd3be08a086c8271a525b2d576e19d0d21a20fb2e3cb10708c44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41b47bb0934ccb0ebc1114bbe384a7dbd5f130e5c39f617db28c5a68b7648a6cac26ef825b6a4f7a5d4a12c39f10a8338227fffa5a059d7e469aed7fcc06ebf3920278f56d188ae01797f99a0ceaa0fbe92c40493a83a874ee77929766bdb4202dde77fa1ee406da24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1c532bb063b165bae97c6be77d8843e9e0a622f576eba27151d72196d027fe9f87a5a846672142fe7ce804f38e1b36617bd734447bfcea4b87d2b98cd611cf50a33202547dc72db6fee89cee7c5945a52bde571fbd65147ef05b3bbf3de5ccc28a641c5458415b97e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa55bfb2f1a5792422cf6f4f38580955602cdb90b1ad06330bb1b73404d364afd3801de73ad3cddc754ca41646b6f407b9a228068f21bd69be39e107b45f16109d3ef526261286da0c32e246daa591bf161ac975b1703e6c376c2be959b1252fe28c09ecf752749600;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11600c8eaa75e961cbdf5be96df26d108750f51fe3428aecbefeddf1ee3c64d4ddccaa0f0a7c2e47c1e09b17cb6988389b979f94223e83f5f6ab7b4d91ece2d98fe1a592e3e987c39cd6c92149ebbce0fd214661c6bb90b1177725b5a65c3abb3c259ed9f28c72d4f84;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117a80ef28a000f99d7ae837b7588cb8fd699bef54036fb96eeadb4183dab765922596e5bec689da03d0565ddd4285b369d865ac478d29e7c94315b8862c017f18c6169210e2fd535c65def1c4f77bf9d6cf59cc8d733a1281e34fb460bf711e5f1c1c98d7fbf7c4eeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h712c5eba712c072e5062caffee50907e56bad941e186e0dd5bb767aedc75a52ba46a93f7869f99314bff96aa2998dd9aeb31a0a249ee93a5302388d17c24fc6ebb7c081c054223d095faafd9c3254151894f4216ba790ea92dce41f02827794cdebd5f4281a3da860c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14aeeffc2fca86e5812cd2c7e287de40f6d56bfed99f8556a46d528194e69b8961dd49bfbcfd1bfe3be1adf839f0cf6fcf46cf91cdeeb3585ee066fc8dff70705de5ada1786d593ebd483da49a1432a4192ee0e62cecb2b4770bb41b411075364350b895e40322babbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0b532a7401e4c9401e14c028ba3a6076ee13f6607eb4a6d93ad5a63b30548ac943d77b47c2d46dc69a14d09a64ec7020474ca7c3989f68329aed47352e9950590e464c8046a56f17539d723000886fc90be5f809d0161eafc2ae57c0793ac8955c9a089f7fffb849f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12fb02d9cecedda59e2d9801ba22429770b3d6381d5a5ddf6e1c7dc8ab1a13c22838c29d7d4fab298b426f7e98506710373eb286d1116dcb47c52c062467001c4caf74789c1617a21ec79673b7f1e14ffe5727ecb3dd8dc95742e014d476f5fd4b9c7dba2f0572f27e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90cebeb17e96236cd7e313a046247c23837e0574c809e67175dfc39557a142c6e5f00d324022528434897185b7f29fcdcf05897941f0e3eed758c1a052c711d3fe6479c301755e98b522d856a3df087fcd291c3cf4d8d8152b8e34af9c3a73e6544ae7d534326c6270;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1aa0dc0b8554295b765ea2a6ba248edaa0d8865b2b2cb4f7dec239b11a7b7819d66bf976cf9b2dbb527cc638418f79a5c63c403a8f40fcad8c8359594d8dc19c260ea4ffe9babe8a6f8a87aeee74f721207c241ec6ffbd49db6878d3f3faed3b43e02bf59b59cfa6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc736cf2827600c7491cd09e0cac3acde4ad24bca77d94d9d172b99037e1c9bfe758f797a1c8903e9463c5976be54deb04cf45646bbea72873a796a3e223abebca6410dfd3de3d90b27667cc87f5ec68785778fe92ad92761b1c3d1a485201d3d7a60d39b717da329d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b015d6e861a1668a7c3acd3454215a11e64a9ade6b9eb3a471740ddaaef64a2b4ef4a143eacbe17dc5057a585621a11e67b9cd03af4c631a8ff967f55986ee7a5b1c7ffbe3c66a1107feec37f9dcb4d2d23a5ff1019593f4da75179eae644c484a316025db7bccaa6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb75a9600b515d2b9e30984206c8f5068688c231c2fe9437bfdea400c7580e2687386fa1d6ba735949d53623f73eea573f53497a29eeb71a0153fa0afbc3940d2067540e87250a470d46b32d4aa0235a96c0aaeaf80ccb4b5bcc4d0c695b356b4f3bc32015024ec186a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0e2df809bf53893647342ee72c70342b9c96e844d988cd242c0756317ec2f3704cbb10cc375855146699d2180633feb835c7ec032a31808f33ec83a2545423b5c6e20ed3a69ca02c994301de218ac2c85abaeb9f831331a0b62c0e345e39b98dcff5c10e5ccaada54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27eafa01011d38995a3164cc812a62c834c54f59d8f76e1603e9d3003065e60635af49b5735f746648e20b61288f129a29a3939d706a75114e227eb67de0e0326136a66cb42640d0ec6ec824277cba919f0691304cd871884782eb104030a6edfb65d0267214536b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h455032349f115da1ca6ab9efced55b6b756146cbf8b0a7bbd68a5d2193f57efff12b866529aacef957df0a280ed377b6a9ebaf30859ff482b3042618999344be963c005539e6231e3e4a16c005af497fa8560aefdba8b299e0b6c9907131c0fce001cdaa2631e5492;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d140071e69f11894f8d01a899c04873f9b2ea7beefac8f5605681e90abf55fe414378ebe31409fa4c339567d829d7f39a1855e1ed63025f58a3cecf953bdc09fd3a24747203baa122b407aa99fd92e051864d48fff09f49493c6e4ea05171807ec435a18ac4a5f7c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e669bf5833c0512c2ba41f9f02f74ddad2fa31539dbcebdfae990c9b5a461437de17b30b6477dd8704719dad744ea5815b51bc531d309214746d1a3550ce357e7ef98e8c9c4538c39dee8641e23daf3239caec44e444878be2ddb3aafc5b385103320fd2f2dac9c392;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b15a4404b413fe335a5e671c180bee73b146fe745b7b60b41b6cc8a6167b0ab1acb780e5ef4fb9e6183c39a1f1716c1f23ad391a1dd83c0f5ef01a4e3dc45a543cfe2f9416c15e630334bd155e6d783900e70ea190c7f631e74b36d934a04d011fc863f59820755ad7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf963684e046005765d7b51f43402bec171d7cc9bd6a19f1db5b692358ab204bf2505429e45a962a0992da1dd3fd09360aae82495775942f7cfc2eb8e2062240909f89bee2028ea88629ca56975aa4e5e16dd4909c98ed2f780c2693236c68f6be99389c1bc0626a89a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57d527294f8ea5d69b533cfb75990224508c9fe38185436cd4e9de169929a90847962987e29b694b30846cc7ece1419101ee4094c508c77b854346e82b7b4f9588ca89f63182d21bcffc2d775162129d56233ab6fba8ddd7a4b42be5e4eb1d21fc23e759e35f974df8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1276b551a54ab408b82c02e4d3a0432dae9dcb6fc9a3d7e73559fd1705c93ac49faa64841c606e1d58d286730ae101356b516e427a9e795b53c507c55fae743e25c7212e91d6ea5b3754c04b9aa304dbebcbf915c1503061db6d7faac738f2150a35620dd016f543b99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e980a32406eff6619756243bfdb1aa4eae1e79c47d606d3be771953d797a2491b84c6c6a3a0f673baaa06146fb0df7590adca122f7c476fc5a559e67064bc92fc8ef237bf5698742524a223df27489f6da19c0e876a70a216e474c83fab78ebda6d8e2c32e2c10ad16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145c66cfffd7077b14301ee0705797acb3b018c15f44a3959ac28dfe2dcc89bfda7e8c7a4a7451600ef89b0851136fbc44b24b5f930f699f779bcd010905a77d7f8bc7b8b12982bf2b31d7e2245a368f138d7001d4c5ff04bdc3a360a2a1340bac0149633992637c57c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h201df970f9b78fda1f34786a266e0a478622a1fbf99d4489f3824d781830d6a1562707d03a898588dbbcd8dde7f3d4fdaab7584fd73edf6f40a651af0d440d84d7cab18b735a7978c2f2c20964beb019ee26198abbf628d2da0ec969f11660d61eaeb0300f9b217016;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b630e8a42502a72a8a7609b03ef523c198759c6844c198efad4555c71df476d086695962481d92beba9d805ae478fb651a5ca3606e327ce85471fad9c6910867bde02c751e1af126a278db47563cf7709477981a4f1fd614e6cb6d3ccaf47ecef73a375b018b9068e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f323a0280056d84955cd7f60245d0d9730c47e92642106e694239d70444152fdca288e4afcf6a0683ee5d2915842b5a27eb5886dc01af3786f1936566e5ae2f526ee623f32b5300f2c0f87ffaae9aa3127dd3d934f1a3b233607ffc4687796281f813b201e2a43045;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e36ae633456e603e6e6dcf62aaa31bd07316e1dea9a0fcf0d1405fd39fb09786d1e5e140d8d771ba4868b0428e8202666468e527aa237187983173d4cba905fbd888aa37268c95459e7a3ee1c9ff91603a2434d74ba1ef844ff11af1249339e58bdad46398beec0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d2d98c8bad18b314305af354ad8e5d466d2e1ac0ba8b934c23cfb1e6d534cd2f5bdb4bd29e581faf408e8fa445ae7d068b5e80115a47ee93a825f218674f39a39663eca7112535791cefb946999441bd5ba8969586f2191f521dee511fc908b044f4f5049a2b4fe51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141d8e0f5b7a13051830de4808422ac30fabab6f82cdfa4d72d6d724e69723b515d89ac725505cd2cec420177a94d62ab921bf86ee475d0bd0cce5a673a2072b310fbed03f82b7df51acbf4fcfaa97d41b0a3dd370fa33c77dca575096f07af1733005edc842da17b7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf94164611bc55533948e58ecf283f682dc4b3f7cbb86ae3cb66d2ec115dcb0d961eb884b82ce493f75e4946bf8d9c27789245494a84a610a58e18c2e9efc58eb94e481b2e0d9d9d33a1b92c13d6ad124c48cffdb8abe232ac12dcee93f8de2e6485ddf75feed33de3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1612d44696544169de5b83097f233868336b6c715b8e37b020b8aaf28ac75775bb291c1b64a0c4d77147f9aea3766a197fa78e15e6cda319ab5426b3379c851d996226d1a1739f82a52cf0af482da90b6981f53a4faf8ac280ea9b703f76f2e5b108703df66a268481;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1276b446005aba400c053dd8b973f80763dc25d7a3884a859791c92fd03406a054fa2c619473046b5cb890179e865c62f20aec8549cdaa896451f7674dc206db8b6a9e9074818a6e8e15b1a163101f648118c4f4144e6d518e05881a1d5e0cfeb5a5c8bf5147b6c7817;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb4f650a7b550bec06ed8d973e1454e8fae6346b067b12e6e2a0f0faa02101da271e0e95b64c22114078144b1715912a28bb484ecb52ed853cfe37b16623f6641bdd7a968f0e69615c18c493abcb01a7ed0b0b2a0ef40f0d0fe2b382421ecd838f7ef816ecd24f3898;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1256fc869584d3e8f16fda9c3827c5f2554253005853cbdc1a7b0316e250d650ca282c65f4ade9bb0e2fbae91c695ff5174777699a9e8c62071d8b011a12b1e33e15fbb12ad0125ada420da07506747831ff5aaaeaf11f8021f881e84e16f38fd474b7039c86fb33413;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147c48ebc825c2fca1761a9dd299102728727bb303839aa0a72966bc93e3e6bae07453d0111e91e54eb4fbe7a70db8065981d192193d5fbe63e5ddcebb7615afd7956d20f8ddaa5cb57791e7df4fa5a876111952b22fea2f07e02ab77a503b36d70423d1d2bfd396e9b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104dfd7fb6789dd62866bb71bc992c3befa90e517611fa423cd3550bd393b3b7bd45ab9a357bd0eb6fe874b18c3fdc37a8a31fd65953762e32d7814cd5403caa5dbc6c1b2a25ba047aa85942b7fea8ea946b1486e86c24199f580cfef593558ff1c80046e568c9bdbb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20b736e8a60ffb2a0d0c3cc014e3b8d4534bd269a11e5beecde045064709659ef9fb262753a74a8917b1f21dbed616fc26b900d007d6a4a5fbbd78abc5a657ab4c4f4d346b5e0adc76e4f5c7e7eefbb42cbe67839852e0f3a5757707ef59af0f0aa3994b462904dbd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1732bc0e621159d285f92481759d82b7616f17743d9cc5b94e3cc5874a19276ab3e343b43144c4528b0a0db6612af1bc4075cadebdc95b5aaaeb8662beee270d1c4b8a259755609928cb75de7385ed8f33db94e57facd4dd56c4d17cd57127d57e325fc7e03c17b1172;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6431e218b12c7435f2b3085ec52307c8f55fabf74bb4b3a48ee874315ef976b0dd490174c92c3c3791687680c902bd5960c66b41e6ecece797b2798431830a3ea8d464ddf5109eccd1d73b1fdeeaab8ef0c4640e32ee09a051ab3bdc262de944aa5e5d7af7bd24a7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6499d0de37ccd8ba0a87dc304ba81f80ed432e8a3f1a3f3c62f3ca363af2e50401e0665332cf7f42e1356a3c222a28a2b3534854d945c7303e02feb65445695c7de56e12c203b3162fa8915dc683ce9bcc437cdbf36e7b3e6fb2657a02be0c393bd71a4304559d853;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c64a133067dfe29afdd9541839327b69b9a36b719a908918ea8a532bf4ebc661682a85f8fbf9385efb72794f45d751b3ec41eb06f80ec4ef24e9de03d6fe543fbf3da9d1a9c421469fe916f532a6ad9732d3af220e8fc275f8852008a11fa3254253b00a247f33f2bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7e87e6408105bb10f7c9d914f1f67f61ad125fc5ee5fc957ebf85263e2a5fefb578eb6ff52de79a2e2469ba15c5a0d80f63f752b44fd17c20bfae95f32d4b99c10f65be6732713d1bddba02b2b61c374d6a69335ba16c24d20401f88821931b5d6bee2e6f65842d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbcaad26856d373528c2f2c28792ea91a58c1ff83aa96e3e7b3814013317d9bd399dada9c29ed2ed9e2a1156e329b830f3d4e21edefa608ad54c184d663ee8036278a9ea4418faac4e1c9fdb6b1545d4c21f4223e9e6be081e4b2195d6cfbc207b83c89a5ae6ff3d513;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd53454c708c4668856255a18600d6396bdc2cf86a6786bac2e420978eb6d15153d0f430a82d96a6953fc55d6475854ba67d2f94841e87f12fe45dd5dc19728663e0a325b2aca54cba5fd7a162535fd2f1cd55294993ff25f187eee190c9dd9bea741dc1d83f8a20db1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60d86cebec98c5b77c75c35083ba0b037affd6d61d6f1b1d933db77f874f87f7d1a777431d3dc98210c995d6056dc79b65b5f03fc861485ba59eca7be410d444f1a4d7a7ec4297bb0e13f9ab025b5a7d4a1c933646b1d2c49e0834d83a6b8cc5bb4fbf5790c46f60b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187649a9835329324263f4ba745e71cf4a782bfae573b1744b9d029cc64e2134a98b26670bba838daef2991573456a0b83f913dfc921475cd3bb81b44e0cae9574c93298318c7e28307f195c021651a612ac253fbaf96d3a470b54f15441f04dee5da6cbc0977dcb126;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f6852eb3fc0986349b6036ce2f6b26766403a7e872c6c260d43253aaac18be7e8d87a73df838af6bc2a7c415cdb4d40020631e572a6a2385b5cff81fb8684b8d6a08d3a1830a9ea1c3fb77d9b3fdde22b40226fabbbca562a00274f65a8eeb3a3ff0f947f0f36d21d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb32fc40954093b7a6dcfa974aff357445cc5e8e4804e1419bafc0bbfb346a48f83773ddeddbe2ccdbe53c85333e61df904d87c7b87b8b609cd07216723d2db7acbe6775864d954ff91464520ed04fb59b3a92c853ae926687c1745b5eb402f4593f5d7c039f61b0d92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ac2a14e014b66bf8e4c2fc050a4361fd996104a51f3fbd706100fabcac0a020c7ba271bb4484ab9e1aaaf3014c8809441e3ca697e11b39afeba6808d0bf7af5b7e7278ecd588cae574dcbe42719f581f344c4a82a131d653d9724a272fdb4ccbf2ce722a3c8da46fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h942f3c77cda3eebdfb93bb856752d9ddcb7fd08041cb4fb1f6ffd34e67a00a7a73c5a11d3c972b734bc67687f51aa2a67bf009e8c63bf8600c94694d3060284187e085683a9539fd865d6db82bb39058d761c6030acf02f97f737a352bfdc07eb8a0f27aaa16ec14b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hedbb6d8b7c00b9862f90c67de0dec15e02f1f233ffeb8ee103cab7ea5793160644954c9a6e267c25003bace4fce08e248edbe8c92021e8d411c7fca94130f6772ca86c3cd0ae1eae197a4a24d57ea841d5a3846e66f6c6bf22506bb8c0b8c5f80b993ca402f7c6af4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191b5b5678f26e9d2eedad1fc329e6a4690bc0d3d4a28d460c5b41246b7f8472eced7f37eddaca907368b9aaab6a870b2a98268e7ab2e628cf1bf8a5536906ce1319a9907e6166e331a96de1cd0d6c8c6953334dbe5b4a70a8bb5c3ee6dac24c3e67a7efbbc48d4dbbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc57d0d98f46164433470c52b021cd3dc88b516352610b873b9b8a0b1d9bcd0417055a2787645e429236b0471ec62b32c7b7b4d82da9375c5489fe596b006f9c2a368a92bc82bb1e2fe8301dc0bf1e3042e3ef199b4b481b1c00bfa4e20ffa6f286c7acbd84f448a496;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1771760a9d0f26bcca512bd40d982ae18a27f6817f725715e5a1de9e8787dd11befa1baef6d9925116d4600531b8b8877ebff3290d87bd94b702ee919e47b8e9af3d83cb14551e0d951c084c5cf2df616ca959afae041f7013f680bfdce08127addc788f365623e48c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15165da9cf1bae274becce3e686d933def0d85e053c268dc0166124191dc24f4fef36ad636decb5d5dd4d09d03ea0e963434ec9f61d9c28acaff133be0d9fc2096289c6ce2c99da4000dedea40c06a164c40a2320f52969ee70e3be8e3abe93a8a581f74ee606849e59;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1522e033bbbcefc59a01b9864a955301daa78a147007a5d3e1a28655238d37fcb3287e622def6075a6388fd8d552a4ae707659965ea9df2ff898c77e0e540e911eb0acd6661f9a19d7a3a594fffded0ff2d5c3de1275d45903523e598548ad6b9210b3db09e6993aa84;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72e2e15a292238848c844f120b87e6847021159d84c35a88f7d313d340b9e5a44ab770e6eea45d55b4a75feb5ecf5d7697cc6549c1bff351f4859f0dfe11966ade729910dac7580086dd3e66eb0a7c5b7116b25775eaae357cef89d90047a90b46b3d7207be9b237f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ada4377d3916d40012466dbf29fe4074fe8236a42e034df563bcfdb61220afb489abd8f0e30129f0270445dae8de7a1a86c4ee6a399ef227b6d9aaa7d1ffb9b46e7a8fbea9995f8fb5f9fed3106482e4444ee7174b449c7e2e7df2fa0b7a694c3b8bca9e25a4a41ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea70c680f66af2a7852e90b3d2917c54d33649af7f6624069d8e139b197d069a9e02bb734a7f089d2d42f24aaf3a34e0f14214ae6bbf1831e3124132ae26f94417db1a8fc3e890006b68aa61ae9fb54e69f8f6394867bf3fbb304d93e69565cb31915c84d3314a6b9c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3c5416560b70c176cadc63c42c1e403c61bed7cd727c63cc64d7ca9df0b9c8a16ca9601aee102d1e8f3a3ea373f916df361dbcf10c353dc3da3fe88d7c933269696bf6ad0ae8fec4ed3c0fccdc7d7e2e4be4ace2b5871ef56b32d5342c26d84068e65aa8aa92c8e50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6a025e31476fad14f85ee93f57ca59864e779af04b1689361fcdc506d10fb521be36b152829858e58edf83db18b0a4cd6716b3c05235a30139bc2ab65b9490a62c6f69cefa4fda0f9e3a3c9c14b4ad93a317c032bfab7d16fe0953d70f3accdef879eedc30e3a9d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d1fe511b477a7bee22f20f7a07c387a3b8131c0146080ff2944828c86329a098d34f1119978fb632a5f7d2b3d1df8ccb2728b08a8f861afe7dbcf21a9a487652c688691c7030979f314f98287a5b08bc3cab289716f2466b527a2773c39bd6aa2c8d4b06d1a717ac7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19effd453a2e415a34a831e7d8ee09905e352c4829ed35e9c88a0207f9d3bde643832c86095874502e152d56c0f9992a99f39cd960e399ea737f77d25811488dcc59f76abed783c0e30dc38a48048f5b3a21d10a47d9e082313534b03e9c88e2af6e352380fa6c9bb08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134747e19c8cc3b65b2de863340b55ab872640be10021ebf4d2b4303bf1f8e190d570b38761a27160d15410141b7363537de8b8683cddd1502eae6ff4932710593af4f7fa0cb5d6bd3120f3457f2e002f277a39ed8d5dd81fc0ecbdc0b1e99529ee20ccbd9da9c75ff2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36de3926ff85f56490e66b35b1e373defd003426e658a301c50332779cbc266878e7c2b9f62988cf3fd2a74829aea24270b2fc5cb009c851db6c473b09357fa398504307fe53a71f2a6582ab041b57c29f02d93d1f8763407fd7e5cd69fd43b45e18d64358c1d0dcb4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he82f0918de202e584f2175e8d74df9ba6a28bb0db11b95e6e3ca0fbdf16bf61daa0174a613e6b9dc11ab29114cc3ea3665d55e104c624acaae6c5f5e19f701a321f06ade22a5f08cd96d21b03582f64fb69f4e2a5ffd2b37c7cc77bb8bf1b8e379fd4f9069a4f43c5e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148ea7b7b4dad6153067adf95ebc542a5bc8cb409978d01bb8b0422b0534011f14fdc01e7bcfd3f082066fe5890acd67124ab12236db3c6a647ad5c7e09745bec46baa6fb811f33b8ad3670a040b523a09c598c62142eecf61f8e3c2c5ab5fc5123160fc0f79f73e684;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cdd167c4d3c9fd0e951a6e3ad86e16d8ec261c2dbc919d783247ec6958f312858473685e73093aebfc2b090b52e67c5e48ec889b4ae87b18de44587e4b1a2b989679147e641aa1e41b5c7f477cb401103327dfef77b04414f30e19aa00b00f389603b7ddc5c8365f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf56af2297090468a5b4db1c486e888f1c0152c0199a5f11de3d17ce1c21b3b2d917cc842d8849d1cfbc2d6a9b95130835d9b224cd0356a5c21acda06b849d1aa92f6a63f7401f50017845012d9e6f39cf0d257db30cfa856c0a67db8425ee89a18a70c2671f09e428;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18209f253d200b1dcf76ab14e3c39cdeec714c61e5260b4060b2230ee4a40766f4576fbde1308387c1cc69394e51c5035feca103c2934fd508140c8bef0bb68df8ddc6e02d55a2f9d9c254434203265eeee5ea57da69810b87acfb53cabaeb81b0db9a2cf66eb20853;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d85d2ebfa4e6c7b5ff08a39df7e22903d153bd444ec603b3014037292d9bb4aa40cc1ffc9c57a4353625246ca7c602abf71d4c28498735564939c5242600b049ca54a33d378cb013ae2597212fc942eb489738e8b510c273ab3a3df62b173ebc1d395aab9ef457ca3f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9b172fb98318de32488abd1c9bd66a07456c13b8d58e00a6f4eb3c3dff928b42dcc5215115ca77a4a9257854e150665f12843c42ff9820da32f462503a2cdb9a8883e5a4be9ffe3904ea996e72258d06c1aaee6d46f5cd330df707c13cc7f48d8af5a026e51953dc3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1407b1f2bbd6c56bab22f6e59aab25649c3539f044edea09b376634ea12e53f45fc995ec9ed015d7494b9d98b5a07669f2939c689a55be5a4e46f4d3f75b55d955ec2e919942b90681e91f51800378269166670540a170c3be4bb64002c4583cb7c6bc3170457af308b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ea0477a7db2310832df394623873aed08c2f7f50fd9bd7591b23f345f1f950536565cfd796775ffd29d2cca04e987fe7297a6d725ad3de6961b164c3329a7bd90f841ff4030b7db52207e2b571a818ccf27d6bc48aacde4f2ce9e425efecb5ba821f416df6e776b03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1504c760831975230bb6bf82288babed2cb53c8ea415136e6b8b468603fd9d7719fc5a977d02f51ab477e6bceba1233fb9e9a4f1c117326f3d21445dcc0d9ac04f72f4ee30e9d0b8ce027e540b2a1f63f7c5ade4b1788412496e2dd5a6190c93bb62b0164d7aa1ffd40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187c5e8f40ddae0b86a4217358c384a487fa14272b0256f6513e56debfefcf9aebf623b0a0afeaa1e49a9d79da6828425dc4075deda832bb18242c22c4be93ab2c50636e9f825ea7bcbc1f01bee0bf9492de30eb2e9eebd57e14cca71948fd708850105d7646138549c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76a581bc07e1db179f8eea09ce2052f0754c8112bafa17bd5a01b18cdf6e5e3fadf21265c2108860397a4c5f7316bc8465c2c22a82fd921fa1aa491a97d912f5c27ec00121092987d2d36f3f42b26b276642c7cb0880a69ae1715d492c0b547b6c87debede86bff4f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadaa81bc0e196192476d211e82104e7ee878fe63fca87384138233023965413410c27e15bc35910373db3a4988313d6503630679a5c59f869dfbf71c696b99f411507baa5503d0b126cb4ea49b5de06bdf62cbc03f6251d12e189ba0731807bf1ed94ab3a49349d143;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111974bd44b7ed986b479750907782dfe8177a21d554615d60311b3ae40dcac5440f4cae6cb413a8d3a8c97eb9ec926298b98c273366261ed771df1a049c9d31201a6be8be18202333cfe38cde1761730d2ee8d9123b6a9485a20bc994b116b178f69bb25272c837d2d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb096e1d4d55e28aa71c109a1c49c395b9dff497b069e97efc29ddd25b53f6de0cd35c8f359360c1514a04d4812f5a2f9e8670e28a2288057d1976505a0db7906e4e45e2fc41b6e26ff228a4886a0a903f58f9700cde6632aad3714f8b8cfecc8b3006dd361361fdb2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14583a36aac59187914ccdbdccf85f41dd665d6dfc0099acac1d764b07c555ea26ee641e278aa834f1e1eab57fe40d7220bbf432144371f10bf593f7adf64980394f68337f733e6ebeb5d6e7969b559082595d773f01e36d9239b9a286775c06ee8bc2e33aafa2e9bff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88c740d506863d3cf8c10129f6fc7500d14049bdf0da8ede13c7a35a4ca42dbc8362b6d33e5829c97b1b700bf00b3f622c6b8c0ef452c4d45a0e681c28bd40e19e56b39a1e12eb40d27a44c8aa2c6b403c98cb6a21bad9c310b6ce6bdbfd54886cf55ba3fde75a1457;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2451ce48c35290a3ade49e5555f2bab90d75c5799c9059be3a810bb32e3b1754dfbe5d4388abdcdaa5351271cf94d80ed55f291a8edcc19b4ea9c4535da04213011ba27578a48806755d37beea61cf74da89bd397b55a7f426a90c116d516ca875bcd8f8bf4577f803;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd62e3fb1076ce4a2693225d836f0fda7fb0060c2f134779b92dba61c676843aa56957f492dcb73ed3cfb9756cf3ef1d6989c24264a23badcdbbe4264672191755baad5af744004b8a3ac67c572fa0e6ec5d76c871f3c75b03514c3301df8227d39668ccad398d1ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f77bd8df0ed74bb2879becad5c20df1b08921ff869e597f1e182e18a6e1f4818ea18ec9c077619e6d3c194cff089d9b9d51b370a3c4555ff74b5a370f1f5e0728f719ac142c3607be9087c8ae4b59c4c6a62123d50de1410ed2431a1ce58cd65716dc6ccceb69971c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a3a48495db25d193d1e41a95a7c3d233364fc4beb95196c548e0c1dba67d36d048ebad3e2cdd94f8a7cc39b241a4232cc0b1201b7bd578e0c210a1f6f206bac72788ebc8d1bf5b8ad0e0005c98b849266241320eb3f736c3907ad6e85cfbd71a8e90db3978c0f0760;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114b23ebe68a097065b0db9ead743700db2f13538529af6e5ab72352a161a31961e00b622c059ead299a6c22f5ba7ede6fa59e18c01e3884c0f259f1cc11d97de3267a8cf28346fa7d7018a788e99ea0e552bbbd5292b37b08d2037bd38b159caa0e8d0813c22a7e046;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ebf66d1cacfac6f0a9a3c9b0d12ea643a7f258116eb8facb3c3be71665974c8cb3addfce2b260a8d34daec8803163042d344a5f3a5b3c311e777da42f619c120c3ed76f9c5f21774c821882c99f63c0b0f140bc7a66ad7e3e2fac300f9f565efa1ee5236ff62c4e56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8ec4828ab56092514264f35999c64ec780ac1fd42d17dc42010d90f4cade89e04e78cd163f9489a40659accf293545df048419edb1fa799b99b75bb60e9479dfafdd3767148b4b88b8ace78db17b6b313f14c113dc7a16b18ebee6dc03a1addce14260f64df5d073e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116429685f53b7e620d1c2d23fe15d58ee7a0c5050658e91c4e354db661dd4e581db4e85bcfc65bf5caecf065e9461c316c8dbfbf9f68e7586b9b21e2ddce7ddf49ddf6ff8b1c28b690461c47f55c7f734c7b9ae79c47f6e7fa80ec134158ca14bb67b2437b50cc8e0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfac3926fbda21ba53ffa1c95e88735d9d5bf2f630f50262ba79e079e0d8cfb3a40f0b53ce3d65354a675efa69b929d2865e1c6690c50c63db0e03e08a0859b8390e9f6bb45020ce68d37ec5ec3b1ffb855fe123789688d1ff859071339eeedc936f9725769bc034869;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c64d05c2acf2dbda565d71a050c51fa5f507b6ff002a452083b5795c96f4eebce94467f5d24cfe9b8a9cffbba0b96e901ffbfa2ed38f3eedddf6f7f8452e5f89c2eff7464d89e478f61744ce92240f342c44fd08e68d947c4304be0a127b53e7b2557705d6f607795;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141cd2f91e20b55a531351f251e2fed7e41ef4253c94bc0ab851cd4917a79aef42b20db2f9afae2f669bb51fa38e7f340ff99f86afdcfcfb7ca52d176879ad9385fa499b4cca32a0297a3a33761c20ecfee2c538e73b564813021f2efae5a7be2b51d47b9c005620940;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e91ebe5ca6a21bdd757062cabb8e8b27702073085c1678722f1327996972ee041a3cc03363ff55e360ff20f798d41bdd68017949cdbceefca8a4b13f5dcab11a2e6644e5ba349dea5ab802812549aba7feea444f8e71fe4e3cab2feb55640c1fd489aff08d7d9821c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a58d9b4c79ee184858cb2bcdedeebbac3b6431c2705ea1bc586ceefb40d1ab2645f8f2c553138ed033b9c41eff34c33ae3626306fd97550d88f4235339db4e41b949046020bde4d30ba3f978253b05cdf1c75b1474e6e01241e18812e76a0b7c6a69b45f2aa0a3958;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e23caca3010d91f1aa369dc8f40b0e06e492bb317a4321e17231a5933863dc4c3242c1adaa4897b71334dd782326a5615c1fc36402b798dfb549d00800fbb0b18e90a7bc1dc2133a044a1b15b17b190a6da64fd532a8f12b76930b7eef323473cf1817ef5a614f9c85;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96e28d5b7c62ed7343f6058dc79c919c978f000dfe68730e3fcbdb11cac6f5981721e76b468837055eeac6e5c4380377b25bdebffa10cde516f2b531b2e482a5a1938de025c0907fe5d1976665554691754336425a8b8e5b63bb787680bb39d3ba47cad3866737ef68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haef03e93b3071c881d7ce14216c3984afcb6444b39d51095a40b2de4980abdba79525ff6635c12a836f6893ca81357b764c7d9011bcc6daedefeff79d25f6da54ebf90dccfa09bb8c34e85de79ea040356e3acc1a6690588770157530f7d3cb80327b9e888541931b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c5e1118c3c055c7170b764b968c38d3090e0bb3b35719caf45bbc72d567c684828623566e8e1759aedd13e4d7535e7f6780bff28337488affd312f6e3a4aaf79e5624824c39781ed58557f190321d108627707f36655f3a4cc34ec2a21e03e3dfe3fda56de47844b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h887f526b33216e1b0088009c21a3f6d9203b159d17410161e3c22e252795b26bc7d2dd088ebd696d32bb839ffc3155aed4bcf4a4edd10d87fafe27ca00b8be20b8a688202dd9b6479aaaefc9a9f30e650c76c99afdc2b8ab7d627626d0c7cde284e8b050f60efa4a0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf44627a5aecd4995d75484952e9fc3c31710644cc98e69c549a7bb32020d2bf6ad07fe998d48662aae780c6e28bb7a4b42c95e0cb09041808deb429bc414ec52c815e264f82a7f0b5f17c9ed8e2930441bfdec0581b129b140dbc1aa351bbef3baefcd141bf2b7149;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157519ad91c379ab91855f169103dd79bbfe414e56272b28f6f25114eeb1496047bcb59ae6e3037fcbb0eeca3ef4660a3057f231065604ae811e8bda37159cc1bd6811a44c3381cb9df1620d509af049742c8fbe699384b313336e2d2008fd9587312c673b5557069e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a57ac6d2d2e27723fb5d36df4f788c1b36c446af1a748d6040b17778a4fc7b9a0d47dcb1acc2121c3e0afbabd6748490c96fa7b119603a331a0f1ba2b8f7194b2e6a2c8e58d351d9305708a3600fad91ae449881c148cfa6e2301764c896889af1b54d0f2854457a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee8c47e8cdaf2d2f3af0f87e163f5a3942f4b9997d02d62719c4acdb76a3b08801f2b4f3da81d45f97fad13b2e321d10aabf2f564da4bb23884c6ed8c1fa8ea0f9e9d28f0555b89a429031c251f48ffc04907945df37c57fc44d002e1b9a8a9e7867153f1b4ba9701d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1591ce7ca968d8485b68107c13b6456197129bc3c4ae34e324a3b64ea5fc91bab6b8ae3da0d68938edcb8f12393b0af5a5abd84343ca2c8e6ca139a3512fd8bc0a8c11e19e5e86a1e53269a13cb7292620318498794b6bde8c0eb5002cdcac489f429f468ad6effc0ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he23fef8e1f547f75076b11ea95eeafa26aa6dfb7986d776fc9ef2c7c48430214ee7f4f119db0dd572753ab4cb8b9fe968cfa0f83fee5617267e5693df68cc6d5b2d0dadc35877bad4f613074ef7e10b51af099a37c6e9397a366614494b893fd50273c9fcccd77bf37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f77a5990503ce4034bde17e8cc244ce0823f0d400af9e4f6592a5e8a16473d3cfb5485ea5c36fb9b4f103901027af5153dca17a2101ccf69b5257608f4d233f2940ab8b80ad406515506fb92fabb1a474b47e97d0556be280b0ed736cfb64ffd1de66969ba4c0c1f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f742fdfae3d93d42e5db2bdfbbf4a1141b40d775ba106f63e95859ad9f6791f8c15250b4caae9f2ab707b7e8464efece07f70bfa48da1049fe2b6b688edd6ff0e5c49acd0f66362c3bccfaca0f6d3a810a6181d295274817e2437ed456ae4ee9834de8dcab6c29e1bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f223df878e588ef29fa8f99c6e8f3a7738b54e32fd4906b9180d7306196eb201652661f82b969efab248627b7c88c5e13e92a6bf9db7a67bcf4cd52a89e6d060ad2c98487af39381658ef6f0477e0791c07a17216017d5e04f39af3b64bd5d77ddf24b48250737509e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e91e7ba0318b76ae6cd17e3f7f7cf65b3f91b2aea6a34dd182cdf15519ada0d73bb2bbbf8e33e6ea8e4186a0678bc7e13810d034b900ce619eba219b02de538b4451f60f5bdff8a9b4e76d583a1ed77d3b6c825e04ad818bdf5bc3860281fce53d2df7b893b58f93c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189a2f6e065841a8b1929ed7d16dd11df25e6de6136d49a7a01313bfcd245271538d1a2620412893b0370fa271c0f6bfec5aff7ee6160ead5fccd7cb02dd86dd2ef2466b35ce116b85e18b1a18a5c31c448d201ad9ac4428ab1279b7dbc420003a3afa1bd469b68910c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1844caa3802c279853022e3450b7cdc1472d6d2770e945272996413b990bd18ef3dd929d8591ce0db23de937ef2bad34a53ae169dc4ca1064a91b9acaa0fa7fd6e4e266b7e3cf60bee1860e7f2e7f49b81e9ba3956ebff1bd99df81a6ceabbcc533781183ba03e35e92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134a21d6a69e78f3a89fa12e134cb34a5993214bb121b604e2db0bcceef85a926b289d44a4b099fd7b8459e4095e8c32bd1c4e28fefa17320d4bef4c253eb4101a39b9783286c87d35f51bb0ab417fc8abae2d76ace2d100ffa7f9a6f63b773015b918a4c186b4d81bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2077966d88ac392cac068b84c9c3d3f2f2780493b02240a366cc7cc9b8e8cbf3e304ea120994bb19d3790308ff024f1288a5a1bbff322d1bd5dc4db2b47d440800e2a5217921b4868dddadf5eb71fee6b3ef40432b7358b7b60c8c49226144c9a6ef325caddedb444f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8b8eda47213ea0b2467519f9e474d69e262f33c0863b6c6afea7a9f8f717fb35d6df2e4f07604e5944963d3c7e1a45449d7d8cabbc43b5b73dbff87c998e2c7e4ce2931347c65e2020adf01acffaf04541ae6397e54caf92ae6e4f92eae24043af19a0a56f663dd3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19130508c80e0ad93f0ad8a19cad20feeca9711a66010c8c3f24570b30bde5c52592b76e9a1aa22ce283a44f15a449ad34372b22edf2b448bda7681d48590825d4647aa6cb0c8dc3a0d1f530a1cd2c99bbc5619653dacf368aef1662cd9adfd9ac4cc27b91eac06d0c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195fb146fe738c207d781b20ab1fd7dbd21189eb110625007073bf87fffc9f3b6ef222214db614dd3787397dfaa7cc1105641e7b3e9b1ae35a00315cb42a3987ae415ec8801c657ae8923a1f29d55cd2c736e086a0ac99771cbd02da949500d08da5447a69b33e012f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf96814c4a7c7a8e0c667a2a993e3929e9c1e61367f951cce83667fc908876264cc01068061b08f41a55eb1dd482a54c4e4fc3e4761d7dbf87d981f68e22be7deca5d78ff694d3e9c40909e185952ba02a17165d9c5a4750039861854572375e32e08ab53eef21ab7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19323f501deb03e601dd3422d3c5c8acbbdc45db9a96784c5a4e1267a2badd3e58826c7d5ed522d74ba95c63ab3645153dffc888fa6699065e887a35f54e704d94409d7c285a326eda84e5e10400e6eef1d43f9bdc2f2a6df9e886a3c0680493edc34468ace3925a94e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h940816c61efcdefaec9413abbbd84c1c7509be0a51767049f878c1673c77606b3cd64cadb7b0aefe0cf342feaae97409acec1b7c45b081ea2ab9c2104951260ae5c4f2634035692eae5ec5d8d2866120146deb10626948949fde8b3b8be07d5376baa828e668ec2259;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h805f860b493d25400d700e3db44ad3bafb19352829f1013c188ee1befd5233b586a1176cd68c1b7addba9a11afc770b4e5d25e43bc02a463423b7b8ae2bf4c84e2d759b2a926268388f952cc97cd96a7293ba40e33f76cc56f6b56cbbd843d038461ee613352cbef52;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h887855c611c355c01428873834f5b4d5a46eaa912ed0ce8104df2f5ea126bb0eacd163f6e4b21adc7ab998b827fb6c0cc8de37a2a1a5d63ee7035f8fb90ef8c1fdc152af60e053c0aad066a1a830ebea562c6201a2d6e5b277353dca8cf1bf9a4dcf1ee2c827d76855;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b20b4e8802bc37567f87318d307cc935693c40850acb60a1c2acd13bb9b7eae5d496b4ce2c878e92f4a127c786da0ffee18f02a2af1f3ef363e08f4aad0372bbeeb022d878986da3a2356e6eaf8c4744529f2dca32482773d548dfb9b575abceea0fd78617fee2af0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f5d7b8dc0fe06304f79bdf357d94de1c696502a892156f3dc5782a36d6890a8bb2896fe3d38f0e98d426f8bcec9d1febb32dced66763c85b732319da4cf00b98982760bc61fe855dd6510465bb2753426240b0291641faede9570ef69af909b5395e2064846706445;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a93dd4d858c9050b9e25ef0833e258adc1bd41a49e693276347213a09e1e79e3aea9131aa863854d3a8096e1750006527ec49ad2e0acadbf9e4e6557d28bfc5c1816975ee56091841887dc92c5beae479864b00c8fbee4990b4e49f76e95f33948282aaef8821d338c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16cfbf3164cb8ec98f030d266862ed3dacd4f2c42394456dd2af38ee7de3d25908e91c133c7cddf2c294e15719b7fa623f98ccd42b3e4a0dd5bdabae385e39f58e117b88d915288afc211e7a2caf64a3b51d0d584e3dcd2f8102ebee499f97136f318f0f6d7426ab8cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3cedef063ba974510fc8703da55691d97786df6cd7ed08b4702a4f05eb2e6e61103b648281900c9483c62acd7408a471e618e9b120bb6556408f274702decc339c143f55d6925d5808ba1a56846bab8ea66bed33c7cf47c4acbaa0f661da523191e059058f4262836;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f10a971b184df3ae1a9989b7ac5cca20e516fe6468c28208cf568383f695094d16ea891227ef7248ef4de33fa5f0c3c314525af6bbc75c0b4918829e50eb2cf979d3385edecd126c12989f5b3f5b1efecdbd73407791ec63bb163cebf3847db45a0bb899406482800f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75466e795e08869bbf02e45916a93f37372abced0606496a252785c7f5242583740bc101ceae2643f1fb7a0f93152e6a85c4b85ab1e3dec821014eb742a8e8b869f4ebaddccbf189f6171077c97c7c7a75e401fefc799a9b66ae4066fee57f9f722596d7ea203b634c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c00235b401570e8ba8d2952ddbd59c7011be9b3d2bd9d12b47d62d9e64150fc27966ec799e5db566043d3f22d52647fe81f68e81aa8be29ee0a3c45be01e1aee392b465a17c5a8f286d00e17fd661e5f73187a68b4a92472d33b661296c7cd96097edc524e737d3872;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2605f55be3cf7e04811224c2b03d3a2c4198f8502bd0676735d94ce4b76fd3b173064ccde8db9a63c48b6a2b7837127a5691be067950aa7e65166e62535db9665f629f69ff2e07b116ff552efad9b7be8b4bed5712663e4cec18d5b5386243a86f940e08f21fd3a70;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cccea77c25acffe5c099e3c253b0a0b32d3100e86ff1c22a4326e04bf65ff2bad833a3590f290cf4501703ed4e9122e640c1aa1dc811f89ab7c7c535955b5ce029aba921e97e40f8071c3944d22716b18ad27b288fc3b0ab9d41cc59011af85639412b9877ae24e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13abb59a44adfae618beefb6a065249ce89dc433986c995cba555f738f60811af234aacb22e7a126a93e6f34e214960a8656224ed25dca99929b54bedbd01a526234c1d04dde90f7db0ba04577104bcba1460b827734b6ebfe10a7c420560736a4809a7cdb9ce20a23d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h446500b9be08f62b6f8c2a8102a29cf227ba7e0ba4deb4d6e34b2c87326b8bed8d43b05c669c7ccf3ffe13749556f8659d9c6c603c9abe7d06d2babf29513c01910e2e5c93bcc370aedcb361ad4740981c84a1c240f59bf2482e341c92b69101c91300053a11edb34f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128e8f3839b058b417051ada5e6480a15f53e677d19b6eab8e447b98f107356c6a6597a109b3aa32374c5496d498cefb09852b061511eef3835b3eedb05cec7861f66c985eb61629e46dc618bbda78bc92705e3d6b49dbfc3de59d9f668a644134d758b9f6ac480e474;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5e0294e0032cd4e4faf17fb8574a502c7d095874820dfafda33cceef85938a7f344821cd2043bf633ff51383d39cf8279cc443d171233ef0bc02e8736d98a0d3b0f1f3fc3ff87526e7acda047e39fded9dca807e31fdbf373203283145ffc955bb8ae69beffab130e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95f56defc032e9edbae5a045ccf4bb731f1f0d6bae1e07f7ce7eafccaf1666234c52becc3de76474e8e408df8c4a93986d37f709ac40689ba29319951b81a3ad7820de47ca9b26628ad4db64b3ab0a766ac2315c2dc83129bc00e279ec82320392451f2dbccf6e9580;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3cb3e8c90d207b21188ede79b64902f2fee710a0d1b24dd9b559769d67850d1d1bd5cbeabfe5aaf692ba46876fbe5a023b9d299e15616b6fa97090ad46d2bdbce63a4d7c77bea8e039cb32261d33d7f43230905847d34042b74b71c7f150f6d26df676605b4736dd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb176c5fd95ba53bbf0122e5f6e61bc8aa5ba2ecb796e1b53e16b77371963b8f34343c975e249729407bf578306b27c4a01628c1f7694ebbabff1bef4cac8ab7970af12a2166b9965510468a0c8e5e0fc7a085fa3913ba8d28a95ebcbdb125123a72b8980aa14dcc4d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h318b94ddb488700215ed17bb1806eb06dde348562b0e67200b1029b97d9988b403f36a4c25e3a2fe813c714bb0b1848023b4cea04a70bdd86de90e67a06518f5d23529e5b8a1aac380cd4e60e4691b045baef0755d1c6b56425c137555a14ab38704ee093256e87da9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76a11454b43a58ce47642dfdf0b96428171a28530388dbc1a9e5c47a4cba21bbe1f336c1667d3a43b3fa0646b96778bc57217a0c490f26761ba8f528d9d72cd20541c17228f04342e7fdc28ea060092255bec3556df8eac89f4163cc037938675c11eac3939d2166cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbd3a7cd744f33c8902f07daa3a65da1b1e23a0565109422546c2243558f00049694c8e74ac32f214b974bf6136004f394c9c23941ea5cc7d0fab752b8b9449f654e51892af29adb765a99c5dec97b8057e30f5964514d28973e1a9827a84841ebe19d0348c01d22a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebd81087677faf6621ef97847836c931a4b9bdc05b78e70d73bd9fc076642b336cf37cf1d9c026f6cd3e9481f618838ef811fb6f5bab5d4da262378cd0b8ab61adfe73798da65775bfb6c002e929e24f59f67936127fcb472d99d72eff1a1e42e36df2bacc6ad66a23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cf4ad9f6933511785c7aad9edf77e799a8fb2beb38069169b51ce3ac69b334d9c11b3eaa90c47078018241cf630c51551ebb23121ef1b322b7239f74e6f97260d3012f2a3f92f89869aae89e5fec913a47b2b2b96951787743bc2e1ab6945d00ec085bbc400cceb2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b0d001e847f85df6229673ec7c60c68b37972cb4bc1789023d20eef69b862145997b18fc98f0662fcbbc492e18437bace9f73910b45a38a4f56e210ef4340014079563c43eb187b651f9e4706d096435f3513357ee2c94d0ef303a9590a3630400806b85d86484c3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32eecdcf3eb036655aacc520bef3de1f348ebed2ddbd7a1a3891f95c4cfbcef3332c86f0be5fff7df3939d9811911148c21d31af14fd9652aa933fdb8f186256d2e77d6d8e395ccef19c770ef4364271a9ee98ee599334a8295e4203d312c4d50348c49b30d24158ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb83262a1d7a333aa3fb2921fdd6b56bbeea4ad75669966f30ea6d1844b61c57ead12eb41faaec3ee7a27d1e21512299fbac07763a825511ee36e31c6a770dafc8f09c12a8de6f0de5d27f7f1ba3165efbb93c3362f816e5539547bc0895753da1a4e6233d17ffd34a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f50a96ae1a59a3dbf5b703d98db51bbf134d45d1643818056cd4735f99a5262d17324c2bfa29b6e8bdea6dd356e22e9800da43f4c9c582670cd2be145e7e1847f51be12c332cc7bf899f9416bb4939cb1f04451fa61b6f45dca4807767beb0bbf4ad1793a56f499b78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2dec30e0d23d986cf605e3866f3b057f25e2ab02b431d93a2545d137364fc78913eb7d555d1b70715ef4a472316b5134fdbf63aac973be5d2cbd03077927886ffdbf6b0ad54959270d4e382819f2a3597b19d169656006e98447598864e45968530ee6a680c7db310;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1570b360cffc261b00d75969bfe554ce23de579ac34861b0c42d6becaab37853d3e7913b5dcb8771b2c15781107c77f221113c44300196dda7fef14aa63a56803e32b7ced7578cf155427082d36740f9fef32a6dd06296bcae4cc2f9ea570b461db75d453370f457d33;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d35628a2cbf1af06aca7f29335ed7d2df4c77295e4d607608f182e013c31efc33bf115dc79e419262f7fe54f59c1f286cc54631ed7bd6d5e4fc7c0a305239fbe5e9c1b612ee275b52288883adf28042a5b02aa72afcfa443d4005fabdd6d04c09aa22366622f0b4f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf17cb4e041b0d448f344aea6e8e7db7a34ca074e654b54af9f01cad5e0dadf257c6576c91b7bfd82ccb53825b162e558e573b10fcc4f33f0c127c9291a0b6a8a6fcdd6a39c5e4afa23c9a2b94fe215d79b4295d32698b09b0a6f59840bcb055552a3018d7abdc5c029;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd14b8ea5fa0defa386977f3ef3251696357de78fb33cae60a4a7f28d68efa6fbbd0647d16534c6210f9a6b0b28ab8b2dfb8c9e1e6856f2578b242a896c5b78b96b28fe82e971bc26ba98f56333096a33761e223aad0964f66ab50247a85249093eadbdac670bde8ac8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd574018eaf1549e97896725d5ff6d8d44bda6162745918af6e496f6582f5421fc33c3b7fc852af0377279c3987181ccf6c0cee68caed4d5eb83e0d454a5e85b39a6f396dc307326c77fdcae5c0a72dc17a76bec91fd390a20bdc421782f20fe97655c5026a1fd1f21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc73f0d408e96937b19e1efd9b1a4225ae046c7380edc38f31b9e0e9eda37881a430d4c00c363cf7af8c59d34e45115c8fba08fe8f71a9756b1cf16860ae2a7eb12fed1fe3a9e64424e5776256e28e4c7d40c5f00b8fbb7a1264a592c628a6bb3ad0cae9d95b89980b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fac06ff9ea3bf5051ef12950865db70392aed40dea9ac144c040137165253a9588c318b3bd383453e8574523534ee782f1c7161ec39d54af9760ed65a6ec9ab3b8538df4df26e8863ec53cbfe6723ecc357330106f3731c51e6abbc6e0f00cc0908bde697fccaaefa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee079493e068462046953f94e8a435732e86758ced254bb96fc90fb03f8f71bbde1842354f02a07072abb8448ec391e5f8874c572df2dfdab7d2805b12cbf8f7dd3679a08c955c9e5793b21f571de3e0b712d87eb7716b3bb5318d86a22cd8fe69357b1b709730a7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde6f4d54dba2934c3301b75ac78aa9c2c61d5b1b39215592a02f6043ff5fdd2edd7a7ff1debe736cfd2277cc64ac2e5760363975dd2e7e1116e3f751728ce10c1cfa238570a27e12493f9db2f0210e24e1581a5a01564a092e6e38836b4568f0fefc313fa84d21681d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf320eb555df444d12cc462611c6c6c235120362f0f5fd20c9322e72308823d754e0610148e9be26f701f1f0e8648d3df197ad0989a53e8441bc1dadb1c54edb2022d54461b890d43cf453a896172649cd82c77906d2a079151d834fb5604e8f4f141ccd1373659b0af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb230dc6aad00c060398306180cb68eea7b8ac8da93ae6815459c85e5e5058247b391ae9bbb4bc799491dabc84234054ea4f18895784d406aa79e7a4f3b304f2d766c11c602c96fcec4b63cf8abbd67443e125e4749b05f1d5f265a6ad4f672efca6a02f6905883627;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e8a37badbad7ab143395463edf057eb5f66f1113771af6bf120458f4d34146a0057b2ea9517948334215811355a9622c1a19c73cd50151f5347115ac8884c47500ec2bde67a1c5423db287626035f8d59b0fe5ced69979bd67893b8a6ba694846788a93077f44b629;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8ebbae009bc5710752fa8d73b16fe00f261e9e8dbc2c77a9a00a8055faaa2c22a00fbaed64b0d5d7f2eace555d77b794ceb01903275165c8211d8f8a3c9f59b9d2ab2cd207975d3a2f2f08040fba7f858af746ed1aa35ae1f892427992af8f3583481f814c641528e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa40825f948acdb8e89d5abf87a893a0966629f2c49c4e2c3faafe1306017e8181b3d37534a6d6ca4a4fc3d708f42b3e1304ebf52d813380dd8cd827d7bb5c6d29fb4561564fc032e8519232c82a692aeb65e73d3fae88fe6930e1b54cbe48cf7dd7c9353105dcc985;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h510e97cac0051ecbaeb5761206663d4b7fb1e8739c2db843d01998f2473b48b7076e264889342d1c6cdbf029b1a5a6494f7015f5af1ed066d55f4da63917b8c601d921357bbc0ad5f757b98dcf11503c93c757913f04477ea2e7d549e189769b6af6908f6deb5a2470;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6515de9a9cb33a1954682f54665e358c802ff800febb1ae868d4031c98e165b0ea773b32a3dfc0a71659ff2fb3061526d6bb0e5fdffb509360d3c8f0b94f64ec0374c38b6b18add2bf7cb570ff47603d6b9201d91dff66692e7a187daf7be089e887dcd66047dae601;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5e16a42d6eb4377fa0f7b2f58ab2a27dc7d5048893b6fa4588f1d3acd9a5bbc25ae4582d3bb72bf44876ba32e63dde7c4a6a907c2d5db9e02cce145bdfdf508341a432a83a8ac8c857224d48a2c18448fdc52f8b8760a68edb0c2671d6a5483051e981d2a3c1fe77d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f79c794d7e160ebb9797ef62446d975a1dec24516ac5271a92211bc7b106c5beb56226a700d027a4939f35683552eb9bc30cd4f2d7088149df2b58c0e40a12442a02e7305bbbccff83da899e066a0e246d4aed6a823753a93c7d83e24766b41f4c6efccb594bf48ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b22391e8a7793b6359d4548d6b9fe304113b01e5c3f4c57d929b98b9db689e13c380fedaf9ac924811e71a46563f03d2de9c34951de51f2e93a17bb7bfeef870cf1d82784cef159724db02946f56ff4c102664ba42e12670df5c5c1e87305016378c0709b70ac5d0ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63155ac1101d7d410670f465dcda85ba8f10b1ccc015851894e02856300d1e0e593b97155a37c0290b6869a48fae7a99e577140ec1c8f44af928a8c00aedff97c9ad7622cd73f09919fb886e156cb20d9306bb38e3b8b5847e2955f561e8b5bb1ce82432a694a0e2a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d663df5fe002c7a3fc6601c5d634073b42ddd2563425086dd98e7897d06c3b081a0feed1bbfe9ef19bd93d6acf772b569aa7857a059c6f0625a8ef1ee448786b4de9bbc33912c348e1023dbb9feac4800d32a7404bb67d7fe11965d932b16e73fe66f3ad2800e86d16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48133de49b92567f1128b209e7139de97c25b7b2116f4a4e437a815784848929496cb158a65c1f4b40f28b9c4a78a7bb57978d099e7e9b4b32c7af83cd2b9435423ea0acb39f04e0f9c0396fbd81152c90f8242e67794ac489d8be313b27bc220cb64f62e1082b7939;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1943922a82800cd5267edf48790e67095ba9aa166497325090802af3eb62105678fb5dba4173a7fd86d4c0da276fc16f5bab183b453e9ab4eb044c40688ed03da0580333309b0b09b11871f2a503a861f22f72bdedfd3edd5c143d378385dc1b4295be14de513cef76e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc961d3a97de6eb013dabb32d19fa1784579ab68cb301ccd1f36df4c6212805e243842ea4aee60e422235102ce2874ba52ea20c83374f78e934700ea11b39c7f512136159267db3e052a3760b1bf51150fe657b6e1e24505d04b9ac593d4c9da132a36dbcce58c05913;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169c4ac4d3b19006a4b92d6644648c62fb9346c0b6539ffdbfd9bdc3d63e80c2d3050d735b72f8eeb504763bc76fee112ef1256e85ff87c4489107d2455c4e90d75066a4633466a3240ab18fecb6fdbbacffe4a997f72574319924026860a3ccf218fe456db40a33831;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9d65a9ae7ed1e02e102fc5871f4ef1ee788891a2e2fdd7782c0bd123bf82244b944ab0bfb8f3b8e113ae2e1f05fd6405a5a96ec6dde3a10697be2389d80227d7dd5cc77438b0e7d34cc8f673b9ea578961ec12f12b7f6dc2eeee74c80adccb727daa5a78181d241b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h577821259457df7c66a84a696ba807151a97613672355ef433aeaf94b199810c3779528a751aecfda2d4ff77d43c4881e0220d2fe121528eb2dbcc1efddefdd86ddc9b342c82a5016ccdd30077c16e39635f863f4a11daf5f389826e043fafb8a132b711b0dfecec9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c1d6e1b64ad0833a9d04fb2b7f03c472d91ba234a20bf269648585edf83aff693081dbfde30427218d34eddf085d70c052a1644b05c1160334403b803847ff253b5bfeff34a137af817517426b1aa4c0c8061804648117031955881c5363e39f4fc11bc56fd0f16ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he610b79ec0e14b664c99644058029522a0ef491577bef54f94305716316cec972c5ad449ae0d21301d36414c2ab80075a7138e4e6ad2cec0d4490f74d9438fdd042194e7a53186520069ac4fb740535418ab9f471dcb130091b23593a3d959063a7d552100306281b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3870cf7a7b30f33f97ed5014cb429d6a75fba0c4f4a1ec7e0ee715f2065acbfcefa876650bbdd904a08973538e95f6909b8b9af537bf229e9fad668903ab544a3198af3b8aaaf331ce4909e4f6f2398af7950a52f375e64130cb9c0b364e50d9e4a075e2c59b0939fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h597400f74232b33110a301735055b63b90ca28338cc544a41dd61e01146dc8f385fe55eca71d474a070d59ba51854cb51c805e2f0474002e8f917e4abb5b026767a7ebb3300ca23c11a13a9d66aec3e985f21cb611802425ed9d5bdd9c166a5cabd2224b9db00c9474;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha87ca66fb7897dfa43923894261adeb232eb4b7e7be97f84b57ced914c665ccff28c72f47c18b1044e76f31346a5bd1727ada76abf9483068ddcee8ff929966ff1298e7d3e973de9497ffbc27645f34f91c826639fdb5aa920954b6502b1e679b8424c6006242754fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96b0a22a4f63a3f370e7aab9965c55c6c53efd6be1dd0a7ab761966b41f8bef9eb95a29b1716594dbd76b1b82edf1df4f5db1d20c6fa639ec72d74e64e3feb561602c44c97186545fa9df60977e8c4c16f782be536599a845b49ea82a56d806307849a42e84d71072;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4893e1d9a27aed9d5f7b86032f0d3652177b1a1917240d3a06e91ebc1c963570728525ea659451cf52859f674beee2be23d0ab0546ead74ef527a76fe20b6c3ff229b22c909325cc424149e165247161e1c6046b6799ca8a6f9a189983a7409bccb255c64ca701c83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e8ff93f6fbfdd3aed11ae483c0bbdbed5094775f8507d3db86c462cc9ad5fa9727dff2bc06ed4cb991424d7857f93fb6ee3889a5b85ea4b84ec7d8b3b00f591a7f315382d8f8a610c97f5ab0a9c5e29a55354d5572a0078862734d7873fa53aeca46940381ba70226;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1454f34304976049573d4898d6bc0a8562ad44d63cec9d29b4c005319febd76ff624252c53d0454de07d05f441c60fae45cbebb0556932c0190d9d0932d3b22be66bbbc9b873bd2009c7751a0f3f35a9754fdc56bbb837260eb30b6ede1012b3e2788275dd857186da3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129f43ebf2fbb2eccc68063b847bcf9e5e4579cb82e129624ddd9564c8bc41c6714f132a182af821174d582b99578fc767f62e20bb13b6a0c5e72469d3370b664d1808d2608e21dd17141e2010e2e368a1e9023b03fb60052f6619e3cee2b767a9896bd03a54f3abf53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9be68236c635696b5bd68a508c656ac13a146e46b962360121401d60747ccadfaccca3925714b7b259ad3e1e1dfe8a04c60804806c0ae05f89f4c9db3287d1a3725a2e0a595faf0f6fb11aedac108ff8f134bce67a94d101d7185854b9b2a9c3daee0e1b1f4079fe3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1237ce13d2079d380767a6b373e8bc7412fcab37bcbd6f3f09ff99d1e0c29226e85270ec449a3d580f631fb2977967b900c86bf5f6c810e1b02e49b33f46ef358d366315587d248dafb7ad84f7a5171dfbfd37eab73a6ad62236b2ccd354e9fa39e005e20f1e6eeab8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0c57edf52abc7a023f014a95065fe2f02041032b87abfbfbd7061329f4807c250f17e1d55733c5de406b45a14b786c7c5ef501cce384482d7459bed76d5f3170f913c402fba52db214aad9b1df755c1adcc6fd61daf705a4788ae96fe8eb493116fc0b2654b214dde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dbd98a072bcde6508e0a7076be3a0721ed40c2d4afd941cc02994835e4fafac34e872510f7dd382bcb64e9bc901c4625464a5327729ae066738cd182baff79743fa4bd9ad761c8252d2ea9c795ffbe6c8fcbfe957d0e572968b319f65b49f1c4920e9780771121ece;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef669e808d71d3367c32eea1880f512fe211ddbba03929436e18c68c79011efcdf77ce7639dac08a229d7e203f7d7bf276a3d093c3794aff2f0b54a8ea39007f616b92f3ed52010845f57d87dfb7ae28c6427ee69b2470256564d78fac4c2695b2bc1ff9b0162208ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bde3cb2dd8ce70306ac23a82a8c7b8bfb5a9f9cc2776de0d9bdc94f166905882ea634780348ed2e5988f396b7358af12c8d7b4938090ad45c737045214b06a97fb6bd439ea175762f2ac37163b0bf6f0d4e3e4456d6ce3c9a4e8870479f57dd5622ce9b966e2391e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acd83706f63204bf7212d7550b2c75e7600d119c2cd529cb5a1c69049efa6f1e563135d8613b4130d84b300c487b1e77d11b3eda3060ca7512bae5450bf32e5e726f9bdb989e999eb9915b2c27b82b8e750920bce14a7120217dbe01f57c7c585968b38f0d27251824;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14dba314c6bcbfdae73964a42118d994fa4d5fd7567959c0ad15a365a1f85dae8430c78fba23e3b8a80b7f7a1b446175d60b8901e8a73c5b319b45af3a4a84847da544cc4006ba0547a3debaf50e97a737053bc5db7763c38e8fcc5656770ac09d081123d05ffea5c4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175bb6fffbd0d4ad4b59fb931400940f7cb5e4bdabadd85fc592e0f13312e57c3a1625efa8cd4adc83cdf0bf78c5e4bbab5c1dd547a217f8567c33aa5f7ae0110fdbda09f30a7528f6a86adb27273feabefe4d7f7e73f24f4b385ee4f20126b1f3c92b6fd19b7a17d68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0ab62fbecddb089e3f2e8dbff03406c097f3938fa96e5462e8a8e58d9655b9233444902ea90d089c7160c6c14f4c1b262282ea6f8073f82a23e6059ed1ad6f8fe31ad1a7b274637b97756c6016f00ab6d61a4613b92e3c6d148433ae9f7032024a81fb415cbdf0416;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h619fc4ce1b21682ef40c9e49bb3ffcc5e4ca2553dd3b7954272f9a532de6b6c9edbdf0abbab4a6c899444b6424463f8efe533c565be2471e08e2286cca1ce28d583504e144a8a456a59f234f83145d4fadaf2dac81c85cf4bde82d6dc828c3ba73a9a86bb24d425f6b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea8359381bd0bd1412b3b0684e48c37e7951844f62da2f488fc95f331d00c81459aaefa54a82c149547b06f9a7038d89949176d6e85afbcd572ea6449e5d3c9ee4593aaaed8321f84016cc343b7ca664ab33e6fe44a7e2af9c3b1f7cae42487756463aae144cabdf3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fce169f24014d385515831913f7cb66d171429c00f2471878595b025df9c84b8161f646bd885a93b4fe6242eeb6d2d4151ea3641a172f7cec8fa2b5c942a00335b4d9ededafdf01553bea54857d8df7b10f700a4aa346a6a44a55bf1a3a3de5917e96fe6db5a942249;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa04aa9ff9b9d801a846aec9f1dbd4dee3ca853e67e2dc066e47c1cc0ac7330f752df65685ffb4b30bb423b430ae461a37c8d4e9b10d8cf14c293e0284087bb86c7709050595d1e302efd9f5f371e3609ef41d2d9ebee18f411f5dd34e2e2cec7b2d99d0b0e0fada2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a0308aed854a9a572c86564a9d3194912f30b445ddaea8e001ce1a137357efb4429338dca53a7dcef289123b849ae0118bc9edbb54c31ba778ad89359dbd6350eafd8c79c190f9c758f09377b3a9742cdf208cf658daf816179f52ba0dc8b389733500baf36fcd3d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124178967f59e470e2b1fa6e2a26c00985875d3ac71b5fe29c846eddc065b084153ead847bc4d6342f22b06f52df0243073e072743b277b8dad58628789665c5a0bd09955802f44058c1637150c2ada903bde294816b6820709477c98c4ce4b403ff0c4874e310ed675;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9364cc5f6948e31a76e62b475b7e8f6ed4fa80487505edb07ee5ec256985c5b5e86eb122fa4c16a4b573df88ab68b35ad5121665b23c20c49f5fa83ed6968a86875f3292418cd22fc6a7d6d90f7aebb589ea54d5c19ab733287fd9b2b471d458b822c0c4dd374b53d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dbf3c430c5c475e9be31746d849de007d587f48b8db472249a3de572c79b77fdcd5ab5ae725180d80464a6e283066ccac5e347715c6117fe0a33a7819d15d4a67b5c533debf776d111b593e8f1277f3fde2a6589271c735747df86104be98e13ec2b2eaeea1e343f58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ca41b54d688de966aeb7638b1dcc564dfb266ca0ef997712d664c36336e650a755b9aec7450a7cabd138645c666ca3e46a706f80af1adf2a8ca1d0c3c7580f7a5ebfddd59f3b2624f5e7b3075fcdbc6f37916e78cf15dd3e7cd01eb0b14a0106ab00bf1962376dc0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b79139f0a8d13caf318ec2572d11052dde6e9dc8d4aea532ee5b4a36b8aafd0bc03b977bf4f82af30cd060f71213f570984527272f725b4616e53a1dc005f6b6b894e0ea597b8db6099c49b11d7b62238808ff1bd0bf88062642056cc5f0d823420141c386da0755f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1888122f3ddca769fdcf69b4bf1d0e490c974a93200b32f12f1728a2f94e7f860a5b743626657f64fa8996b1ba91b557ca72c1c6b34380f68734d7b7e5d6c19e2de934a8a22c91e7c04493f45c2865b737608ed4fb30a4fc0afe1023665f51ca1f4be98d7449cd291;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1a2db64cac3dd69c81d70b80bbaeb7a61ba776a0fa29210748e71ebf5c9bda18e433a2fca6cca66b439339de7b24cf1a20bb3613f6919b46564e235a4a8b3c0f15c7c31826f002aa4b556caec0bb8f1cc629c2dcc4a16841601d81b1f0d9dd878c90ac32e40ce55ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103e2c7f086612639c79c5967a650e876259d7350e53ac722c6868781d42f29e3ee366dafb0aa7c30f16fd87d38e2a4c58179d326491d42ee2bf3fe83755ec56a19ca5da732494d084379d0f9e778a84049e7f31d82c69d01b566edbcd012fadb7ca6cc716e97dc646f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc8a560044ec7bae18a7d584d52064bcdf18910b01b407696f214c0686495a004ffbc86920b33e66309ef2d9af8d40605d4ff7cf1cca6f503b9e199d04fc42962620b081580de0254f082f9d946964ae2852fc3e5d9b3111bef1f619249fd9da84b86d5bc88cb0c011;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc794a91d8f618effe431e4cf5865dc9f95d41dbf1b2c4e159bcc378f381461665404ffe34984d6ec1ef301949f62efba4020b21313d773031633472489b5de9c6ecf20d66c6fdbfaf803b7d67d39aadb11e61d98259f1cb45106937e3d6b2d815f341937aaee732f45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106f8789d4e7fae6c0a9464a5109b25b3974c0bf356640524d9c7801ce6525611bd9665dcdc9b71af8b00471e904208fea9f2d16b7cd46929ed5ade50af035a3f45e317359d3091cfcaac38ef16f9c526edbb8046281f680bf09271abffea997fd5e323c62f5408707d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd90367e2daa0f56dc058a321e3c8bddccde677b05d9b6ec8cd6691fb8195b473e9e2539dd6da10f7569a9266298ad47a6ade97e1e3d9ad9fe6057f21d17bc828afe42a47db8fd2de671f3b5e85b155cb172e939c2f71c69efbaed93ff31cc62a5bf38e995d391096e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf2929350ce869fb9af42530c2b0f2ac54ab0b5c5ca2f5dd4b9773fcf17802623872c2557104879798586ff4ca436ae184c29946c3a2cfa256f12bf11b9e736b6bb6484624c31b8961510066b1c0cb26f33115bd63418e75b2ef346ac5f5723192b9a98eb035ac2a5d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cf32e1e22ac43c0fd137ef9240bc9fdbaf6640d65409d90d184af1dbdfa78cb69fffe4cdf402f11830f5691dd7d7696d0fe520fc2dfddaa9af07f2190c34d35a11e07c906775062f0444409a750091253c24811c9a804914d2e0f59e144b6e3d2a0297f439bdff671;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137a3386852cddb57ea3e5f1b59a2f5a9f9b2861aa1ae174fa3e599bdd3add9e12d18b34d455b698e92aa796a4559cf0b7755887fdc9f8d9d4fb439634bbe103f2daf5550b8385af9914cd1c5c87988cd95a9fe47b4497de2ca9fa07ecfcc47644fe3a1f02a25ef34f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f34274327c6084e3a187e0c2a0b57b61c4cd832a16fb10ed58c1b63ea7a3fd7b529d0aac38d9ec072933377fb92df19130d50801e5f073f770b158588ac03dbafb1749a375a0cee619fa6049b8ba620099c83af6d315e0e6536220bda6c2abc34f660c2159aef2fc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bcfb1423af8261ed79a7166d8929d98bd9e4aa0c891c3f18a9c2c414238ce460d37099ef72a2b2f9690ba611fd4606219d59fdac5c3e0ecab035383203163162f268963cea90d49f7287c5c90460d3a82cbbb16f26f03df5aa9b5b393b32fbd5681a2559cd35b7eaf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1425dc76c48c9cbecaf9c1f3804e324744c2cbaf70fa36a48862923bfec34fab6310763dc50b105bbebf2d111acef4504f5e0031116e8b1ad99d748f62c85312c354cb14507066ac0de8c60298c6b6ef4bfd0f7539280beeb56cc5b56d84cb22d8e1428d2a01fd87e27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e96aaedd670d5bbbf589abe7203d61f36dcd840ab6960f2e855c3fd8e9f3abeb4574c3e8deba9d4742913bc50290b10c4dfc84cc0cc26231d65d838e5edd30e7bd89e38bbc2c3b73eefb57c44d3c64d6e886b7b82844587ea8245a81e9860149775833b9269f66c732;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69d537b6500f389f979d53004460c241dd7492cff83119d1fd9624d71eb13420e49c15698b3c1448a25ff19f85a83fbea32f76c5ff01654d249b6df1bb6327b6ab2442361322662b00784498923ef157f0a48366ced70ea483aff7ccf112f4dfc9f6b11539eec4051b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff4a0ea0845f6a278764dbe9f7f9e6cc0a6ca64a900ab2554d8461a34f36af234ebd8710a04b63dd4cb77cfe82f4c8b3a97d9e5f9a4e787b66ea01843653d961bf5617f0940c7ae34044b132583b3459b5f84786f58486f7aa58f1d75156e283274b7d261713f40301;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d124d6ec36dad3ee1a5dc4ff23040b1c2748a930f019e8d9eae0182a291f1ed18adfe9748d6a1a4236b2b15252bed6397cde639d6fb531a350534b81638edc01d2bf2dacbc2ff4f32c223abf0897de5c66974cc60c62d716b5126667223d7e3ed2d458a2cc318f661;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf22e216b8561d8b322db410b01e5895f63932bb3372da2d7f79115d372bf9d89c78224f5c3ee9114ced6428de63a6d5f2b75f443d6503d1b7c86a419a6912f50043988c6373114b6af3c9d5e8c379da42b807bf87e87ec3156ed7eaa854dcc84f1ffbeb7af75bab8c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143b948b8d4b28c94f1baf2428e2375054cd7a9d48404d30fa8f278fd87de0af635188d2abd639898fa9bb4d0db19f593ac9c5b65f03aa24b0531af89ffc16ff65b448adef96435465a4b57f252d242f23ee42e0117480c7c9050f5af3938233949998e6a2e906cdc51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f51b28c1a5eb09140daf10729ab75275fc0f54d06d51f3f9d56146e09525d3b774afac3ceb072ca565d65f50f779548f219517328f48172fd56e03bcd544fb36a3cbc2c8e9423b673cfca83b56e478a3f61f8fe48a1aa133d43bc04f5c9656902d85990df47834aa47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b22d82f42735358211298dd6922f49c6303b3589f5e867a6deb9de6c78cb5fb51ad6e4c53ef64afb574f0b630329a33cc8e9240b3fd0a07370f998b07a91af92db09b402e41fc8b93d40e5019075de8c0cbc9fcb0d54a953f6d71a6375c690cc68a8675d4e17546aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd16a01f7a41581223af08ef1fbb76cc77e676f1934720622bec8c6fe255e636ee36a925ef49b51fcc89413d73b39bb445da537f5d46687920f24edd87235119a0e592697a5443e407823a78dec04ca91288fcf920c0ca6ea77e61997a188e6d95b2c11a406dace69b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e57acec784303877d81bc0a92992739d96d2ddfafb24bf0d8ef745386a2f2c1595db2d27df2873509bf6e7036f2fc807b44a2aeeefac55a4c162a36105bbf14dd2e711b29867463756b37dad7b5d38ccca68899ad5b8aff27d27d3c35e2235515c518c3ede812bb28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195a23f94c4e991497a4d713eab4fd17ef4226f5165ecbee530e77ef66d1a83e5b5f7ae1fcd3136703e3d69e258eb0105cfecbed78a0fa5eb8475f5024cd2fd3de859b51f54b854649da5bbaf7fdd27ef7572f18653a08119379840904bacbb2ca51d2b7edfdfb17315;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70a1ef114317155cb18127bbdffc73515ad1f2120052351adc468cca791510eda04b463f2a1329d9523b104aeb897fc46494f080bb4e7ee8b1ae93b3e0d8f852a45afacaca196e16c9a57969306a6601c35181cf29cdabc50719d82ed14a496dd00fa9a5a4aaad55f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16105d34b390a121e63ca493aa3cfba27a22dafa2284f64166e26c49c871abddea20ab39fb71c3b77100bdb4df398bfda247e342d93f874ec16c002727860e7e8ec337ec69e1991e2c1a7cdbe506bd4df56d95a44061b4078cf92cccfc4ba8e4736ce73a1cf657076e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e05c56f456c5bd0ee73afde94ef3d61c587934cfdc6124f442d48fb008f9d20d175307537f2e4462b33dcd162677406dec7bb7f11e89407c9d816f564db102348092e5399d3fef84999d2d7f9a0f34f339b4dd843a4bdd359b0c988606c23d5892999bd26fc688901;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171a70d21e61fcbd207788f2b22bf573a3ba6e94f52d844ff49d504582a7b984f817ad23f6fc0353343586d070b7726ef7b9502cc5b9e0f34a4374992e46fa52dd14f80a4e297fdbaab5ec068e5c22d570437dc53aa084fe7240b1b5947a856768a8dbb8fa28e07824;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1907a498dfbf78df552fa03d3316396b9400a4a93ee54fec3068a8a23aa80eb08b5e90fdd864be148e42a6515a2ccf56f8e079075cc286c70494861dae478d5670066fdff1281ba17ee04447751737ac4f047ec9cc953f4fe6b30ced6a11c80a4605a8246f8245cd97b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h846dbc7a15847fbb0369322cc9ff415abc494bc4a98c98eb3d0a769cf3e4d74f0c5402728aaf756207e49befc10e6d1cd1fd1976ccbbb2c242517315c732581ec7fb75f7c899aca488be5ac225b4dc432c65c44d128fa659178c2cb3298ec8928b2ad2fde21440ea82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h750f2565665c773ecd439c987ec25dc14acf017d269bbd1d0d489d826a833635041772f6bbb45573deb43454f85d2a47387d1a201ff309474167fc1debcdd51cbd08621b782e18dd5acd47d2494998018bf931705043c587c35d4b2991b745e3729a635f9d8b4e4f07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bcf4816f580973830ddf81ef6e4deaa97ab0a9612830461313224632b532f82ec77e9f4bb88f88113353fb84026472393918003764bea8720dd22fe32281eeca6bb39b39be4f62649d4147802f4b719f48fb5ab4532053e92ab177572a25a9283b997c792cf9e8ec9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55edd6430651d37df1df1fbe02f5372c6a941cf32da076251012d8bd6410a6d9f97f5a2d3c34d59ac9551479672d89d4d4d7060ca8911301b626df8b96516e0d3e11f3d9793f9e060eb543a76468cbafc3b38af2babde19d2228db81d5ff415783014aa29ef9935e77;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce926b166c125da886ea3e9fbf420066a8d3706a1e231f919280e7b4cbb0a3c3b7831bbddeaf265d3d194545aa59a3abb1baf0fabee400d5fc39b0fee0093ca53e68b3289c47336d911062b911e9370d4daba4df9596c7d2067143470db82da1cb8305ecd19f120365;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec6966e260c2f8a944b4e28dcc40f8a74241dd26d285e1756aae55b774a6d5426179ced300b76abc1bdb6b67a2d1873eb5d130f2842b7b6516ab84340f4a6db2ad7b4fe2f02c8d24e276e980978b7d435793d5fd49fec7981510a0e9a2a7418ab4065df29db8ee5dfa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c3bea2d4e89db7dacf6a57abf3d81c97a82517fd59bb277a2ce2824038b9fa3605f4e188070ca2e92a1b8758bee6e03da8f665575ddb160149e7a1390470d9face9a087705965c851439b5c1b54417bbf54148fd3ddd2cf566e8e60d5dbe8b17664f18faf5e2c2d50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1315c346b779c080de139104de8de806dcefeb8843a9b4fc1972a6db17c845a18aeafde35f55375ff5edeb01bf4793495f366d019df15b9e528310d1c1081135429a2e87aa8da8a4504673726a9b7230ebfec368578c8590c92cbc61e24b48a3e2d101f267c0eb58a37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb398285046be42c4bde075819f844c88b35463d501880b83c949a48bad9cff415439ef387d8da61f552652b7037089de49819cf764b08ad3f0b8411e6add9bce998e113a500f21170550ca8d0b7c4e604a7c3773ac0888dbacaf3ed1e2b98b194e24157f656327941c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5433088f0603e2d0b2d7b638acacc34bff8cb445d213248a588747920732557123a1bf3bced543c5bd51a9782f01ffd58a8c06f5c08a122393ac10126fc4df73f0bc9436b702ce9bd7254ebd5ec0907304b4e993cbfe8caa221d9ada4448c654306aa0ac90a6962f42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104c3cbae780745c52df71517a3b558dbea0fddcfe2038d3f32b804252b6b6622a9cba16f5739480ca88d894363318c88dd7e6b00ac4157321d7f886d39e59b79b039a6718c870e38b21d0f7dfd3311bf3f9a046e2b04a7e7b82412a6f65aa274be73e2a310170c3266;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1136a648f8729d3e8af5264761bf727b62dd4728afbdc41346a7a9ba437113106bf8edf8b4f83621c72f49dcc52db70d0ce4e19bcd7861b3705b35b70ba4ca0732f7de19282f80aab1d1250b845dab92931b170c65ed2df04aa8a1e90e00b0473a4ca32d1b858b5ef6b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5082674c7050c4d263a4236e3111ed5bb3aa6e55abddad75c8fca013cdc99b8c25199addbb1b750ba4365a5c6316d38d6ac9a5ec062af3fa14665f9bad366dbc99f97f52fbeee9d8bfba916a1d1af937ee2ab8b3800dfda9715432ea478ae4017b4a390ed79ff902a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bc0bfddc32581433493776f6147ded192cbeb3bf98d350991e2efe7ee83956fa00aee24f13ca68499ee3ff4f8ed9d6af4e07615e3a9989a4840b96aeb5bef661db413c111fcdb2b0e33677228e1aa7404ebcfe0a39c9b450ce9cd5d153c368b94ee82f6119fe1f2d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27ea8bffb6fec9513795252e80276a322ce464b6cf1ddfa516c1d34ba5e0a93edf17d9226bb91f23825d7cc9a99758dba42fdab055fc35baf60d986ddff4990d61b078cf7b3ad5997136b2a6698a557c7ab9bd0ebd99b167745dd9a69e3e1b6de11c4ffa00148576cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133fb7372a05468af01ef6f6e864f6db28ed32fcc040ef6e843b0eed523f4b65c0e32bac794405643cbe1925856215a8a96f756ef85c501cceb8e1f2d786e52410664d6fd9108aacc0930bfa69b76841407e371b3a76f4fcbfe3ea9d39ad35c5f5f837a690eb80ab16d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155de4e4c1ec39d7e4886500fdd67da32713bd5eac12de523163b2f945583b0293c4978daa43cb5cd703aef065356b34668e2492057e5ad8c6035020cc6dea7bea82f21614419a708df0dfab6afe0da70a4302661b9e77513953deaf83d9500dadd067638075e7d3eae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177cc15d470feea8d8f4c88726bcc194df7e0fe5e9be8ca3a1f2175b83aba162767bef5425b457897a4fe5f44135c9b740826d5e0966915a55d63deb58e2dff41edd69bcfee00c83ba30044f18cffc4c32c28562d61f419f4be66f4522448b52dfc9f62ac19c4b1fa72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19db8ba6039fc02e9665866bf5cc17b6b7ef73a92623edf08d26ff2b5ee97a2a7d00c6dc8de4f0234f01bdff55df9b4adb7ebac8a06a064bfc1974e7b22b8f0d1cbeabaebd2c398620f4572de78ea63ca36ac9deecd99f7b98f83e0fc5323c731d70dac0c180962b61b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159c093d33dc4b1f1e3224d0205dc60931d16deaa83deea53a3a07b76447131889878699de450943b12ce243c739f27aa7024076539b6f7d26f19702356c2102839ef51d86d16e7d8181dd34c608eb37f74ea40a990f39de13e22de0a77c066c8659e92142837a18c81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144a61bdda60a51a42ac32ee3df6b1c82798c2cd5f2390cecf5afd52446f110a28f09538c90a484c0a922dca3ba27e265caa10e27be44733d26d636c2ab266425caed66fffa5a38d833b68219ff2663764835852118118cb72fc52fad76caca4c872f81b50fa269fc08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h278a102a02b026c1cedc0a8486e042d30e57694e2970da1992a89067318945aa9a51e99da5040aee4cf6e14218fb2238e0daa555c20cf11159eea73f270d89ebb38ce848629c7277cc0d2959706e414d888d4df8fdf6f5d9d5b100189f7e2070fe498182aa394861da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bb0d5e5a0389e3191b66a5e28b585a1c2585e35e7a6f9b8f04faeef3828101e71f84fa0fa6cecb44e9a7e27f9e82dc99fce1ad9b618f425aa7bc64620d272e4b480ca128b92af485c6336b283f2c5f03531e30b6e70b304965e7b91f09e8fd5e3e901bbb053cb12b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d93b0591f640eaa0c8f8909eb3bc5f1a3fe301f9ef99a677ca45eda9f855ef69457973a86e8deb48e57be054b52ca030eddf4fe7e6b0760a4ca5089323308b2adc8b59b1ca115f7cc378772f62f9212af6abf002110f6f49f39df6cb75187f8df0cfda20ce104560d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90ef4b6856e37723791a256a74f0e01545ed12b92283e90b67f1b2fbf948074afa22838cc3659ad02436229769c5388f8107091c5a458b10e66b3f395d56e490914db1bef77701e02cdf099893a987dd5e7031aba4fc2809c7f655b4e33b299e78242f71b1d1cc2d81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e61a69565ab5f26d4a58579b7d84111e87d74d3f01985fb35f874561ddbe47bd991914436b386eadb5cb92cd2dd275c7f0b47d85ab2c6c4a05184749a76d87e6fa18603c55cc2ec934c240313228e6e20385ec7cda09287576373b2b23b7364b5fb04e495d5bdb957;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9bf5ee8cc29628ccd98e934b60c4549efffb0f46fd0e6aa67052fc8f636faf275214de61086ad3b50e28e28be6fb71756e70fffbcbf027b3b1950cebb5150e7ac2b1e74561be9c23eaa263506b89a4dbec920f7c52c110a70c92e8bfd406bc8528b75acab72da5826f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a76051b44d670e3c5ee0bcec571f8f180d8d6374ce299cdc4c42c621c55924db5e22fe921c39f88f0cadac3cf735eb6354c4d92300d03ef20c55d562d231b2009dc677f1bc2b5c17c79c3ad4f16fe1eec19852b68970a0483eae3f184227c37b7c212cae2d7f55e06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126bf6fca4a01fa9d7e05475167b56eee43f94068f03653d44d25785b6309677c6981c0500611d8135328f167bc5de61ab5c56069ec47141436fab7c4a7370fd220d72195cc91851d1cab8e496d4f897ca69e82fb0ea9fd7de9015cfbc3f63fe767c25b9a5420a24e8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf46a76e92fd074c9339f403943e223edb0cd9a8f89dd9e112a5838b36beb66566e8b9267568343215b9a99ec69e3ecc3e1333f8a5f3867497e1a240d2a343ccf6e9518b0728af3fa9dd4b084d623c77f7f7a745f03d3797325826dc6b3a3e69a5cd60a4f673a4afcad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1598dca80577df887893721c9578a658b610077cb350103564d374eeb6cbf08814e655b66e7aadbb02d72ede5f991db377eb8ac0f3fb87e59d8cf5d9574da5a41eb4112088c2ee7512bb49773aace45134b0b03876dc6ae75f490085f1783b88b20e583a4e800f189;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he76c2bf20905d476b89eb41ade53e544b6b3cad74329e616b2f288f794e0501291b308569f487c8840cfdb374897bfe6eb6a7f6c331d94e3986a358f324a8edc119dcdee5901a7e3819050546e2176432e79cbd9ba51f70d6f605877f2b2deae726e52924e1ee4d8e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fcd99ffad9c8e5a65faecd10f06af9eb97ca7c22de604db18a791fefe417555f8b9b9d93482b15d2141661e56b0ae920554abf9d9f8aee82d75d93d67a95745675b7bf0911d874b54d3941d6bd9bfb47486011199c11da41b8e4bdd0a1bed33976a1637ea933e8be1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h659f5f2f37a53fb083c303d1b6f3b18a3174c13c08ae4090b3420a614cba7325ded4499968768c339bdf55a9e1f3dddf188c043310c0d9880627ab1ff5f6efb95c3eb304ed731006fd8c142d3e4f244ff193ca4f1da9e6cc1090aa6b47f14e922cd183485fd4b32e73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe5c1f15ecce87a7f59afff0978c41b04d0b238195586ead40bc141fd16b75d3304118844bb7be0fd872a31e269d2087804f8ff2b8bd00c4bfcea4987c9317425cf90dc60be13d336653e946dcbc46b8d4255b7953e85dfc134cc07da89fe64144e7ee96b7fb09b4fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h455f2195c78242b6988332a3f18281921710bd719defe2ad8e5e23532981d1cbfaa3deb99e2d2243501380656f21ce71692cee9f3fedbbf786f0096f491a477de68059b0947ad5526bd9ee531c36a0310b4ea44e8dd5fb99c02ce2e17eaa10defb92914409b6898e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a9b2a847d33300b4e5b6bb74e425e857983dbb3ae7c40a2097ff9063599f7a004ed06f0e94d5a34e9ae4f855222d27eff4d6c21134f4ed03681d866a33d837bcb6bb26fd97b15fb57ce780beae471dff7fb2dc280d94734ed3f18b2d157cfdf318808a1cf4d53959b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f90a870bf146d49dc7b87f4e89d9dee7c2aa582c0c96e0a085b8972a041128bd5e72cf6fecbdefc25ac49ee46292ee2d6a0dfa6d73e730fc6e84d081eed2eb9815b062a55a6916ac731d20b763c23319cc01d17bd9917d904846adfb1eeeaa8ad633c8886b4e71fa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfaa4638b54ad92ffee6478b53ec18e2d531aebb3895c0423fb0ff80e740edac4ff201db9df28a0122013521b814405089c5c1bb71ef7a68d7962bf72cdd0a4def0ccbeda50d0af05ae63a5c60942b80ae1b17ba25267aad3adc630327b7aa085c5f0a230ebbdc98ef5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc7a0b4829b198975e358da1da1727ae9258408b33fb5bdbfffa09cbcafffd7ad84dddbb549b122bf51de1301931a2c77747aa5e8f4a7408559cd784b24ecbfc96aa9d3c27a19529465a4855e19714ea06b3e0709c47002886da9b5de59e7b915437bc0c29b0e9b505;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1338837d11c43fd0fd6be5001e2ce380fd4de061031e3a529f6ca97c4e43fd0160b23bc1a99e3530b578a5181b6ac2f57b3dffeb6f5c5d975b427a123ca1d4e1c63b4dc7cf2e87d298f087cafeee2fb9a480cf878605a20ad3056806114f3a45fccd2788d50e2b5a1e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haac4a694cfa43e58f886b3f9d146db4c0c0fe076c57d67fba5668b72d7ca3619b33b6ebd6878aaec16aced4f3cac2d3124585501525aecf36cfd61c624a405f77412a5a5aada3ee1cde56089ede37ca1a44866087f6f39910563edb8f2d57a598389c2710d1d3706a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48efcc560c9f30531060bc7ca34ea80bd255d87a1b4be06939663b453212fa6da803870b1af654063f56e56402c9ef670cae23e264bb9e1467478ad3f292f49bb99de52577236ee792a64de56689f6ac37f4ccba5ce857c48f84f43306d1d1e24743ad548026b5fcdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h590742806cdbcf1c8e47e0d1bf3bb2122f8d2db42ce8307f5a7296dea46d75b00cd49e7ecfef07e35d528f0d96679452960ec3a8e7a81d52404b4395f6d788d089d7bcd525db53d633da572a580a177e37bb630e2fe352571311ecd1c39f965549d7261018e33237cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb28a43995d4736ae6de6fc2027bb6035f3dd7adc24a4b88cb699bfd7be24b5288cc4d1fd7e8a37dc464c00fe55c07d0565064d9f953c7e6ca1d3507ce99573f4dae1d21f36c3d2d7952ffae009e615eafe5ad56e052899eba8939819c45c73fbc4ee559b85245b2f78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e09ca45a4096c34bdd1c4e0a1cc063b8a0b473ee5c8e98dfe5bdbbca66228925f0d829a8f3fb9b58dd2bd9f3e674dd3f6c08dfcc80fb88ab4b4da39b120a3bf400384978f952720895379f16979980d64bd0bab1c75f6e181295c345c5568ccfd9829f612697868bef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bf5253e6ebd500dbc28c50828b20e989aa0db0193af73b12858f04f524167123cf0229afdffc2f26d852d91e193d8e4a2f7b904d56d620c44b37833ddd09332904c78e8e27ba5923cdb72eafefe8d70035676f94f95ab63a80d1ac2b43c432cf817ddf5172094b0ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12efee4d233298a87a7152e5970d44ccb68d58303a923af6888ca43e1074abb440d616eafae23f8247eab32a3d9af6f290e3a9e0bb20758df62186fa2526349cfe794d2533f46a408c3a7b431345d76660e5b07c80112226e7e4cca8b14c7558e86e96a7582af036783;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177803d26e8114646420aee97b5cac3719b4892bb739d306cdb26a18459c67b88aeceec5dda4e6842c1dc3e6324ca3f9144a9db2449e4cd7c5b50f54a4eb8e84d618eb5a3fd171fd40f9956db6aa821d32c2db498ab88a1e283bf068c8bdd58c7ffc93cd869e80341c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b559bfdc806c7cfdc00542bcdd1c68201fd8e72ea439ffa4bc273e91a13ea4dfc3bb5a2d2e4dcf6dfd36239e06b5967e765e4e7ca3a9f49b0539541a772b2e1d227a9c6976656b9bccfc655a39136dbdbfeb813bb376d46c6d4a4b0fb4066665263de7e49d416ed5f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36c56a15f02e11d3bbe3881f707db23e664193525944af8252c99724f09610dd22c73a6e83bf748b6b9a5d4646114a4f2de9a8e9696b52bdac226d0aedf60934dcb307afb58b07e51d503502a7a54f9da64b15cb245179ad84779c10777555c686de44c9edb8eaab26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1823cdec75b2a1fcb40847d573e29e9eaa1f85ef036d15e64a1a1a3c201aceb3f2fa34b425dcfe5f4b2caf796b416ba99556c6b7c0702ada83280f065697c474f2833eb5ce6290618c009a35c0449c98dfe2b17469750239c3410b0421fd1128953d4536836e54b88d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100eb7456cddd4191901451e91d48cfdd9ee9fe785363a2fbe4109711ec01bc59e90af9f1bc9786fb1402a17832c27e5c0541e8374f271cb5b255fff981471b1ba437dd1b47709bc64617316380473ee130c1ad237fcd2394f20d4a9f796eddebac519e3d7680af0b9f;
        #1
        $finish();
    end
endmodule
