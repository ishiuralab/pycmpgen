module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    compressor_CLA32_16 compressor_CLA32_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA32_16(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [14:0] stage1_0;
   wire [9:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [14:0] stage1_4;
   wire [16:0] stage1_5;
   wire [18:0] stage1_6;
   wire [11:0] stage1_7;
   wire [13:0] stage1_8;
   wire [14:0] stage1_9;
   wire [12:0] stage1_10;
   wire [10:0] stage1_11;
   wire [15:0] stage1_12;
   wire [17:0] stage1_13;
   wire [16:0] stage1_14;
   wire [10:0] stage1_15;
   wire [8:0] stage1_16;
   wire [4:0] stage1_17;
   wire [4:0] stage2_0;
   wire [11:0] stage2_1;
   wire [1:0] stage2_2;
   wire [9:0] stage2_3;
   wire [6:0] stage2_4;
   wire [8:0] stage2_5;
   wire [5:0] stage2_6;
   wire [6:0] stage2_7;
   wire [6:0] stage2_8;
   wire [7:0] stage2_9;
   wire [5:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [15:0] stage2_14;
   wire [3:0] stage2_15;
   wire [11:0] stage2_16;
   wire [6:0] stage2_17;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [4:0] stage3_5;
   wire [1:0] stage3_6;
   wire [4:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [1:0] stage3_10;
   wire [2:0] stage3_11;
   wire [4:0] stage3_12;
   wire [1:0] stage3_13;
   wire [6:0] stage3_14;
   wire [4:0] stage3_15;
   wire [2:0] stage3_16;
   wire [7:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[4],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_3[25]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[5],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[6],stage1_4[10],stage1_3[10]}
   );
   gpc606_5 gpc11 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[7],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[8],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[9],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[10]}
   );
   gpc606_5 gpc15 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[11]}
   );
   gpc606_5 gpc16 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[12]}
   );
   gpc615_5 gpc17 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28]},
      {stage0_6[18]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[13]}
   );
   gpc615_5 gpc18 (
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_7[24]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[7],stage1_7[8],stage1_6[10]}
   );
   gpc615_5 gpc19 (
      {stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage0_8[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[8],stage1_7[9]}
   );
   gpc1406_5 gpc20 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[9]}
   );
   gpc606_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[10]}
   );
   gpc606_5 gpc22 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[11]}
   );
   gpc606_5 gpc23 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[3],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[12]}
   );
   gpc606_5 gpc24 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[4],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc615_5 gpc25 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16]},
      {stage0_10[22]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[5],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc615_5 gpc26 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_10[23]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[6],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc27 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_10[24]},
      {stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage1_13[3],stage1_12[7],stage1_11[8],stage1_10[9],stage1_9[13]}
   );
   gpc615_5 gpc28 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_10[25]},
      {stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30]},
      {stage1_13[4],stage1_12[8],stage1_11[9],stage1_10[10],stage1_9[14]}
   );
   gpc615_5 gpc29 (
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_11[31]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[9],stage1_11[10],stage1_10[11]}
   );
   gpc606_5 gpc30 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[1],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc31 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[2],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[3],stage1_13[8],stage1_12[12]}
   );
   gpc606_5 gpc33 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[4],stage1_13[9],stage1_12[13]}
   );
   gpc606_5 gpc34 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[4],stage1_14[5],stage1_13[10]}
   );
   gpc606_5 gpc35 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[5],stage1_14[6],stage1_13[11]}
   );
   gpc606_5 gpc36 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[6],stage1_14[7],stage1_13[12]}
   );
   gpc606_5 gpc37 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[7],stage1_14[8],stage1_13[13]}
   );
   gpc615_5 gpc38 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_14[24]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[8],stage1_15[8],stage1_14[9],stage1_13[14]}
   );
   gpc1_1 gpc39 (
      {stage0_0[21]},
      {stage1_0[4]}
   );
   gpc1_1 gpc40 (
      {stage0_0[22]},
      {stage1_0[5]}
   );
   gpc1_1 gpc41 (
      {stage0_0[23]},
      {stage1_0[6]}
   );
   gpc1_1 gpc42 (
      {stage0_0[24]},
      {stage1_0[7]}
   );
   gpc1_1 gpc43 (
      {stage0_0[25]},
      {stage1_0[8]}
   );
   gpc1_1 gpc44 (
      {stage0_0[26]},
      {stage1_0[9]}
   );
   gpc1_1 gpc45 (
      {stage0_0[27]},
      {stage1_0[10]}
   );
   gpc1_1 gpc46 (
      {stage0_0[28]},
      {stage1_0[11]}
   );
   gpc1_1 gpc47 (
      {stage0_0[29]},
      {stage1_0[12]}
   );
   gpc1_1 gpc48 (
      {stage0_0[30]},
      {stage1_0[13]}
   );
   gpc1_1 gpc49 (
      {stage0_0[31]},
      {stage1_0[14]}
   );
   gpc1_1 gpc50 (
      {stage0_1[30]},
      {stage1_1[8]}
   );
   gpc1_1 gpc51 (
      {stage0_1[31]},
      {stage1_1[9]}
   );
   gpc1_1 gpc52 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc53 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc54 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc55 (
      {stage0_4[31]},
      {stage1_4[14]}
   );
   gpc1_1 gpc56 (
      {stage0_5[29]},
      {stage1_5[14]}
   );
   gpc1_1 gpc57 (
      {stage0_5[30]},
      {stage1_5[15]}
   );
   gpc1_1 gpc58 (
      {stage0_5[31]},
      {stage1_5[16]}
   );
   gpc1_1 gpc59 (
      {stage0_6[24]},
      {stage1_6[11]}
   );
   gpc1_1 gpc60 (
      {stage0_6[25]},
      {stage1_6[12]}
   );
   gpc1_1 gpc61 (
      {stage0_6[26]},
      {stage1_6[13]}
   );
   gpc1_1 gpc62 (
      {stage0_6[27]},
      {stage1_6[14]}
   );
   gpc1_1 gpc63 (
      {stage0_6[28]},
      {stage1_6[15]}
   );
   gpc1_1 gpc64 (
      {stage0_6[29]},
      {stage1_6[16]}
   );
   gpc1_1 gpc65 (
      {stage0_6[30]},
      {stage1_6[17]}
   );
   gpc1_1 gpc66 (
      {stage0_6[31]},
      {stage1_6[18]}
   );
   gpc1_1 gpc67 (
      {stage0_7[30]},
      {stage1_7[10]}
   );
   gpc1_1 gpc68 (
      {stage0_7[31]},
      {stage1_7[11]}
   );
   gpc1_1 gpc69 (
      {stage0_8[31]},
      {stage1_8[13]}
   );
   gpc1_1 gpc70 (
      {stage0_10[31]},
      {stage1_10[12]}
   );
   gpc1_1 gpc71 (
      {stage0_12[30]},
      {stage1_12[14]}
   );
   gpc1_1 gpc72 (
      {stage0_12[31]},
      {stage1_12[15]}
   );
   gpc1_1 gpc73 (
      {stage0_13[29]},
      {stage1_13[15]}
   );
   gpc1_1 gpc74 (
      {stage0_13[30]},
      {stage1_13[16]}
   );
   gpc1_1 gpc75 (
      {stage0_13[31]},
      {stage1_13[17]}
   );
   gpc1_1 gpc76 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc77 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc78 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc79 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc80 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc81 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc82 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc83 (
      {stage0_15[30]},
      {stage1_15[9]}
   );
   gpc1_1 gpc84 (
      {stage0_15[31]},
      {stage1_15[10]}
   );
   gpc606_5 gpc85 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc86 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc87 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc606_5 gpc88 (
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc89 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc90 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[3],stage2_6[3],stage2_5[3]}
   );
   gpc606_5 gpc91 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[3],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc92 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[6]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[1],stage2_9[2],stage2_8[4],stage2_7[5]}
   );
   gpc606_5 gpc93 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[2],stage2_9[3],stage2_8[5]}
   );
   gpc606_5 gpc94 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[2],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc95 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[3],stage2_10[4]}
   );
   gpc615_5 gpc96 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[4]}
   );
   gpc606_5 gpc97 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4]}
   );
   gpc606_5 gpc98 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[4]}
   );
   gpc606_5 gpc99 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], 1'b0},
      {stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[5]}
   );
   gpc1_1 gpc100 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc104 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc105 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc106 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc107 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc108 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc109 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc110 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc111 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc112 (
      {stage1_1[9]},
      {stage2_1[11]}
   );
   gpc1_1 gpc113 (
      {stage1_3[5]},
      {stage2_3[3]}
   );
   gpc1_1 gpc114 (
      {stage1_3[6]},
      {stage2_3[4]}
   );
   gpc1_1 gpc115 (
      {stage1_3[7]},
      {stage2_3[5]}
   );
   gpc1_1 gpc116 (
      {stage1_3[8]},
      {stage2_3[6]}
   );
   gpc1_1 gpc117 (
      {stage1_3[9]},
      {stage2_3[7]}
   );
   gpc1_1 gpc118 (
      {stage1_3[10]},
      {stage2_3[8]}
   );
   gpc1_1 gpc119 (
      {stage1_3[11]},
      {stage2_3[9]}
   );
   gpc1_1 gpc120 (
      {stage1_4[13]},
      {stage2_4[5]}
   );
   gpc1_1 gpc121 (
      {stage1_4[14]},
      {stage2_4[6]}
   );
   gpc1_1 gpc122 (
      {stage1_5[12]},
      {stage2_5[4]}
   );
   gpc1_1 gpc123 (
      {stage1_5[13]},
      {stage2_5[5]}
   );
   gpc1_1 gpc124 (
      {stage1_5[14]},
      {stage2_5[6]}
   );
   gpc1_1 gpc125 (
      {stage1_5[15]},
      {stage2_5[7]}
   );
   gpc1_1 gpc126 (
      {stage1_5[16]},
      {stage2_5[8]}
   );
   gpc1_1 gpc127 (
      {stage1_6[18]},
      {stage2_6[5]}
   );
   gpc1_1 gpc128 (
      {stage1_7[11]},
      {stage2_7[6]}
   );
   gpc1_1 gpc129 (
      {stage1_8[13]},
      {stage2_8[6]}
   );
   gpc1_1 gpc130 (
      {stage1_9[12]},
      {stage2_9[5]}
   );
   gpc1_1 gpc131 (
      {stage1_9[13]},
      {stage2_9[6]}
   );
   gpc1_1 gpc132 (
      {stage1_9[14]},
      {stage2_9[7]}
   );
   gpc1_1 gpc133 (
      {stage1_10[12]},
      {stage2_10[5]}
   );
   gpc1_1 gpc134 (
      {stage1_12[13]},
      {stage2_12[5]}
   );
   gpc1_1 gpc135 (
      {stage1_12[14]},
      {stage2_12[6]}
   );
   gpc1_1 gpc136 (
      {stage1_12[15]},
      {stage2_12[7]}
   );
   gpc1_1 gpc137 (
      {stage1_14[6]},
      {stage2_14[5]}
   );
   gpc1_1 gpc138 (
      {stage1_14[7]},
      {stage2_14[6]}
   );
   gpc1_1 gpc139 (
      {stage1_14[8]},
      {stage2_14[7]}
   );
   gpc1_1 gpc140 (
      {stage1_14[9]},
      {stage2_14[8]}
   );
   gpc1_1 gpc141 (
      {stage1_14[10]},
      {stage2_14[9]}
   );
   gpc1_1 gpc142 (
      {stage1_14[11]},
      {stage2_14[10]}
   );
   gpc1_1 gpc143 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc144 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc145 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc146 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc147 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc148 (
      {stage1_16[0]},
      {stage2_16[3]}
   );
   gpc1_1 gpc149 (
      {stage1_16[1]},
      {stage2_16[4]}
   );
   gpc1_1 gpc150 (
      {stage1_16[2]},
      {stage2_16[5]}
   );
   gpc1_1 gpc151 (
      {stage1_16[3]},
      {stage2_16[6]}
   );
   gpc1_1 gpc152 (
      {stage1_16[4]},
      {stage2_16[7]}
   );
   gpc1_1 gpc153 (
      {stage1_16[5]},
      {stage2_16[8]}
   );
   gpc1_1 gpc154 (
      {stage1_16[6]},
      {stage2_16[9]}
   );
   gpc1_1 gpc155 (
      {stage1_16[7]},
      {stage2_16[10]}
   );
   gpc1_1 gpc156 (
      {stage1_16[8]},
      {stage2_16[11]}
   );
   gpc1_1 gpc157 (
      {stage1_17[0]},
      {stage2_17[2]}
   );
   gpc1_1 gpc158 (
      {stage1_17[1]},
      {stage2_17[3]}
   );
   gpc1_1 gpc159 (
      {stage1_17[2]},
      {stage2_17[4]}
   );
   gpc1_1 gpc160 (
      {stage1_17[3]},
      {stage2_17[5]}
   );
   gpc1_1 gpc161 (
      {stage1_17[4]},
      {stage2_17[6]}
   );
   gpc1163_5 gpc162 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc163 (
      {stage2_0[3], stage2_0[4], 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc164 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2]}
   );
   gpc606_5 gpc165 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc615_5 gpc166 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[2]}
   );
   gpc615_5 gpc167 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc168 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], 1'b0},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[2]}
   );
   gpc606_5 gpc169 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[2]}
   );
   gpc606_5 gpc170 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[2],stage3_14[2]}
   );
   gpc1163_5 gpc171 (
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage2_17[0]},
      {1'b0},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[3]}
   );
   gpc1_1 gpc172 (
      {stage2_3[7]},
      {stage3_3[3]}
   );
   gpc1_1 gpc173 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc174 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc175 (
      {stage2_5[6]},
      {stage3_5[2]}
   );
   gpc1_1 gpc176 (
      {stage2_5[7]},
      {stage3_5[3]}
   );
   gpc1_1 gpc177 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc178 (
      {stage2_7[5]},
      {stage3_7[3]}
   );
   gpc1_1 gpc179 (
      {stage2_7[6]},
      {stage3_7[4]}
   );
   gpc1_1 gpc180 (
      {stage2_8[6]},
      {stage3_8[3]}
   );
   gpc1_1 gpc181 (
      {stage2_9[7]},
      {stage3_9[2]}
   );
   gpc1_1 gpc182 (
      {stage2_12[6]},
      {stage3_12[3]}
   );
   gpc1_1 gpc183 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc184 (
      {stage2_14[12]},
      {stage3_14[3]}
   );
   gpc1_1 gpc185 (
      {stage2_14[13]},
      {stage3_14[4]}
   );
   gpc1_1 gpc186 (
      {stage2_14[14]},
      {stage3_14[5]}
   );
   gpc1_1 gpc187 (
      {stage2_14[15]},
      {stage3_14[6]}
   );
   gpc1_1 gpc188 (
      {stage2_15[3]},
      {stage3_15[4]}
   );
   gpc1_1 gpc189 (
      {stage2_17[1]},
      {stage3_17[2]}
   );
   gpc1_1 gpc190 (
      {stage2_17[2]},
      {stage3_17[3]}
   );
   gpc1_1 gpc191 (
      {stage2_17[3]},
      {stage3_17[4]}
   );
   gpc1_1 gpc192 (
      {stage2_17[4]},
      {stage3_17[5]}
   );
   gpc1_1 gpc193 (
      {stage2_17[5]},
      {stage3_17[6]}
   );
   gpc1_1 gpc194 (
      {stage2_17[6]},
      {stage3_17[7]}
   );
   gpc2135_5 gpc195 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc606_5 gpc196 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], 1'b0, 1'b0},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], 1'b0},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc2135_5 gpc197 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], 1'b0},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc615_5 gpc198 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc2135_5 gpc199 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc117_4 gpc200 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc201 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc202 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc203 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc204 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc205 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc206 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc207 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc208 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc209 (
      {stage3_10[1]},
      {stage4_10[1]}
   );
   gpc1_1 gpc210 (
      {stage3_11[2]},
      {stage4_11[1]}
   );
   gpc1_1 gpc211 (
      {stage3_13[1]},
      {stage4_13[1]}
   );
   gpc1_1 gpc212 (
      {stage3_14[6]},
      {stage4_14[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor_CLA32_16 compressor_CLA32_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd340fcc339af61888ba31a45d8689d2f852fe757785583e7b65ab7356099aeb4026b42e135221753662a506490326f2fb7b4cc045816dd9d784f25b4caa0ca22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfcaaca3bbc1acae3c9e24c4ff889e7db89c54bc1c63351323a346c68067b38cc7a753497ad466e0b6a92a040955bb0d632a7b995a629d4286a6849c9fd1481c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h228996a6132ec9c0a7ed207c2e4c8eb40d39a45bbc29806fe6827be63e2b796159424ef825516cc0eb63f198039d3f335660e32f5a3ea21e66bb7446bfddd905;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h60e6c011f1f2d027f127c5a6a400f7d769f0d8a32cdf6e03b7f49ec1cc3d01c5281f504e69746726a57df7c40d6c1a702569221de6186f19647aa27951438a92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf8019e15e2fe6dad85f7ea191c694919b119446cc7c4478d9d5f359711a5c7b41f0f65e68fb2448a56e0935cfdfce5d8b9966b1327e4c22291ff404da9cb40b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h18991ec9187856c1e022540382c49651c6cf5c0c0785841231661134d9e673a9ce51b6e1603516bd25175233cc51527759d0ee2e87ff6f8684373c5a599b7ba1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h530dcc0cec715e50943f4a1bd9fa7f5e133c24f69346c5e8dcf6c0cbcf939dd90ef734f80ed823ca06d15ad8b53071bd19e521227b11b586d9951162381b3751;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h255be106a0cb13cdfa51a32935480ed8cf3ec75b43af13fdca2bdeb5e14fe3caffc10371bf1ad57eac2184f505c7cadf4eb9fee3cd3d7fb76ecaa12c84885d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h92c26e59b81d892167096b5544d3deb04e9d27f6210fcdbfb431a5cc4b19046d4affb519481acc9d4e4573b645881790ff092f887af5ad50137987f834dbbdda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb35afa7f791c4bd5b8db88f242f18c78cd9891fa256e411ecd478a23f40049498f4bcbdcd68c10d9560621ac789a6040ba419828e20eb9c5596eb523e6c80ec1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha3b0c6ac790b5855cb860185292d9ffc27dee0419690ef65dd172f185bc885c7304ed28ef3abe4fc4d79d216b07889ce773d5a5c1144444096174faa486142b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h744076c61b10f1f30e862d22995b245b8b29a0255d223b5011cc86b596a50d6c368690fc6c150581130de434677fdf9eb66e5217443b9790ff188cffc2c5a1e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc93ace19f11b805e1ee2a85a749a6f42b0e9736e9087b39d0eb106d7a92061c2088008b952633a6d372a4940dea6199a4faaddc4941161f76c1b1e788fe0beb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h969ab52174249943b071c9bf0e075892fc81790d24d29c1abb40e6c447f05bfca022f04496a53b2b13743abab5fa8e32af7ecea81302e75e491246a9142eb733;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb4281bc57914529b55874ae78859cb2ea214db1b785766cea55d060965eb0438fb10693af88939fb3e311012cbd67375c3695a47e093bebd30eb2f6135914bac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h54a0b1d4d13c706cb9e276468962f9fd24381c297b94b1653715772f8b0ed99318ea99f5b317f7af11ce878dca4b5f96d3e17aaa5efc74b731c9fc27bfcbb244;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8ee95aa0083f7fd1330973fa80232660c008e1610b3cef88faeff74c5eced67c0509b329e7c2c82b6a9140bc1632fe199454eee28111b707ffda1adf3f50efaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf3e8f54547670279c1c94edab1538c8d783986578714f42ab0b1a17c9809eb5ef6e68dbb984bf0bf4301a38f380dac7f3de95b36b59c69882d158775e1084b7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8ce171f03ea404a10873f88b73833f265738c40a6fef75d8bb83f92a54ff5ceb15c504abe2032ee7dff047130e10b8756efe611d0e5078decfdf0768e02c46f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h52f074e2bab0176b870bbdd4b193d213ef2ca696700a79e058261dfec50d6436fe9b8c9d9600e419f244542eb37eb53a56a7da3527a3761bdd93747cf1be9bc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hca5ae900ca1fd6ca2f34dc863d3160cdf5ff6d120e468f9040b9ee0d0eb2b2700c903e9ee9bf1961eea113381a468e534987663ba639dd89b1e3f936b884ec1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h73c379b10f5a1a98a3dec39ce18244f315074d0742092175a81387ec4395ed7f086d292ce79783744ec4dfc24aeada07120ab37c07130cebf340f90f1615a210;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8a6ceab4db45ccfe996521cf038d203001e3f68d8c17e8513a8a0bb7e1bca2feb37627222d7d93b62db6ed80b2ce3d9b571bf9ce454b834acf90d75e7c186e47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdd7ba34de27c1f23b55ae2082c7368515a3ca3c76e0fc4740da365d4b74a78357ddec8e176a4ec8f0507a69b952f0f58e0a2728d3ef1aa64b8b32df60ce228d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7533c677046ab0d6f76e4faca477ce1746af8dd285b5999aa693ed67d4efe1f55aa40f3e30434005e5942ee6edd2c859104b046b1e204ea0134d8cac71469fbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h773019af64263cac01b34fa00823350eeeed4ac21693861cc1caf57831c7740471e3dffac6d467e06ec3cb2d072091f93cf64587adf79f5748e01397ed0c0685;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hed9307b0c32ddedd3445b784a7ea9d976ca08608c17aee84e3edb1cd6ebdebaa5fee494af207be61f904da350a1778ee1e78220818937022b1b607ec6a191a55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h99d356ec5c6289f11876133336baa568144caabf6890dc1ea54f805a45cf651c7ce7dbfacb32ae2686177eb4065025c5f9c810ce132654167f1b4c5626719743;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he6041755bf56d009cb41b4c98e3c838db2929874e879d598b90ec0626936168d2d2fc6f3531538e1df0b2e645f602a388417af83dbcf603eb18b8fa33b2a228b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb8e70c428f27bf23510aa4a223234802adf1c0ee1f5f02bd239b9dbd575a9fec7273562b6a723936e1da79cf6949a1c789d972f2493800802fce6f9e9607ffb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h664fe740fc76fcb6f39741de1b148fafe9de01c66a3b4bdbe745c48e50ff2c18d56cd719d203a2a8e082b8938d1acad9708585ede9b4577d28d6dbe4aa43bf4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb7a6e41f133e44c4782b87b75bae7166947b8747140cb98581fc4c6aaae10e1bed497f8b19d4cfef64ec9bc79db6b5da8e7514c0542e384fc204c4bf9d8f498e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hebf164776361df1e471671cb51fb45fe42b2398f2e3dcc30f6bd19b460c35b00b333b11f086b2459f1101646444e856ae0cc140a7b7a7a6a8f9814bde9c070fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hbc5228e5ecefb9b2b67080f5b5ec84bd1bbd1bcddfc9352a5a77176f82f3eebed6ca336c9cec604ecacc3cf8842457d0683cc215cd51613a9394cc743208fa02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h617ad352b797685f3a7f4f5ade985eb429abd5d4748fe18abbc29c18f30abe0835d2bb206da48cc8134c279a2cc8e5efb60d1f3e775da44a3a44c170f4d8effb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h457db230cfe22c9ed4f447b09233ad44f252e898c58239f7adedbc8e318e9627fd342485b1d4e21cc973aac327edbdb0b4e0a0bf5bd06f6c3f8a72e52a9956ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9c9ca3bb6233392e0efe8a41f8a1bbc866dc816eb3ac507bdd48ef9ad665383bba627a7c326e8e9e899e9240965733e33ad958d0e676ddb2e4f14addde6acb94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h953a9c6d36a7600bf9a2efe91d04a070392badbe132fa1b5becbda674ad385a5645e9dd9fd1a30704394e0040abe3b56528298719cd5e14198d979fd40910814;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h34112fd409dc7251e068c1e51b3cc7bfb4cfce6e59ecb2319273a74bd1f350afb3c90de15b51803aaa46a8256047849dc92d2ece4911f0e8fb8f8c568a4fe63e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2e8ce0bcda9d5688adfcf1df6c21959f3280bfb0a416067b1579aac92bc2d448773a4f78a7e1931f91d1a120f70dc226806ad1a8cc1b9127d3aea1e4c9a9a9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hbe52143e5fceec03f2c6e9937780e4b7dffa15ab23bb1e9af85d9941c69276474cd884fe615b69e46a221a82be8673a243b435cfb4cc56cf011cd0ae35220a11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h799750afc1fb25030c267b437264ca15fd246fda51baaf94c4206c6bb4b0602bdcefd38a829cd53a6ee54bfb1417e307a54f1f5bdfb3c97f6c85e5b7c1b49921;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2e9718a86f5ffd029cbe42bac39225ede07766778c37de586b25895648b441b847bff8d4ad14b4878038ebeeabd514e2249de29ac3beee2d62bd500218dfbac8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haa3eb812715c53fd657f55f2ff1c6c41d8d8efbde9a7e5734761b5bc5f16d36d060c8b144c8172984120eb1193e6fd00a24d0e1cfed0f6c91df7d7c1dbff1078;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcc7ccdbf5e21f53d3f0c6688d5d8aff256e97f321f95f4589dafda67a108ebaf32d4a75eda26a9f18324de89bb51abdda808fc5ee6caebabfea8e3fe54a85a11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7a76a08839dbd13664fb2d0ac09e88cc3cbe3ab7fd21866552ada78e62f932751c5aa9f8eb89243eba8581f91892096f1d7ce7c840c7e3c75c0804229ad623c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5a77f662a831004a7007047df3fe2ad874cb9d142a0abcb0634961ca4a94ce1c0434fc8f4a8792b6f142db4922479eccb5b499328ff4be715ee390bbf754bf06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf204d03fad0febe7a37f98e0592a4d166d1c46f45baaef6bde87b91337e39e24e3ced1a53eca162152fcf88c25cb172dbadfc2960b506e16d2025fed6f39b8ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h15dccaa5334bee0effa1db92be1e3abc448409c65a0deb714656e06ac23243d2735bd8e74edea5b3c3ceef7447172c24dfc90e6734cde51e83f630397032cb6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc73a728ee8968efebf15f026388ab17bf8fab2b0316ad973c5c631117ea2cb9f8cc19d757cfdff68d9e250a95960bc91724e1f15c58ad7d081abfada0c1bbf7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha1c30c1eb983aec3a840a5210b5b93b0b6b4331538b95229e4f12906784162bfd16f9a29d2819772e0e889ff68c17b127fb6e7497c61cb920b57bd351dce879d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h403d173f11b9e5041f47baefeade5f6f909c51ab722365fb49ae259fb32d2786ce723d25b5634e297667c10d4c5c620994b2819dc4a40d321b3ca9d1374a08dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4f99bb349a020587d68a9978814e54dde3c79d6f75c0a5a5b87db9c5aaff2e78ca4bf0b90220e3183873cdc51276f22fdcf8caaab8e1b09d219579b1f08276e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hde13f151232da5d52a2e3d5355296f9560dac07ebc890f4ee72bed1fd25c64b32446275c14649107ff7933a4fdff7190fa21e3085e339f561eccd9401fafcc7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9c555d4a2f7114d7270fb13ff7dce43e9573b3141f9a1c1d2496b67da0431c7fa9ffda8d52f5672706c8ec9cd33ffeb1802d5f60b906e0e52d2957d7dafd82eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4d0408cab3cf6497b0b19bb98a9f3b44ba069d05c9e9e63ae7d370f29c06468635d76da67642c8775ef8b8b0f20d47d1b46cacdd63e5db26bc9a80338de58c3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h55a51717368a30b12bcbe00370d370fbb8a02140762998bd528d8d2ad53b09d2e1f2dfe03e95d1a93071cf2ff4d74cfb756b9cc9b4db0f05753b55591ec5eb77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h97d35a4c7f8f0e9b7872ef8f1c73dc916948682868cace1306500ebfd9b2f83f2f88b08bc88534dc625c7a91aa4df53390be0be44ce84aa0928b92ec5d789ecf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hbdde572b3f2dedc0bf041d19f3234805b9e2570dba9b35537e54704b0404a9c5579c6f5aa7ff446d47af41815777ba59fc5433b96927f9f2176a0ce11e642640;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2ed4d98310a042864525414936fcbada44f58a40e55925c6500a8b61224b487977bc6b45bac5b26d5bd3ce62974949cfc1803177fb8a0b70445a3d9cf5fbbe2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h924fa9f8edb190d005acc3b7027f19aed7770fd099dbcca1cf0566f922d00e63601a5864bd2eda28f5294ffb5670c08df77e4ee0bd436d1ae32c9c7fe1188b11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3674825bcdbebae4be998cdaaab9896c4aaddc1f649b6c3d85bbb7ea17f9a60cd13286dadacfc6ba98757782e07251283b7f336783c240b632797cff6c3c81d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfe803a868d06cfd781e6ecc74986a0bad05f426ded165208770a066ca1e534e021057478a6c59f24c6c40a2ec30687698a7a7a169cd5486144b2c65d1753b0d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hde9044e31b5803f57e38028de06d1b28bbbc7a8de549dde733a496409c1e8d533dee5a744992098a4c99ca6c5670271bd5ddf3fb36a7301e7a1de3fc1b23396e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h41dd6a57525dc4f495446569d8ef2cac9146f989f4dc72efece79dccfea21db567cd5231980b3e16a9faa2f95e051ec445f4d9fb96fedaf7dcb4d816dedcea0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h301d1782e9b8cc39ccd114ffe7f9ed9218ad03934b00b2162241bb9f12d63c47cf51053e1ca3cd74cf5563ed6af75c3efa3d4bfccc61669a19041ad70316fc97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hba5c65084454bffc8a5a76f0b043a8ef549deb308198db64e214428ac1de9f867727428ed2c65a6944619d9bf57b23e50822d0ed94b7481ceb91c3cbf7aa5264;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8660afa3358e8720e62b18a15f32bcf84e18cd1ceb0b0fce9000737f08a9b9b06c981247f81dd20fbb8419817fd73782e792349dbc8e9f965da066941d9c13e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h454823bdcec3c7fcd6e25a7a53f4c8559e62689c9f9f4571cbba27564a3d23850d820c74079225462b231d8f3941d2754c3c5b6c5354e07865955571da90f556;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hec5fe2331c608d93aae6f72d7434d615b4f9c3082e32c0e9300e9923098bc7261aac08ee1828e713551de05c07c706b278a6f95c8a5f2656f003824725e1b96f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3dc69bc9351aea54c820689f3e203a3cb26af5a9352cdef562077f2ad1670bcbbabcb86bb66b4f741979d1a9d46192877e246a9bbae766417fec2893f3ab5c62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8e74269202eb778447af67a221072639d14d9fe6d0377792244fce6665f3cdc6bb051090bbbc3c0e842a6f2385451d8200c886a2f9e2cd4bb818f4c9bda8a1ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9e86f21e3edf3691e8b1bc2350e318b4788986fbd0204788c85612eed45170da81c0f5cf9626adc02bce36eb2018eb4d73682d9aaec39f59a270082aaaa81adf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1aafa548548049898c4bdead6a6c95fc8d8c313b63fe8be5ad4c02539bd917765322e0cf3a92508ad6ce3e299c15accd03541db034324945835c6eb41f96de7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h49e72b3a64ad803b9aac6a0bc52c65379e11e1452badeab9f7c4644c84b28e4c7df95a0331c4c0b39d941ec6ac809ecd0a64eccece0787b687b3503b62962d3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h943b73cb6f20740239917b93b81934c9c65e4efd7be599ec51b4e85b45e3bdba1bed21a0ee5ab10ae70fa0fddd6cca3266093c9898158ab16f90522e0c00876;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc40bd77ba9c312b49d64528de75305734985781b8e519f2e0f8ba84074fd6f51a023d6bcd066cb5e987e63c552516193985138f76d3133068b96b70c70668106;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6c8698ee0a365833d23e53316beb65aa208e96f4d9b5cbc9962e732c7bf9c5a181813627cdaea18eb2e030141e82d313935aff1d4f96ebb59d3379b434cb6224;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2d13622706156a48d35ac6fee27ff062751f3392c1f5d9e36d3c699daaf0ba0096db54edd3bfb0214637bf63292969255f7d5383f639de18ff8d4f8ef6301201;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8e4969c1783cac506fe77491d107a1e615440f96f29b319c6c5b036c60c9e31e61b374fd1f8f02d0576db9824fc7d2c608419afe9b2a319d2fd39ba618a1669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5398f9d7ecbebca75aebc5579e462da51ba4cca2ab83dc5fea6940c9228fef818ddb9d561aaf7b73c44b3cd6897462b4cb95218c9273d8d9ee8b8786b1bd8c99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd928bfe1edac89565e49a22ae31285d306c6b1731d547e5fb6a5865a8f77db663fbf63535ef60229c79bb6be30943fecbf931e6b2dcaf52a089a9fa22d7094e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9e3baf397a791f47acde23c661f4f500055b544fe62371582958554adde076497aa00db32da0c578aa345a14757a2dc8bdddf7df5676b731546abd4c2a32eb80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha875ff273379a7b3f35cf048c00537b3e3de721c3d174f5381e8e27ad3b8571ca0ac60bf729955cfa5d095b47e50085523771320bc1bfe3b646bd9f3969bac9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf31bab01c59916f84fed568ba7ebfe5d0904d3a7d90e953a9b699474a0182b9dc085f113e489a420507cbdf5f3affb52a6f5f7368ff0d6edcacf1354b9c628f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he5bdc98d3eac048b8cbdde539df15b520f7dbda43feff1c664105135bb01f9c68376d5e88198ba7270b5d4dae0ead404abe110f243cf0a482f672c0b1cb3178;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hce161df7acc9fee8a4840cc15785d0cc0290236280f9655c17065be1664d0b17168e38a8eb67d94d75fabfa2de6244edc61f101cd282de12e27364c0297dd4db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd1ad1f3bc4711017138d38d03ca770fbcc3fcd42c158487bd04131d4b275d5a154986be7363915e8fdbd1cae62f3bcb591bce3ade684372d274839af1fe18b09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h49757a1518d3fde782f738c280ed2ba0ffd8fa02941048b7d32200276a6516329aa205eae1962374bf926b898465fe35cc25fd9f0ace24c887fe9bb4b3504a41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h57fb50df9c3f3c2deadeaaeb4fb3349c0fbb23b5b7c5578f13ca787782c90db1ced1e657e2dc47045a236ae62f25a77ac240048d93b52f05c597ac923c0a2ad1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5b75e7ad8327973fa4a729f6b1ef444b5e59722f259714a386774afd957ff6a2cf3f50136edbb9a2865b3322993047502cc66cf49137c5abeb65ae908acbb24e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2be3250edea377457a25aa5ef17ae55cc8ee73dd82e57711f6b72090cac4e90da3d5fdddfdbe999e26693906b1383b4c06a8ce65ec5eebbe14e2f90287a497ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'heda6dcbac82dac242dd38f1f6d4574b275c3a2c58696f649dca8e831b64434351ebb836f6a4a9eb4e55a9c7e56d5b711fa80637a5707cbdf8a6d61d6d12dc4f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha35198f4b55376d3e9968389c14ae28c97b80e627bf9b46bea418f6124aee6255111364e9b9f92d15211337266ce592e2ec477d4b96a99fe7c686e20c27f9b93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf06b0b4313af9fe248c313e042b2e696ccbadc4732ef7e2bb0b26b8b5a2bc3ac7d041615808aad8d20d2b72e2829f91eacd55ebeb659e965b148dd0a7b32135f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h11eb064503d5043037232ecd3988446f108d0f0ad80260b235939ecf06620c854f67b1b67102eee8a5b4f95aaaa65f325d7283f3c48a5280bc365fa87c3ddbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h273aa62dbc2ec108c7f220e7912177bd9cfec0e9d807b0a02c36488c973feeaf9d799eacec4cfb39e4e3312aec94edc1bd3025ebe6174ca46a79a0f42a16b416;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd12bf5f11f5868a9c40f3efe3d7754031eb8f54fbc7840b17b2b5b4d2317cadcf6161313d22b0b252144a479abf76333b455eee7816ca41ccaef9e6dd49e7f82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf045b5327e8cc6193e3f0d8a0d933c2ba8277aaf0da7b96dc955a6a477f37b50e3f1367c29cdd253d79d7fa50f4e516a3a4520fb81dbb4be79cbbfa298efda2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha5e8648679a0133acbd316872e402a1198b6a8426c7b787b4083c51fc0f80eadf500d94fd539ec74ce22122b84577066c72cbe6528d47b07906553e6d0893af6;
        #1
        $finish();
    end
endmodule
