module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [28:0] src30;
    reg [27:0] src31;
    reg [26:0] src32;
    reg [25:0] src33;
    reg [24:0] src34;
    reg [23:0] src35;
    reg [22:0] src36;
    reg [21:0] src37;
    reg [20:0] src38;
    reg [19:0] src39;
    reg [18:0] src40;
    reg [17:0] src41;
    reg [16:0] src42;
    reg [15:0] src43;
    reg [14:0] src44;
    reg [13:0] src45;
    reg [12:0] src46;
    reg [11:0] src47;
    reg [10:0] src48;
    reg [9:0] src49;
    reg [8:0] src50;
    reg [7:0] src51;
    reg [6:0] src52;
    reg [5:0] src53;
    reg [4:0] src54;
    reg [3:0] src55;
    reg [2:0] src56;
    reg [1:0] src57;
    reg [0:0] src58;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [59:0] srcsum;
    wire [59:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3])<<55) + ((src56[0] + src56[1] + src56[2])<<56) + ((src57[0] + src57[1])<<57) + ((src58[0])<<58);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94fc854d654da0e6d55a961571543158fcc27dfef2654f3b906627ac84c183f9d32336fd65e9db5b4165236aca62a30628abfd875675db165cf0a8738681bcc3f355b90352a0f4060f3924091009efa9d6903fe4b44c3e7db8beca72ae7aa099f890b0dc4c5958ada2f2fc24487a432c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5625eab0b3dad86d4fbcb8a7285f92766bc9aa12e1c9e1fbaee0cee334fad8a3cdb5930c27105a9af6221e94ccf198393f72e6050d7ae2a05e03d24270266f2933199768296ead9f6a47d79f3b0b9b181bbd2e94301120b172ba049299c8d3dfd69076474b35af8ecdcdeba7676ecafc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d285cb3a0c6e968330ea5b153b04e3ef66f2a135be93396b7f1abbccb5273984ac61841aeaf403fec373473a4bda97476f52a54599b12df40314d1b0ae35e067bb7094a05f8170bc00baa09867eb0bf7274ed3df5d841806c76bee50460015b57aa17af0b0f7929802079aed75ae4798;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6423f3d7b25359ca1694086407b9efe06fa5cc60d35e836a8136e1aceca889a1cd162c314ff948aa4136044e169d76b7ac0f23adf92f9146992c3ab38ba1b560d97447c209004063b747cf8a6149dff1edc3efb04c0791f38bff6ed95e54d8a606e1f54f3f72c0169e0f08a2d656848da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h572a541e8bffc0fd3d94315fcfe972422a593647460b901e93bae253098de8bb10e82165a35ef6944d081b19f3729a782c188ae5cd2269654acc4cf6be14642b19f5c80c6a25de37f90e05fc86179420a8f671f2448e44bc0d25a2e80455f2551b66c9671b3d591ba635e1e63642b2b2f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61c24c82c1ffdab8b2a96cb7ad36d45fac9d9e538b644e01c44bd6d3e95702379ba406ee4dc0edc22fe56e26021c4f39f25eb7c643ee1c212ff0ee86b52b02a06ca1e749b46a3d406fa291d128eba9b53285f8e82753db1f480edd67171102d2e4b9ef73e34d786cb0dfff55118aaf5df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aecd0e3317ee4c44379f514e9208ab4fbd2352d850e52071a86b075e4f14241c44c07b3fb4a463f65eec61023d62397a3a968c269c2e65de6c6f9b10f80ea59fc2f6d6ef1869bf4594aa81dd167ac911a3455029fcc0f34244a66408d3b43ff465ced10a60f497b46e1e452fec87aac3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56babeeddf7d33adcebb3654baed6e20abded5bfb69e18a6cdff3c4540573d35ebd08bd4570adce10c7968eac2d0f43484d975e6dbf7c0214d7de4e2682221bacd3c31217e1589b38aea5888bd5cc9d72f28343fb798602e90566e5ab7b65131756fdbb2eda13352c65f4aaa4056ca7ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3f7023eb6ca16c7b3fd879cffb01872a77956565fc44e5a44c633998b2b2273f4dfc6e66fc9d972c7100aa066133cb08a4eece31f2917e3085f09383e4c3392756b7bdbe8bf9581a50e55daba93b28ea4c580ae1e47465b6807ee8cd8623cfbd70e37df93e4896cb431aba73ff63f8d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5d0976dbddd2353e80023a1ac8ee7ae61a62c5128e61f1197e98eccfd75e8eba4c1f279a73863e674086bc06783ab49d803bcf0151f2f91620dbe5674c103f7a1429e04aaee8699a55cc614b45bb93c9c24405b8749b30fefc883198ffa6ff78d31ac359edd7c7f6a35c23675e71e3d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe5886c8586ba401fedd83a0546750f585bfc4951971ca8480274792cac19d2fac03dd8100712c371f4e3a22af59885f15f2c2e72bb2f75b131f4c9e24a6bab1a6c19df352b8de0027541a4e6641d6c6b3e079b7cbb9330f8b4a108cd62973c552a7e0d789f56f33da0f9d6f74882a0d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14d1a8abe5214b23222cc44e12dcb84e4312e167af9823dc0c8f3ccdb379dd15010e5323105147dba93656cfafc397714c60b16bc696da73004126cc1cdf7061815b8cdbc7b99c4ee7752a9638d1fec0ef543e53b6d294e2a3904105b9add04f50ea3a7c843f276a5fa74d83b44f2e677;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd4dbb7e01b7aa23b2e683c7dd21003cf7ae4797c9e5ca4ae8beac0bcd0e88b0996bfbcd3ccdb34c0d01e95e39033dfa6f6b4ebaa0d5c13e3a062e78f50b22bd700940172fa58017465f8d52d972f28ea4ce693c3243dea22bd9f97808ab96baf6b6ee45352d87511554f590095a70b7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55dcfc19eec9a34b34fe085e640bcfaf9feb28a37c41029bdbb6a185e2a3bfe785ee2001deb5495752ea18ce6d011b0c3da72248b594d0bb386c615cc66bc68251040ddfc25d24cd35f0dd9d74c2f4ebf314e1a2d6b4096bcb304e7dc644a13bc46cf13d53a01a3df68222702cce4b7f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b0ac6eca68850b6f694942cb2dc275551f8eb6249f35fbb88090b7cdc67f2ebbed4db321f1f888efbc9a686cb938a30336327066470f6066604d8f29732ca935a32948f7f80b2615de695ab5a3331c71923890116f36f537bc2e1f08c7c22e4d54ae3d6a22e9accb3b850429f86f66c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd6b1150eee8fb45b84b1cefa7122f0798e4b35e8fa71d17f9394edd2c1879ca82665728aae4f24ad9d8e0a82e69193d825c1e7f4024ea95faa9d4a8dc3c2d46c915229c927103ab834318649d01890a418492043ed5588169a3f0a4310f305abab864cc7e16c7f0a1f745617dcac8b94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7be636f75513731a3595feea5259ade1f095000b7f9c778823ef45f2a398b749d2bc965ab33c4ee2c632beb7171a29ce865ec9031f3e1a1da8c4194d4e84869366c3389b9945e804d44c4c26a9355318a50577483e72aff3fedfe4b31754c108e389de4e0c13b52e1dcdb12c3b114d523;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cb870dbe4f4245102bbf01baecfe677aa95009b688ed54e3c420b36edc07c7c9ee85abe652f935af988e8e4770b89bff7d9faac1028dcbb8e1f1141cdfe6ff6f1062f4fdb8a721ac477e1a7f194d49d108da5bb2e76ff7e4a95b54bd1ae0853015b6cfab3fbab6381f9f010853a04392;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedb930d490296bac3c915b51876d760b459e2cb4e0add01af7bdc0c3ce423eaa9d18e0aaf20c4ef1fc29eee6bbad195d8c8033788f7c93ae6121f7b8e1fefb0cde1a87da7329e512cf9c3e5e1f75fbb72bf78e7bc04e5d87b3388bf2435e1417e124682e62a0745ae77d323e582fdc8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fcaf65c070996ec46a1f92e4e6691b78e0d2c5677b57945d80ada741cf763525815913b0eb1793ecc2302a5546e1aaf56dba899cf3c5ed32d92feac359fdaa8df0a9b09a078ee58b92ba3e6b38c4986ae4cd088822b749379b205bce3e90e2f218ddbd975da00ef18074b6095f8ea4bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7014f864cf04a0c9160c81fba04d429c7a24787e4a4723b76c0f387c30d7e4f0853c4f9e074a5afeadf51b91e9b872cd04bb495371daa5f11bd94b8473cddb6221eb0a31e3c7d4c5820599eb1b00a2bb547176edd2d563416f9518d35e66545cc9fd06efc94d8382148dcf182ee5069e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40c9b7b0bacd871125c05410700c96f05b1f1caf0c746e6d859e3322a91db2e3402c1090d2de95d717c3693cedc8160db9ff007d06e507fa854839c131580cb699ff6fa545e6992e21ce8b3f4f93f4dfe418fcf10773f86b8be8ec896d1afd0e9548c5d89e7bfa71e0f74a3f10d7d0ce9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8e66bc095491974cd5a188e241ecb767bd502cb6a44822cbaaaa41164ff6430eabe8bbb3b414cc73b6329e68570e4f7c6009dc2fb778aff78b2cb0d1afea0799a9f7e5fa165459b6a366e2493e24285da55853b69b5fc0d6f4cbdc1231f87d676bcdfa57bce715527b18b00139f93737;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b42a6e42b9cce2b93f9af33bea595016313a04c549d36a016d1d37f0b411d21ce226d8946dc9061f4cfa5fdae8812224e2d7cb1b05f97334f1f4b7ea5e7cfd47a2bb6a6d4448cd440499760301476787d0dba1c3ec443e7c8c75e635ea7c41e3b42b34eac89049dfe7fc732067658077;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2c524c5de34c682ac514c1e5d499bb80ae59100667cda1beec8981ad53a68d473649668e59850141d647c2e8a2f9cb37eda9defb5d6ed7f3df7521cf76dfb60be1f4f845d3fa8f14ce411747961eb2b99f393c92cafad555b12ebb81a9af097e5c188e2effbe72bb037e480b0362cb26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75a44cbc0c2ec7d848fa8ea61a519cec57e20639ad340500d9710caabd4a420d741fd0c33e98e69a0a5700eadebda5fa0915e356572703c4c6a6c1c7c474d30af2050abec83c0513520c62023918aed01541e50ee9b1e6d5fcb96fdde457a6a7b21a7a5a010290a0665b401773909c861;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9386e9fc3cc9d044888d4e6bc5cbd160df11ab1a736e1e6a151525facc1736699adaab50a933a3ca383c42dc927e54b77e3b7bcf16f6ba7b45ae392b5dcce66c709f60ca23f01634bdde7b33ae3cec26ca0bc3648b94838b67f6daa0f1a2aaa48caef8a41e625c607ea178747ee2d461d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1060216bdcd090e5f332e250a77ff77d0852de677a71e522456aa28e83b2b390191679485747ebc01d164c7323283df0cc6ec59bd18ce8b1a904fb0aba4579cea86852e51107a33ef430ab014e968d09823b43c2803be66c9bc974ac9f8909967b60ee4d5b3463b2ff8c31378fc42e5cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d34b7fde61e8121ac983ce4f25d5257829f90a283488b0a6708bcfe17e390ca319bbc40a3e356f5fec6f2cd28900650e10da483c5cd0c4f9518cf3e63c326f030ea442169b98c7f04b58ed1caeb25503ab961da39b4daf57fc5b41ebff2be193c6b352422a826ef5f3d02bf9ef8849df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a7fa5f40f012f43a055556cf795209f614ceaa3fda5a942a627154f74688c92dad456698288880520bab06ae37717f763f248174ccd723563facbd3ae5daf7da86ad8aae2f8458e00ae2fd8084dab8b12935f3691a22c7af10273fd1fddcd8da79d8f2ac3b9c0fb1c52259c2c0dae321;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2adc0867734ff5c5c5d086e4cd309cbd3e1f85c81968efa60ac1732af563a6b2f5025b4dbf8b8edec991ba9db96fed045a4979633ae495502ca038c4a8cf64ef9a7563fe3de424f7d9c2f3294b5f376511a686763e1c8ad98d00667f63f3a6bfeb9ff6834a31dfac556947aee6bf30f98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2764d8fdd231af77437469cbcb67f804ca621f60a2c2702c5672c61ce96c8af309de7c77067ba6c6ac4be83c19d91addf0a160d4e6983e6650dcebac2fada2044cb1846f86fa589f60d5fbc9138f827fa9f0e9117cc9b70df161b67699520bad6c52f35dda7462efb84e60bf06abba68f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf996420de9fef293dfc18cab1a721f3adf5b3fd6710b2a0b27618f0a2b529d7cb1fb5001bf6dda647cbf9904f279c44196f73bffd031689b4ab92eedc57c521ffd76b1005c20290bff909c9b306e3362b36ae681d78b21f9530e54f740c0f0da6343ca077107a46d30ae6b2a6f3bc30ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8180665e46e2debfbec759db186db2820476ed4bd2beddec44eeb674a6be9507475e64da8c5da3965c45a1e54c105f7c30a1e0dfa4eb43ba8016f51c554861cdd8a300a49c25ae0d1d6043865eeee9ef7d86cb391df98b235d10ddb7fa4fd7724c744ddfa7e6e47eb7a9b7607843b4cbd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9caf3c609be341e8dd15211059fddccb89dfcb337d512a5c2ba43699c24ece7ca4a000ef0b8ba7db2b8c3711674404c0de368d093a47e62aa1595a93b52de3520360f87e58c9753451fce7ad44a7db2697294d9743692364917a78608ab32b244070dba4a5dc6272412844bb04e22f881;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc27eca88f2b0407e0c6be6035bfb615ebde255ac2f5665532e1b97e61f91cd1ac2dfba2937f601688e6ebd3747a97b0121787e3fbb11e6029e219db79e637280c9218b1db20c61ecb2223091c4831c7af0f8d8a723a91bcb25eeae0fcc567271aecf7f348cab661009e83666fa1f0492;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf722f1415b9a46ff7fda7291e295b65160fd5b9416f1718c4fefd3d17f6fbe1c0f1230cfac7c1c78e1030b036ce619b765b38f6226d1febc88b6b37c4d35de400d11847a38f115686bf3ca05e7554762ce6934a0304b00f30c3d231ccfd134426b1a1655aeb179f02736a62aa042e1e03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h545464f078d2149f54ebf8033df037bdd9307e53efec64bf3fd4051c00fb7575615d0b6f04ab780eab3ffca78ce907ee552177008904c135e74a415d40865ffab062e4962a9f30fef67ccfa9fe87b801c52b9000a53dd034082ef14f0b420fef6a97b491e95b6234a2b487a6ea1c485d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc7fb8f959b44db82f09e24035afce55cc5a9224b65473e0ab3f56cbe82a517c723d393896e6b2f8c02187712fe59071081173ebe2487fd74b26122a44df601fddceeabab37e33bf8ea488e6bdec59620561fe8e3e9dc07dce6fda9074cf35d98a009b875bbaec46d831f440b9cb4c627;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e1c0bd6cdbcf62a250349f4937ca32a6703a336caf4eb3e53b574469e1a1148c2f2e7a34297a46c27270fbff89ab56bdbe18355c939d6c7bae4aabc274dd89ece1811e423d4a4247ad6187e6c06c6e9cf421eed8331035bb1b9886f23c783a5d7c0ec02ba38e7796378d77a09d81ca5f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78d8a8a68dad0b146f66dc0205a2a748b687e636a83ebda24bcdfc3af1d6972f4617d51ddc43922c75ac0d2be508d08c55b1dd3efd510df7eddef0fb96df44e6d820b960dc3b5c589d8ef48e8040fa760878f6c29762ece0a0186eed72bea04f850366e495a6b034b518a564aefca3a3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca7de8b0206e12fb0e03831ddad0dff42367338b4bce466da1e5f7d5c69503174f2d2575e3ed23627111c83b4243f651e583155c1d43fa8c78d1d95800f05c7d1d68ce8596536eaccf2bf9629c7f3d9a9213cbd55c9bcc8939fba4655dba8f9b8f0d11996a8f4df5786a3ada9d397b42c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97ea065cd4e370e6b8bf04a04df43560972968c95bb2067980e93dffe022c6f40e0b9c4d00a3ef29f247c8966407a68e437c8cc4159f36c154fc29d2c9ce85635d9f811d73cd462ed048c9bb03e8007e33b61fc8c802ea3eccac07c3acec7a8d27714fbb902bc07878f08788229a5c565;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e5ba15d1f3936f93649dc9ab5961f1ceff9dec5bd02346df4a9908e20bacc2ccf7a8cc2efd5667a6e17335305ab79ffbc2da954b77600e856b541ba352c834b56fda6a7bcdb76c54db57fa54833f0c3e176a8c7869399838d7bd88b22eb1b9a8008eabac1b823435a3242867cc3b6347;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8904b304a15575e4aa545791fb9a98734aff2a427f0c2b36c55eacb3999c9e1aac3b1df5e5c09633ba8e16dfbd2449b427c2f4e2058aa5134174ca9b3afa0c16575e87af4590a3d6e286cc0ae9e1828971f7566e0ca1c09e74bebef672f3277362187d86d3e3069e29709006959e61401;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4239f319116ffda43c474f259df3847eab283163637c914e1316689a8c5581794d488133ab70f152b5174eaed60419fd694d8854ecfb5a4845df74fe7aa6f1e8c21db8ae2012b19f8c3a8ac43dcc57ceda9e3568255552d7fc369d02eb67793eca5f2f4234d3ff0fb2e1804cf522260d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28c6192d197ee3fcc69997a7af9eb84129bbc4171db9bd036958fc8963130b3f375b9e5620752a19c68316e0c0ad15dcdba0f62703dbb695da6bc95e3353300b77c446d025851416bceae9a12ba037d7f6d3fa9caffc01b203b53bbf35aa3b9bd23d403bc815a611d9d1fdc5c5c745ae7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc0a8f0efcda6e7026a6c75cb8e731e5cce8f894c086df325f26919f61289c77cc8ce7f40f45f2f9d9891601a3d0cea9d472dc4b28941cc06162937d04993bec71e9f1ef7cd4bf51d0057f4e8dc361368be4c3b1d909cfcfeba3d820987a58cf89d3d3848d416ea3af2cd867b01bf210d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0882dd043f4bd9b9d12855862bb9f97f59b215cfbbf1b29d0de3bc93a1be274b6f4b44cff934a4cb320add3952659528cfa642f332b142c7c3d089f4a5442806663f31fee71666ccc4be4367690e9d434d176247ce71ce162fbfd1c6474d8e7c9ab13ee9c959c0b586547d2bfa0e9f19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57e2d92084a6545024e58a9e58bc088c9b97e5b54b9d98cee38686829e9bc1a51f573d7fa298c2f3b31c37a5543f53a84f007f463cd4c2eb369f125603d518883cd398d7722fd4861f7b710b2cba4837e65192ccdebcbc6b95b9351867136716b278d3b2920c469dee91a6a92ca305eef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca6974d2ad1d923db9b29383b3e5cc8a5be08b99b1a360f6d2bcc41236b09924273c5d5b770e384ad5a9b01a5b2033696b42e48985a7782389feff55f2abf45737fbe7be12468d18cd4ddaf57c9114a7cf7bdfc322d5a06bdcf8813ca4114f8025100f0fe79b80f6122f41480c20b2d11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h474a6a1a7dd7710f5e4d0d510038e3d8dc4fdd24f5643de9781b1e80a34f12c8e4b989d6ab78fc82029e96c4a0376484a6755f0b11e0088b9b475fc3a64ba09d95359aa1e89cee174fbbbb48c2df726cecce12fc99f4908a692c3a8ee3cfd6c7f723242281b99c12ab844646832097c3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e37054100a85226d1237b47f975efb9821eadf4853495f1758a6cc5607346dca8373ed28c9cb28f2dbbecbfaff4e029354b293519f1977014881a83eef2ed10f38b44cc36e34e96ef87faaa180cd75aec6e4e26b601eb510467899f901342a80427056b979c58f6765e2e63074f1d115;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fd3f831d4448afa2572930ffc1de2cc34d6d571e4231ed22b91c274235debcd71b680ab565e87e92be5659d9f32c44ea60a2c35ebeea18ad05fb59c1699750f9671a7e22feae8b52aa5eafd887f974a3db06c71dd1e1de501c6b0d7e168e3a0bf09ff1c528a59e13ec951318532f5d6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56131f21ee61ec2bc2b9940ede7da8e349369cf41ff77a24d0ed1743b7e87eb8dcbfbaa1ef028f2005dc307dd143418b656090a031a9af5c8c2c92c7954ac4b648be90927d217be1d45db3a5a70ce45cc0a60f4ddc4cb90e159e9917d184eff1ad4a0026ab7675909f4ef8156dcbbfd82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaa7d2aad2ed02854abefa21945f08c51a108c4637cadc086da89c4ca2fdda7838361f591cac5e1b8ec5e35edab294dbf00dc36324f1fd34ef8a8395d78567e96d88b077db2c1947eebd545e196f3158d2d613d4d83c83e99fd0136a8b03e9dc1f0e675185ad6e965ca114ef13e9d8eca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a51cec6bf81b2bb5cf2f77a3deb31f942f98ad38b06dbeecd1da3f7daff83669101b2d8a080667fb398cabe58142f87041df445d26640c5c3546f2d00419a1fedef9ff6cf9630d2b714e89a057ad2cf3bcf8d7db6a7b2683f6740828e00784f02853cae42cec62e9b1ef87d96f16fc52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2e55daf7855ac0079914a600972e23ab3e31b5702f4f6902350b4295b2490cfab14cf91c8ea9c98b13f39e26e46218992aac072a046cde2a82f43a5725b78e3fd7ba4cff27bb8890bb00b6267414a6af5aeaaf39f9323b9722683020bcb4a2f3806c0aed5b4e5b3b2932f50f6b6d1d62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e0097e96887e7c7315284b0190a56f1999da31b5c2802ebff0b72f80e9d19eeccfa5a11632a01e323e529bce4aaa040580d51b6c0b52c7fd5b2ed74c627da3280a0e6865dfdbb264c91b6127cc1c3edb1ad01d7dd06bc718d8c12aa50049bf13ad8f980594cbe73bd996e71a885692d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c0a78e9b0c03f2a71f045ffa40158ed6525c6778746236a1a0b0286536c3926fc29a7ac8835b2f3edbacd26bb77711c8a7d9ac2f6cc0bd33014df9abe5e29330b740049268ca674eef5b3607b5f3850a6689ff2caa1651fc9c2f4f0066104133c7a98cd793c43e6edfeee0a27472e832;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd966b9d57cd67f323746194cc606a6e309f3c8f6a50481f692804796865b75392c4a8e4e5f9c8b06717fd617c2d51032c5dfafb23a17d480ed7f86feb975356b819bf9eb6fc478885398d8d0f43922b07a1eb381fc4bac8b8076a17cc32f74316e8b453f99fdb7a56f322af157c53b702;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50df9755028d24dd6e4414c48cbe807ed0625f4c1e967758ef1a13e0799ebe1997b51c33b0199f9f3c766eab97312386708ac57614aaa1bfec7b824cec16a2549502af0eed54c99c9d969cf4253b127e7213a69894d5c73a9174d3e1d29af87a01ed995d3113d36fecdc4bd384bfe9371;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c492997a43dbe68a47be576def3142656bfa4dc2c0fea8951a035027f067d95285708ae5b0f9fe18ded25ab1f7a2afd172255633ccdadad20ddf88b1515b159ad814b447624a45c672b99dbf1bfc6bcde314aebfbaafc46daf8d2de86e45b852cf06e0d28cc75a0fc5ea5726dd3751be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d75800c212f2e1cd4208da5a18a6e42d26fbb7d306f51ed4bad0438b15ec976c7c8c2a6cd9b1abe04cc1c79f33d492723a81231cae0d997ce68658f11326686f770137acccec6306ad8f46892ddf0b49d3ba05c59d52641ba49aa9305f9dfb2c8fcf95058cdbb6cd37b25da55aadb8db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50ad32f9ec0a02d3bf3b63d19df61540434bb60ac93fbed0c0e7689854c57cba17ae7cad0c02e5123d850764ee21bc58732e47479ee7622042b68317679d37806d2f7657f8158514015847bcbc2d11baadd2327c184457f753b5559ec0b2b2b90dbe7b6e6ead3cf521354f566173370c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b24f15c44e71c4e538c3b85fae5292b42cd7b6e1e94510499c377a202441c57914903557c5621d174a2a368a103003a5100a5f84d1736e0aeef3951f688b1ed45b4d0fab5ac36f6460a12b67635a0bec5ab67913e97d6f1080ae83aa58abc7bc678ba66754b995ec41be041583358984;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaf3fc75c234848d9894f41af1352875e40bd4bef72b12d5de2ed44efa17ae23030f13240aab57e9293ef1cfb8e821fa1dd497c0d4dc1ad4c3a58de8fd605f51242bac7c19b96d8dd0d542e7bf08a833f7d1d1ca1fe48acb2951ed540e42cdde11b501bca66b048413e47c3d27601f79a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda055f1d0468c2cc66ce995d210cecd548a7ca4383c2bdfb0764eba444cb019d8cecbf060aff66ecbc284a123099d13c9714cfef2c7dba73056e4c04b86d6888bb437af0cd2ac3c4119aa0d771d124147abf1e91f8b40c6396d133eb400f64d4c18cc6657e146ff57fbc913977256c1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9b171b9f1e819e12eeda559b166447b46d425639b12fe271751b03e936ba1ba76a40b030b6e7a82c0d7bff658e5412ba05f2836998dff3fe78476f6f767cf93ac2839273804a7450d46fc55f823ac8b7703edd65d85e18764e8fe985c07546c1423a89dd9fde5d203e388c226da598b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd579185ecf61fae8b73e7bd3cc8bd49a7474cf9501ac21f7c70aacb76bf3f4bc7fa4a3a4a9936eddb9b16590a9b98ffa8f5ad4f7862ae6d6d0b4153ae0ffdd58729366d6df41e72b660724814983b672e9e70ebbe53357da0b0cceb1e5adcfdf91de6bbdb9c0df1ba26db783746ea4b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c9a0960216862b0709165efd896b0ae098cd419562458505418271d11f7f312bfc75a3947e81e62979fa047a484d8c3e11decf52392bbabe08a7255ffdf3461c93e2f8ce3f41d82a38cafe76c7e80220e170daa83a5fe100ed55f40adbaac44cbd5e7573ca6baf02e3d232b73f4f0e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9906f6cb0c4eb25f394adad49e6fbb01a371f39698d5fe47ef433b02174a8a6aff8affdb8942b80688810db14a56000d996aae579f5e3f6631fc4bd19b8de5fd82ff758a428844d2348d9a1f940af75267e1c65679c0bcd865e0cb3ededbf2c2773c0541e015a0b76bd5273a1804cb093;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bd801fa13c968564dcd8fc93b7e156e75e352ff9041f17c94a36ba3a145e7da35081f03ce99081471a08e9230a64501c859a6c829126e136e32147906f03cef539ae61761a4d17ea936fc3921fc33bb78cc75fb54e1a45073309e39e82bc870497f74084d1098383e64994b2c3f5c785;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5209a81b233ca231d005c8abfb95d69e7f4d9ca4b3571aa9381460ed7e8164312cc060f54dbd6c737fb7d00e43085e7dc145262d6f13c6ad7584719f61ec3186c5a287debedaaea9184a798bd9b89923939de36ee13a619ce981768ded66470ed4ae0073b37e4d74b3790b1aa5d1dde37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e563109c4246ea5798382b5adef6dc9760cd058f3f3a6b915e862af6ab0597e97397ece221718a4ebed4ba6c79acdd6f0c08070a94a0ff596dc521f869678ce3e419489ead8615a7e2e55c610308ba92ed5d8bb42a0eab9038d0cb288bb84c316ff20d5effc2f9a09e0f8338d01f636e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3e321e7649edb0fc87c931bd2d23d9d782888bbc1ab3619b804cee08fd09a6bce82ae7b5bba9865428696b3ae3b9fe92f58940b6dbba1b5dc22364adc07d14e179a1e6d219fa9a44bc1a6a2d0a8736ed634f63ed0a820e7bc59341b11c6b2ef6730f0230107537f64934a32cd75742c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ce002228e41d2e4057593a0486a9844fe88a23eaf87a9305f020fa5510dfa09c3944f68b4beabf323e3d924a89299a1ab5cad418cf64a0e931a6fe378a5c01422a1eb39dd0db0ec91cbf99bb01307e817ca8c2ed4ec8f5cad118260e9943cdca66cbae538d357a211317a13a89a423df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h731dada87b5bca7c4795f339f37bbacd3568f8448cc899ed6f9dc492e22230d7b48c347f5873f93d806851f7db29835c94c8cdce0697807729186a9aedb0a84dbef40f8113a0ac674b8d1d50061b1ff05e6136b865770cf6ef1c87e03ec92ddc23a88e664bc2003ebe2dda7e404acc111;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40dd517c13a77ac6775c2400f2345c35ab14bfc53d3784cc174814cf64cd2f06f10b76431f41b8b1753ea66f9060c2a18dc2aadccbf19ea8f1accdd158002ef3e708fe79358b0e484c2c0d07c3c2999181ba59013c7adb62a1719474339085293718093b606ecb74476a293265e307a37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbad4ca6484b2373f52b5a81c4cad04aab33fc8213cc21d5f64a87efa49acf5e136fcfd758c0a774c109f9434a13fb9b8f72a822f778f43533157a209dd653416f3ba6d60a6449a7b73d9d170e642a5a2cb775a2bbe908b664d8fb003f86dabb6d28b408aeeda7154d6a2e0b40510ffce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc195ca05a1003194f851ebc1d040c0478fbf03a1a92e0e06c73261357c5450e3c283739b30dd34c4789e266bb8cdaaf1d274f14ba1c4c6d5807e19f25515354010a6d12c679e36d3ffb965eef6dc0feaf63bfdb80daa66a5ab7a2429d084c5ae06b735bd2daeb8509719e27c8b92fdc0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38fc2dd77f6336fb70eb8919efaa5d13c99077d21be6fc928dec8345cadacef43e554ad2e8068e65dc407bafeb3ddd5dd6e0886bd8ee72f2611968d90bbbbd59e96ba5a18d81ddfc66c7d4c9f01456fe02d3b05f01956abc4341c469dae1b4f811a42e23b30d399d1b48e25d2019dacd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61b39b29e4c9f7d66cd6b3d08f476c3ebf2bcdf641e962a8e8c7bce4ea42e73b52678a1cf6be126a18916a061a5eb32983e78c54a6a51f76179463f01664d264828c221ff5493998396d96e29f3916c49626ecb4e0ce50a57ba52c1ffec3f5dc8e762f45bd81246130e077c5f6fd644ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec9798834ee632d8ac2e6d94d1e0934b101beb17653756f54f6a9c20208861b6d88943c72fc5b4264c7fb9425f9094f4fc96a6d5a8a5cde8cde689ca7b04a1bb2950a09321ae25234dca860892486614c33b88bd901740ebc7179c26e07507efd97a19d9819c7dbd59a4e99e89e5935ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h266952818e3d49ef6a764715552c0331a6b932caa69682a7b3f9063c266411ab01253c1acaa83e7b52d3186b246033a884f0fb1dc049f9b319d2a720d08bd6f3f547245b25e3520a6ae620f254deafbc1520f7a0e07203a18955a680930d40adb72b441f09f5ccbcee6b02a2cc423b241;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0e75df189b02d8a7581c5172ef1ef41ca703c76c8f4ce06af92d7d2fd9b0205231491a0610396225a27805043c731994e3dc4c29ad3efdbe412459caa2dd1fd04ff31097702d666a1c4672c59104836f2c1ddc3a804dde4cb79c08bc78a2bff9f8231ce2dfcbd4cf20b181fc918f6095;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d9ab432da3dd8dfac307674948259f9f9a1a5e6ddeeac162f34c5d5194f1e95bdb77837eb385053ab466ee320ce0c4dfcd4c9e5321d792424510a94baca81548521dc2879a4d8d8c7db298419d61d24905e71d0d4f10ef552625ef949b0eece778bd823370b9587be07b88eec8035daf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he22d0142dd67bbadf9acec8b5b419f601f8b2071e42c6e908d9856c1d886c3aef43d0a816477ce5663a37d5269e153e74b24130460bd462588ffc9eadc9cc3a8e97ffbea84f1f72f27d6fc387f9eb571a99a0d89c929a792de3b0f7a758b4954989cf8bf0499e2c800feb7d0aa5d348c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha24356bd00e70e4237d414583aee1ee8d5590eed979c4186da7cf2ba9548705b6819eee7fc6c12d455e00c56317df8025f10e68e30f126121f7e9b5e69dd019ebfa19ef0ec2c495ff97e1746e7eeb54434b0d4f243c95cd2a2e3cfaa8615c740fd636e691232b5fc72a7aa47563db8652;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43d96edb22df198b7eee6823f19da5d13d2ebb03ffdaead5e1907191699792ea4c5f2347d5975b6238d32b766ff1a4f69758b44178d05da181c159f0351f6e908c361266c620e9629f8863c5e54aeed96196d5b17f1a39063eef8698d7b4e15efdc3e8f6090bd93798351986487aaa93e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18a491ffd678e42bbd09a4c0eec91c6634142fd3752823104e2bb124b658bcc8f597275aca9cee16bcaeb07648f9f363ea2a7a5837460c2edfad132279e41aa7b2fc71b651e07aabcf26686e3be6c0552f3a9a8aefb0695ae8bf72dd898362889ce4724cd2290936a3668ff9c5232640;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h299f516e20ce8314b28315b82ea7b2199c14ca66bc3354ccc90fe4f9ccaeabf0032901233b7ffc94ade324891d565d714e4313a7e5b841a8d2bb3ffe68a66479d75e750e0fe741a047fb2b98196457bb172a123b0d9948087d33d551c2b6bf6b475a584cf2e60c5530960a3aa50acead;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12fcba8b56c93ba52dd2cb1b72fb21392f16c2855159cf753296bf55f0db26ce8d3c3e2e00ab6358affeb9cd512260940f8e578ad3c750bc3b0496a9bcb2f6c4882d0d5c1b98941a61462b86053bc2a9994ffc89ceaec7ab14146eee433be9d16916e51ba19af48e426a1b3fb867eb852;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9c6a7d652dee7cbf7ddde4e2380a8e05d1c8c9fd98a9bf6fca127fe41f6c4f809181a018a2cb958555aabcaaa9b86ecf2ef1d65aa189e9aa8e0bcfdc51b1f37fcdb80ea463a4ebfd887bcef3835914afe0551a8ac4b38bbe68dee63f7c0bffdd0e736c92c5627915bbdbb3a984ab4b20;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ee0b208da81445025beb8f8177340d5b121acad6b2127291e48527ca914a1f81253b63d616988bdb0afa624baf9043c9680a3e4c78720837513a36a013d551dcbeeab2cddb197a000d47771252968ba2f7bcab2a45d48afbfd8bd99c6522c5cbd6a5e0da4b2b6f4018613e721ee4092f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ed5cffc3c669c70bd7ecd6fcc2363d5ffc63aa8ea7581c46810ccd21bec7e20732054e19d9f74bfea4ea881a5a273638f8d94421f0469070a1b0c91450cec1bd750630f7d627bd53c3ce0c4b3fd75332c53f2642a702095248ffd8a93d59715141099a1daadf82c02fc6382f3ec6b02a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4b91d554f4392a230f4e041b5cd7d6c646d0e10f46417dcb501e83587a1338632563594777123b6fbf5b2b7d267040f7005f10447cd31783d272bedaee3a895983096f36b4c984ac691b7b72d74143a9cf37ba18db52e49cc39c4403ec71a7e5fc8a470cf03551d7b5f12d36c666604e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6b11de6dff98931a7e885c84e86226a5bd8850a64b7c53c1b87af6ae0f5d2569afaa217e16c1ec7ba94d2d2f4d4f5937e7e011cb3e9444fe1fadc928a48cf34c75c43494f045e429a3a02b7be4bbb8d946025f80a95a80553450539455f154cf3b8adcca3de5a3f7f885758268d6f1ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77267d92940f15f5c1c49f87cb0df87812ba6ece64f0a0c46110fd3dd08f1160ffc2006ab57f571530cd28af7e719a9ed16d720d249b3a32d985e1b082238201c7d0bf4c78a510e30500b25636e548f2a31e6f7cd0d4bad74e3cdb4bf08fd64c86b15f2301a39037f75417929ce062a56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2602c4a9eb066c8bddb02a57b6abec049ff2891b4c77dd2beab91a3664e1a7e16259806368cad85f32da27579f9f95f5d7bae487bf23062266f77d8f17d62bc0a4db5b25fc036a1978dc1e7f125ed226f34fc04178070491d8feb76490846b7c748fc00f2a55216e50b611eb2f1e8b5e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha19e560e49b892cbb09fe781277de287a2d893e825cbdc827f26668ada95c10e59adba10cdc4ceab7ce8990959ffd02da7dd9c802fbc08241c204174857007fd20f539cc8619a7e86db9df677dfbc13d9a316164d41695320a059dad6ebfd132b4045674350949a6f20ceee8caac067cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd54c36aab04a99b457e0568542e4b3d677bb8c3062da03d80fdf5871ed9a6524abce707af4146a3e0a142cc19dbf957dec0e3329a5d8f2a449c017da94059f3bfd3fb77d1ccfa7717381520987fe30e26ef466600f391d4e4045a4b97f077dd5ac8935382b200b8811b8e0a5ad30384a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcd45fc56345a0d963e95dda1b8e8073e3f7f355111dbc44e7c38baee8de7b52ca4640a6ed2c8a2d0c553f753c0f2b4ed6eb813e24e42200bce0530ed72fe6bd0025bbf863f1f0ae37b439421a156938b2eb36323b43e58aaec18c0ada9f1a921ff3fd691f1a835c08356b98fa423517a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc1034b92ad43a739fb21941ed205d76127920558944db2d3b64ea0bd09cc7c6f64ca3d27eb5ab9779cb3e653a22bd810688434e95525f5eac90770c29ae9a4be02f39b47b76b9c2c38253068268ea9ee6b8adea8b198dbc0919013db92f442d14cb5fa5391d8e9e98e3fe9ecb1309f31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98c185cb4c794451edfb2f06a6b25db4218fe282299c1575fc86f3bc2890d07d7b4ec7b89a9f1e096549011f4fba988fcb27bc4b09e0150aa262b84c160c8a3bb4813abdb4574efc7ad1751b541877b5d5819db8784513952784e440d5dc4b6be44c87176f072960e171230574930c0dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdccbae527c9dd571838a9a67edb75f93de62fba45d7793b6f1a7947ef6c0fc61a8dfafaf4df63b219abb2b85b40ad18800f31ad49216ea893bfb33e7ff8027c69896fed75d1caa1bbe40a1e19e5d002af56ebe1fb0a36fead105c926aa21409569f0cb0884fb7fd6889eb6759dd667b89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14890eae1d28ec63a72edb2ff44e01096fdbeb8e836eec58c3cc8308f2f919a617c891a1e2211fe926a736184e4a67e9add0d201b71b02522ce01f3a991d736acf5aa2aef8b44cff262e955f9bedd963544926c4f9b92f828129a25d6a8b5a343ee57d8b37a20649c393d33c55bd0473;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde40e0f179b883a89dab9eaf7475529409f51268a5a76185f23d48961df3e8076c4193d937800f286a9bb0086893363fa39765dabe2f0b2359f6476d9c8ba06183eaa64b8f75b929e33e881fa188980f97ec361d36a8904bf61e6c48fb9c9c8874ec985f241263215a105d207d571f9e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbec03f06c9ebe23ef60bc7740b232e9f2dbf2cfcb5009e111c9bf84e61a81e084b0197e7f2420b50609f30c443b886ceae77890b398d2da59b0ea6774117e1fe3da5e4feb9c246872c35c4d810e4e1ef12dece0232a5d034311c7df3c095098c826dd268e8ce0ff98a4f12a271f984497;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he226a9f8b437855a5cb44c5ccb859228ce757da1152e171b183c4802a6b14127fd6d7de1d6c07c45aec2400391d4985c8d43e5866bce34d304db59191d87fe5ededb60526fdf715789a492b4823e9a9f0d674556010b68911b006afe1b4db5284413c2245a209a4477f35916dda54e083;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2fcf3a653de3e019f49d5471df4ff8f63fac3f036821d39a07e45bd2c9deb2579f5921564d79a433ac981ff705c6c2ec182a70c58e0274bd90f160345c99a99bc31f633e517cbfc79efad385f8dfb0527a9cd53e2df560125b61d1d9e55f98ad8d0d2abd19b4e9641a8222d154b05950;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h965d085560a968272033519c1eb4be399931d6c6f3887f72eb21a2617d7138a9803b7052c3c26692f1e47516b6a507ca4e8dc6d2e7f5f7805f33b8541c3d53b62471840e55a1015fd203c60e27203eaf8fcf47b36076a0dfdfb8e64c1f8962004bd5fea3d17049dcc007f2a5fad8e3f46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ed4fe2db1785c67cc790105133f668a3ed2a4c92f24e023a8c8ebe40e3f0650a065e16849e7f16405f6669fff2749e3e852a24a55029ddce662a2a75f5082eb00eaa0847655f961e3649aab858b9ad148108d1e71b026df68e2c8a59324798c6350990e718a15e1c5c8fa66f034e0c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc16a98d5ea1de890b41d19a796bfae773e76af0c4f654f19e22bcc3e27d76b5b2da0d3e02ab49929dced04502e303481fc58b421d1b655463a869b83772d054135005011a9b75045d8fdebc0510545ce4ad309e1a731cb1fd37ce4b389656650685d4c84b3d4aa0a3b9e4ea7cc1e93fe0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h144eb13641fd346bf1e1d5868b6d25fcc376e5f501ba25e2da58fdbd1724ddcdbc01c289dfe8be1ea5b18152088e3a9df3265ea6879411d1a2960262ba0032acb6d218354071e361ea91a4bbc2966ac1a758c0de5a6b9f1172e80cdbb3782b650fc4c104385ac2a719dc90678f0857de5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48655fca2894cf9b60847d224fc600d80f51386938b6769f30491c3d9d0852631e761b2404c22ea874814eb4c138118ff895caefc2e989f41dccc6f31a5d93ae7843e05123f263a9797b5f96154fe5909d7daeb14bc3dd4be394b8c1ef515ee750a8d1ae203d3e2997bd196b879a6ecf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9fbcd1ee57f32cac0ac4cfaf96c718c727b9a5b961176531a0f42edd5990d2ce1c979c6c38eac8fcb933d7edac1cfb8fc9a232469001601801c02448243525f0f83dfd50e5437ae572c2ea2b9fb3065b796fab0675d765d84e3e3bac5662564f0a5119956c83571fa741c85879e95b0a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b0cdf586a48739d5cf7208454c21deb64f6dfe7887a17eb1e5e2cabcf6821de37b5965e9570ce7ae7787df8344aade490118934320ebea26e92c46925e56dd8a4b0e947f6d112cbe34845fd5ba2fa1f79e0b7f73d5d7a51006a71ccf20cc8d91f7aab9a9e78a70ae2ee3b20874b6e988;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8fe942af285f873c630342108b38fb1d680934f561df4af63e8d2f69794a3dd793ccfe6f9b395e0295fdedd0b4a2fada7ba8e881c1312d53d74242690bf09e739905ed60f67c2c737104e9a1d2b8411e48e6dd48b5eb2e05da6ee1b4e734b9e15ba687f1261a572b5481c4afd75753db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3c4270c306bc9fa001f029daeb068ae8ec4b8a2474209f4cc7d52d1ba377be1965349e7b02f0cc00956bcc85affad3bf61c6496642a33fdbeaccb5aa9dbac1831e6e4b43732ca6e093677428cd974e1a6451ceaf1a2cd910a1bbb087ed0f2ba9586ee268d79efd845563ef154f519664;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f814386254578b76a8c824dd68723ad319d390b761c6ab7099421ed89bc2f3f73e46c6ecd0b09805f849ef52414ce79d49b5f4af04f4d10fd2dc0a8bc0d31fb8af18fc3a41af4f1242bf04a3798b2ed873ea36ebec6a2e6a57a9297a35d71dfda39fd0116782308e7a860cde707a9010;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd31ac9b13dbf8689d6801c0e65cc5744d93b92dfee5b4ceec8538a64b158ddcd653a076610b1d116eee9bb79c82aa2920ac27c39fa3abd5e280f732dabc91030a8213f51ebfead7c55b8c622daf4a8743e473e91354101cfca3ea37fe476438be628b258cd70fa194ed410624311584aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8bd2a9e347d8cd20b728bb19b7d118a7c7925a18162e63634e5322ef2baa76d7065e917edb22a108c147b19cc1b13787aa42a48096aed765ca27dadb87c6a22f99a981993ccd5be472705f7185acfb5355031be504ff0fc04da32fb34bfebe9ae78a841a4744835682ea272834533ce0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2467d04f259797c37fda5b61e9dcf4cc0631f9501e7039155abd049e238bc9e1ddab0a0c73bcd61c0b6932ffa95bb4d4203fad6c50909900098f0c36706fd3d12c612ef5ab44cfa49650acba6e31af794a797833856f1195b0d4465903eaa172ed4753565569663312d646365d66064a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf19dace4e4fd2a0fce2e978119b3a615b04b54620b9886c552aa64a8e35e1c747f301a548ea42f3b1ff32b8a0ecf292fc1811f3894857840a0eaefa57d030b84313e9afd3a81abbf877b5697cb327be24e2a2f0b14193665d0b02937d3ada4904072409d476c5cc9083043186137b06e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h547bbad5f99b11bf05ffaa17b3a9afb79347903c7d9c68d5e312ddfb61f5f5e50cc59e0a965d28348f9bb61993778371d327133e3384ba8ff9288a32bd9769e920ab2a903d980863c90d0554255a85533e88718322b042eaca2359078b2f19919784555b30157936479f72a4e5f8b61fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75de070a0ae2938778d282a4d3de3d2edc8192a1132b2cda0d23146e479d90c724f27766654cd34e66ef1800b6bdb78a4406db656080bb5ce5dfd861f081a6369b03b2180751f42734115f5f60cec710c7958fbabd39523b5fb13136b9c9e290a6a9129d762cf77ce77dbdd986df91b2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb47b60effa6fda26ba913ee1eb64d33ea69f664405bf85227361e93780abff4ffeebacaa326b4d431c7edb2b46188c3efc45cbfffa465a10003ff97a2255b43aec7df44d16476cff01569a556dd4a86693396a7ca670adbac006b82f3ac77ace9477e2d2030c5ac44ce5d30cb4e91e90;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h437b394f3f688916a7ba524f234ee200e0d3cf4dc9d6e342031b7b9b2f236d4588e4d8b0b328b205b3115a146b5676f32579824c94077744c612a42fe70b2352eadfb316fb7f6e0b739549a7992cdb9e9b4217655a8169d112edb0b371e7a5e3482ab9e505cb3d9fc219933478f19b7e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57ac2166d4fdf640a06100aea1b9291716383792afbc1544573a07da423d40e95ee8ca62c934ac522b163fad5696d1d8484ed3251593e9d6dff4e922fbd6e4f6df1ce9a163b082fb55c8da31e22ce58b385610bacf20e2d660ab1d5aa113c3ebbaca7d787112fa05383a651fc9303c4e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b74a52fdaaee41bb4cac82a8ed4c16a608d657076ce108489f77674fd0df5b3fafda577f34082a30ee7b464d31a5b48705bad66faabfae4cc55d0ea661766d1826627a4e2b8478645f2ce000232121aa468d8d35dc9c3dd9a2093ee5fb20484521673c31c258e10c532722504f9f9df6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51f36873ab8f5e37b431b65d3e708760dff251faaf27ce49d8d51d79aa245da39181a32197be6af28e65ae8bb8076bc1f2ccf9aa297a2f5441bf79341736574bcf455b49f4853f61bb37a8a07811883931c132d3cd877242ba3e40ab9f768b893781f5168f572405342679d2f6fad178f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h767a6d5ff349cf7dcfe5644ec569227c2019f25ec8b9cd1a16595418868a05ddfaf95dc40c54715d9927c381846ec62a999271a5f3f93af4945853d2b51dac5882d0ff928906c386b01ef65ad4423756ae1f5a641d1f0a4a3cc9f1ce73529c1d8d714277fa31b6b0cc79588858125912b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffefd5aa584b734ad36454074e5ee7b27185f61cda20fccca586bcb56e808cf7a723dc34df9aa6f6b7bcdd3733d108e73b0c8973196ca27d3d4ec9c7f86881b8fd8ba344f4f7aec1f4a5c2e0406112ef537c4b772b44b287eb0118698aa69ca3fcbdcd5ff1d6b1b16882a2a2ba131f868;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68969ffcef4c7d85e3d896c4743951bcc2770fe991cd54f30e59c5baa539cecb717ac55707888411f5cd607f92886e902662a9eb16632a4822ead8e039cce3acae97b38bf30652f1157a3e2b0724dc96a553a5ffcfad1d5abe55d93e1246a5243b2c44f73a128b8d0f241dac843cbe9b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85faaaebeffbbd12899f40c6cfe8e5b13a8e048279496d47bcb7fd1b8947d45a81825f158180f4f4f231b0ddbabd8e2577fa1f5b65153843ca18f980c17c8bbb4d71859560e703b0835f7bba875f3a4513ecded5311e782bcbb5e2a7b59c8c59aff5512be64bbda92a1a3468dfccb2777;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2750232746a63e979ceec6d69b970b44f9ab3b51538dbb62e677d287155ea73d2865a3177e9c562e3ad6ff3f9fec9be76d5b279755ab4e6c9379efd8a2faa06f33913aa8446a99b2810b4ac846336683105eaf6f329f9b0c62de796ca81c58b10ebfc464f430e575472cc00020865d4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3478c4481a401776043ac063515b6dab3068a23dfc2bb3b820d9b458bfc18ed98cdeb2d2a6ffa0eb14b63a1142c2192118eac909430f297d080832c8e125ab855fcafe9b8d1fc2d69e868c6f111b600b6763f279a01d2870882822a1870213f3c199a3189802b7069b044155a7cce13a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5aad02e103db7fb78ab8a6c094fa47e1676526a2b6d4d68d127ef93315af59870a12b80361f1b1d3fb961626cd8074963c46d8955bc758178057d5ae817a45d8c5ffbe4ad9e6163ca2a5de39fe6aef15ada903350944937805a9113553d9d91ceaa4ebfa6bce7e3b5b7166c6db7239fae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc70a5eb1367f6d826d1d73abe7202c42068ab37c2fd5470e0c8c3389ba6757fb4cf13d1b581bca30f014bd8e37da8ec32c3f461753dcfd3b7dfa7a7b8ed4856534d06172d213a9fcc3c7bf9fc294badb263de7f23ab1d9acd6a783f9cfa6d248addef57cf2afdf2e978936948dc4f8839;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6922ac5d184281e42e0c81e1d036d5a97a9d3b7444c373d8801299401e4721469871c6fe0ec77473620be594190fa429243d9426c0a9584c3aa6a1b925748e2ab9799d6bd64f99ffd30f3d7d4afd5878b72a81dc1108e83ba47e1c80b4ba7c92a5e76221fe64c24e25325ad9f9763e84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4377ac700cc090f570f9a50e354e7f968b755b6ead382633b82632b488c0dd7f117315b3a40b2d7e0bc5f69feecf1d06189c84cee6ea872502262774afef89167627d3af37fa3775ef7930277335108cb060f7073080aad087b67e51e2e121f7cacb3c0e864a96622f11f71a4b1120784;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65f67b4d5f9cf8dc79b4f1dd4c6bcb687a2d83eb455c0209db5c172e05fcb29750e4e9c5ab0070414b6d7776a4150b93a096cbc6712e0e947cb0c6ad5ab965280d213e56e1404d8050f0704028e9878a0281e783f2cecd187050a36b73c91522390e62fb46fe0b8cd798704406bfdb6d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3b6a6a272ec392c596b1ab1ae71e7d127e3db52d043a6ff0ba957165190b9631dd96c8c4415189cc223b38b7aa94abfcf9cc281528637aa956fc20d3b53cd4648b741c8009302fc78002f51174d2a2a734624f1cfe0aed7397038eabe3dccaaac563904fc67eb9e3a1572854aa70412e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59d5da0f8397da412c440a4351b69fc823c561697d113ba354e613ea42ecaee8e578494c5dfca780a81dfe208412affb1d471791e305b8522f9118fd843859b85bc29cd5b44fcf5c782f84f594c8791ce7e0dcc85bb85caf6ad9a38606377d604d281860ae6de751646882d1c2e92cfc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b3c4700bffe6e22cb85df1ccfea27d3ef89d6b42f920924a0246ba9934c0b52279b82822852cf6dbf84fb8dbd1ff3b93d00532a318531fe36e75aed94a767dcfb9e17de5a72123242e3108ca99ea4010dd5eb176874e1aa3efc8fa5e3d3450f6c3ae5a55ecd15d68fad26e82ca28ddab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfdca7acb08c72adcc824f7325f4c75b1cac396cf29557805df4316ef91626119b2e94133ae285db2fb16120cdad72ccd8ce40a66a317d5edc9f65e0533a3db41385a46086337f3ed89e8b69c956dc569bda1877fc79750ac464528e3f8aa4b62d5b7354e69623cd1364d792edea89196;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73535c332e9a5776356509e4497ee0ccc73cae889a50c0a65e5f55f618554ee88a43f435214967d23192af50f3e7609b1491719c5f3351456a2137f6a05b4abb914332d9a5893ef9745dfcdf56392058b9af4161164f3e353b839ada96ab969dbc1280efdc88d443dd84bb9737d2933ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce41b8a6d9045e7d57c8123ab461e8e2666bc32ac452e837357691f09a8b07817f8c0abcdab6ab503310b9a476439804f3f9eadaeac3b750b6401f595c67343285225cd42ab3920022c89d0693e5f2f79e040fadd1a3370dd891f2252028435c8d35688f11a28c8f13950ff0b9da6a507;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d5d8177d895c6d148c6aa3e75c33f5428f63e597a6d6fe6b99e5ab73e334cf868f05f6aa5548240dfafd09a4156e19d5fda789b11c34571f1ee1fa20ed9b11c2fe340327b19e699b09f07458e26ba0528823017a8f04acf3afa8413c3b4cd52f4fa0bfd63ef7604323c05ef4aaeb1c99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd309e7a05ce7e96887ce48604fb774123ada63af0ebf3777d76a71e11f3293ad8f8ff452a8fecb413350bd19a3113374ce0e6050ae0f3b632cde5c9af6e3378b637a262733c4e8876db8ef2206f7ee6328ea53185fd4938e2a37549c6b59dafa8f9367bd336db089e56507279f903cfb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee27434fbe4d1232ce27ee114885b203c423fa63e37a3f5872c2b33f83d9f780c49c92af1f94f4691f70a6e088d555fd8548a60b54e9a17dcd99ad21b69d34f5b0f93e22e5ca14dc939e77ea77ebe7303b7d1fef9f56b513d4281fc439e6229d7ea9880546473e975c79393abd51b276e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c351446fef677ebf5b0c7c116278cd1c855ffe580b36a04dbc0877e96a1e09219b5790ed3adc3515f73e7af6e21ad57d1364fce8675ddb3ad1f378b208ee1198052a3361764522537e7956baf243a51346461c08c635cce796e43cc5ac7e62af4d18f4075c48bba230f32fca6b43ddc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd22f9c7c469e6ae0f3d629fd941c48d010c1db6b7019406e703278572fe50a332381e8883bebeb413b05ecebceff3f8011e4b8767280137271ab57fa2d778470a4414b951f64ca2411b4a5d54e15a1b061cc5bb6aaf6d09f0d398ef99a7554055f4ff14bd4eb788705dcf9576f6310544;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8e39f09dd15e87e85036adbd6219556d064acce29df24e2503838eb94b262c7ba58bb1c8a4e4371b8e96b54f1c19480fa4d50549119943dfe8381fae4a71857e68363e458bbb8b4f5cb86e6ba483f2ed02280a6f0b2b326f62b5d3e09efb219f7ba2bcdc6de4cec049f0686f33cc6eb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed0342bb456341e1ad503182b1dcd0e102e1967c3cf6660f50e3cad38a9da55c4ea3a7f943960a328f77707014ae349ff3068029967683041d371b568d698c508604f6818d66d7e8439e2cd447a5ba1770d83f5a30bb4a3145a304fb07eecd4dc26ca90dd62cbba98f5750d9d641e07ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf3b6e9bbc46c6babb23c6c5d9512a7e058c0c5535de1df25015d6112e407e72a3de758ba3c11d281dfbf490b711eee6646557d6f3b8df6f4257ed67c484d370cac9fd370fd3b04962f2ae76fa365576d9c15d6195e9de2f7b14aeb09669f4807ba57d7446a7255a3d0be3dbb927d8178;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb822aa7fd07075ff35271e36786bc83dcbf03edb34f1bbd13fd0c22e8e0d476f400aca2ac27c7b191177c99a9d0aeda9711853c77fa80a76e658ff493717482fde1b47fa3ab6c562938fc364ca1492384a4878a5eefe60b927787909a3172ac0fcc3da514609fc6eaa3ab102ecd729b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ab2bfc204db50d15d31d32d268eb8e7566926c28a91a914738eafb0686f2b1c6d16b76a9944e036e85c8ae715694cc2d8d17618bda9d74a1a5f7cbe93c7bfb895013af7e6b42e46e5831e3d6c4c41c690bb4339d26c47437fb3393b5476cb9fe3a6d68bd223d4f278d24d752ad475277;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf40ac8670328da00eee6276505c4f5b090d8ee64d4180d0915678ed8499bd0d5a63bf4a0ea9e8645af8feac91e46b6fb8f54e3984aa90703f1639bcb86c32aa95a98cfc9c347b6251888cf1e9d21741bb93ec08edddfc1796b088ff1b89faa27a7aafb640aa10b263e6754eecee050a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfcd3bf2603c512d3f6a6dd5156be56d5deb7587e16ec986dfc9b355f0d0365c8ab1846ce2f14a5b69ccbb34b84e66a879642c9c4958452491c59c9f1f97c43d091cbe80262c3b67ed2657ca7b5754faf840c31c3d7239dee058d2967400d33c45fcec397a5984a9482b32ff1909c474a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc553d97807d83bed667d7712c669a5cee434a7523a2c120c654fd16509dd047774c1e949e95feb4c95ec277f4607d7ad4f289b43569c8b21a4ba3f7ad5c71cad9a8c306f93f4e1e42a7d8a9b9fc94e4fb494eda28dc3630a5398184617861fe15293a259d40ba58fbf4c181577d3e148a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8cabdae4da400a6890b7b746a0d33b7e44c95259505d51a7330e9b58a4c404c8534e9100b00f2947d67629bb3814c3c605e42455ac4e332237399a48f930050d2bbd6f7530705ac6a3aa8b95389fcddf0760470707d33fe38609f328531b83f378b7eed4dfce7f98a3a0627d0b33fee8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3f877b39191c336fce86c5eb9680dadcd4be3d117864c5d77eaa093416f047a3fe0af01e502e6eea81c136a7dc50575e8b0dbae84f4c939e6cbec921948d5f3447c73269a9fa777a946d220af0eef839ade6d6e8abc77d83c3a304866d89655573e16f75c75673c8ad2cb4b25037894d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd89f18e5248f2861b328fdac5927cc41fccdd233f087a72f33707c370b23754af9516ab3300f78c143181f93aa802aef9a56aa8a61f1e1c84cfa6f614b7dda704dffe6f7e49bfd936206d3912b7363d29808daebd4c7bf956e7e4e933636bdda89509ec0203f33b0473fe2bc25d5fc27c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd238edd9b2d9399ad847d73dc1443a9655dc05f80b12876c10f88293ca76e9510469e45890b493fbc20c1abc75f8f1d401bce0c6ba8c0a0379d7c3643b54910b11c00af08b8df77eec26fb1298eeccfbe92e2d9c512dc2daf3470960b0364e40e7cfa688b9b1a97912fdf427180fb7e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba684c28dcdd8e992881f43c60a07b3b4a2d10cd22787294a0b72cc02a2b546dc885dc3d09f012fb4a1dfdbfcbe72275dcd7b0ce1a8dc12100ca9d4ce36157b4145711d2ea7b75b381462608ee2fc930abf4977ccb406fe3d9ed57b297eeecc0a0f7913a828347c33ca21426b4395bc4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed8fe36246df8a5c62ed5f035cb68a4479b12d8336af317e4469a4c5613b95322a8c8299b4f62f325441fb34383e5fe7906ffa1831f6e507a7639aad9cda0029983b558f81d57f73dfdf53cacc319c882fb38f04650b4ef779f7948752887444c4aa0b27ea69268849ba1914dd9b93969;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3deb847ac89b3d5b64d93b7c756136098c2518e6bd597a55e5ce47ef07c6fc6f10b21e1ef85e930de319a03708b1ad7c9962470f0b76a68ea34b5b27d10adab6d1ac7dadb65696f5ce237c8a6c298dd1774d00412dae3635918a57dd5b7926030169ca042fb2a4c2db960d7ed08cff9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h386b80122ce276dfdf976828f45c6a86dbeb2b7579863e3aaeffb32d5eaacbe472b7b5a530eb419509fe5bacd1469189db1497f56946e21d9925d057f47b2320d65dcc06b25396695747bb934cebc87fb158ab25635cfd072aba60c29bb146d9214a3733da7b20f67c9270d7da86fabb7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57c62fd8bff380146295758a123515eb1ba089e923c18d307ce1e4ea171ca9afed872ad425d1eff5d50e38a6cd3ea7e08dfe9b3a4b915fc399d830ed31f067458625cf869e02de45d77b615a156deabcc0239c0ac3101943135a929c6453d1e2495cba6b0a9a7dca88315903169653b15;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd983ddd25402d04b6244ef17f00a8995529e2301210cc83f2e7b919160547d044e217a42a1d1bcd65c2de2779a8b059ffc1e08019752f4a4ef4dd8c77e17681a9da05162606c0c742c953a63ba77bf68e0da6ad958258cd8aa97a3d004ce4b739f480f46ef924b9a6f06d6e4eca673e8d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff643aad4187c1df6912ef43929446e0f104aacfe3581fe23dc0660512e23d4d453fd408a13c0f1d0f86b88d198070cbc3731510736fe6d931043b60df3c5deba904f780a0c33a586bd576a4f7b93ff606dab838cb5aa98641609315ae563bf83b500ed0ce8909446390d4069d64b0a24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1bf2d920bd1803865c8ca38218e516d3b64161527977973942ed01ca4d58f14a5927fe37edbf1617801c8ff63dae42abc0b11fefb0f67508232f3491cea836ace68a44642487d2aa02a3573ede5aab4cf891de03f085b15936895ceb0a443cc66ad41f3a92dc681ad683fcef299aef06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa3417f4d2b04d5910d12baf1f1fd75a2645d5cadadaf455e8bcfa0b5337c840d4a25787b10c9a218a355f65a8f42fe9c14f9e58130e45cb043c4f63b6689368152643d2c1cc3c3300a5059597d15716752aaeb8368f66d25ae1391508301e071749736c3c0c8f9291a7b1eac5d15f631;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f17420f859ba8b2395e943b15da16ea482e986172c89b33f276d20688a1c9c9a70954efb0970f04b3dfa771c5b259724956a50fc657e70263b73a89ccf0b5ff3f3234ad1fbedfd538021348790875e860be2b6b510441d4666cac6e4c89fdfad90e95318f3cc619e41d28e19663f2299;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc58f8bdf37e4fdff2debbf1ae09d0ac6445a5e873a028ffae18cb0b6a69a76865db15d48ac548ecc947c8621efbdebb7a55a284275c302bcedd3c65cc6113f5022a1afe7dd55721b734209accea6c766cff70e02468710a0b4752da9e2acf5c164fc8fbc2dcc225903177cf90ed42c055;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19b018dc79d26a42b001f33123d4eb9a8250406b6284ae2f2fba13771c642c348a682c93e516d84e9e5a31f0e8269077620a64c7223345896fa16586c7f62b06a514c7e35f16ef25137ed3863db7b507595150ccdc81796d6947483bde0d9fe8b4148ae1e7c978ae08755bb09c2f4d1ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf90fbcfb20f45cda8d5a5266b5e58cad72246c7bc1c24c401baf58cf09e66df34389903f516e7fb73e44a71a0e0c8dadf24a63b704153bf5d748d654e81517cfb1f50202c869d1c887950ec6acbba235c44fcafa279c03a91e587f5660bfa8aacd834f4dd6a446efef92b3d14058fd662;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7d55a29eaa6f322fb4a22d82df46869f3916bc49dba26d9ab3082afaa1e447c2be98a917e0dffaad4f0463252230d50688887474c1f1d1a5e87632955b017bcd15efda41d789f5cce259661c9f96613613bf270e36c8f44fdc8efe8734663cedd5f73d6e0e36a9cc966d0e772d6dcb80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f005d56fc938d45afb8201bda96ba597dc8d8489a4fb395bed03915f33a0f9665c37327b04687f49dc8c00e91a1811e99a94c8c3e8a95b6f9ef166da59bac5429c789dd71aa4039cc5919fd44e1c1d0caa35898bc95164f56e236d2c20fe87d4a38ac1d10ea6067ba0f5f49a0b5ccb7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4188b072d4d9d1b3040d356925860558919ed1cb846525ba8598ae9e6fe467192595b2330ae6f2ec47de6f5967fc3f7015e062c786f7eb935c554a9a1ab46f20e1754a05b1cd1c91cb5c906a4c37cddba95dd9cd42d3057a2457a8f893168627043c807d527723f96324f14d3b09c38e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cd6377b23de56d367744ee08c165442c637e92288bebe8918df7f8719745b2230051edf1b8af6aa6b687e388f367137f6e908a9d895a91ddf211b6e5fe404ce577e311f4e73fcf45c4926f83b4cf9b034909d4b77bc93ce0edeaa3f5982c5dcca4293664820d709954d20e73ce31d75d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h542ce4e61e6fa7379799fd0800a6c8e987d9d382af70fb317c0124c17a6af9ccc894436dc8cfb7b405cf3925105834cb3d94c81978890e0df7391be6f0470da3126d0ce576825c06a0b91c8e3f115cd5ab95538759fae6a222e669263d5255379fc79b51e349ba3a1df49128fbb2fd753;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf83a1bffc6d0285f218174f02c83084022b71e3b63a297ed323feada1feed7cdf12f2591b3815d29cf0fb46dc4483088dc40cb91490541af5339999ff5c86ac7ef66a2aadfa385e866f62c298e41de4bb5c02b2ed4bd98ddb0e39bb8cf904167b70bdb0f903716fe4a669e4371d4c6ac3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf45c4f432caa34812a1e830209b5bf3524fcee289e5ae8b9a2d21d433929d208616d543d4a1b543ad87ef696da160f898f254ae659fb992a973bd0de54fc27758d6faa4a9a0e0fabba60faaf537fefb4f80cff03e92372a3560de516b13db05b1955a9e57a69c72f07d72c158fa7b682;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b2fec665f6f5fc6241f851b6e90483df5d7da72d0adccac835b76bb488700a2a4a88814f23373dae66b8b829dad55136f14d4c235e587a82f7ddf3ffb330407335e34bf79e85fe9b4d5b780cc245f88a76b907b2f7da1524a9970679cee281cff3b7f5ea4addc8d96fcb667fab86c616;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d79f96664f76cf304b905104dc747c74f2c69ec3222a77dbc6c4954bd7216bdace3672dd9b37db616331aabf6726e39549f8e063e7c41d9f59cd3428a44c6106debe4f1062243f575780f90c111d6fadfdca00c6825f674cd300bce3a7a9065c0cf8f79365b9b99c3446339ce610bb49;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f927e17dcfdab9b2c5cd4246639fc02e9f4817eb6d4a50b3c075da72c2e8997c2e180c2b88f7989aa4ed31a7c16937ee28f20bba5cb38979c00ea868b88d5ae97b653ee45e285726fd0722e107497bb06bc4b182fc0ea3d7e8a35e6cd87362ad3e9d10150c1448b64926b054e20d0bb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h429a70d0220a978967bd4fd713c1e0aeef5f2a3fddc0c1108830dd7f17df9638650df976c86c2d07c777abe27223e343e29d1b7a0b2c88f8d315ffa34652cdf71a9102a1de53cec034be798c0d34024d05eff50d2a03cf3a225e0cfc87b4c66a48cbbbf7994104e740bb9d4d7b75dcad4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfca107229b5e2b7f00cadea2913b212e32513cbbc5e3ec91cbf7072c39b88802d46310d14d816420f475354b0c50cc202e5259871ef851f2f69ab677d842f68a525c779bcd694882fcfabff9f65b11ae016d5863eed1c2bba45b4d5315b905c64c995b5ad9937b37074716ef13a4b660;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h461a390f9139d91d5121b3ca4bb9654f30e62c051ff23ca15dfda41c95e968025c7317a8bf2a9c652f006a24f2eec25c8b7ec2537fea9448e8ec0503cbb580174f5c22ee0827bad723d85be1be1ffae711ba8ce256b63534b3701afe74413354622ee056daa85e486808806b5f7862f56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h327ccf946d2eadfc6831ffabfb99bbda65340c8370c3a5d617c7bb5f6a5bad35a3adfa0a618a9cd024599e1465e71b01d8e703b645a271cff45aa5a64a4e22e67597aa0350a7ddc375beff37722f597f4b816e0287dbe012ede87dfc7d680f3841a72241f02be4a64e873587a117de21a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f277bc447f1a67288b4a26a1e1988d6304a5cc41b5deb3414fc0160067e786dfea3ab6289dcdeb958d1803a8bce836e0890838b7b26700f5d89acaf1cc057f950f8b221de8b4b91e4be6a6f098df78c3c7401ac287bf3a2e876fb24ef1357c8f839717eded5f53bafb0e65d961b9d77c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaa38ba4c4b63884283d9a37126cb89e7a4d64df90fb21040e308d0a64e3ba7c4e205be6a3000f2b5ecc32c614575eaa96dcf06571d379073907f58bde9f6ccd2af83e105965b7ef118b923058f4aee4a0ace97d7f726d8c804a8e66044a8d229bccb32eceaa93aafb7e43ddb2ddc516;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c666edcab6013238572fdd249ff6e0bb33320b9dc2d140b8e86b61eb1a387bf35341f48481d7af42acf533d4f4e60b22e7015842a27a959be19f3d8b8d24b1ead2eb7b695b7bbc287947cf670dead0106bcad2d43714c24fa99fe6c68bc90d8728bd8511cd8ca40f470ec3d6cab0a77c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8110c4ec5b0f7da830f607fb7152d267ccfe8837b0852e8b968ef7ca401b0d6d7c80c7c2032d66bb1e492cf65642f700b39b6f0294cea801dadd14a153ddd18283b5dd5396084541c846ec8b36dbbe4de4df2e29b384842b7b3d5e7f8ed20f669413eddee53d7621a805fc26d26daf3bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1de4fb2990b90abcaef42e1668e266247aeaddb2e2e67df0299f35222ba19f8e4d548261e690d4eea71a956de94f946118277498a80194cb2da93565f2b1cba3972567ce362f8388f5c0a6354566051403a1caef06ad16e22a3670d165bd643e5822526fad9c732074964a3cb0f84961;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1eecb82e63566241aa1f07758f6701b899884d778aff29970f9285246a183bb0cf96476f5e672a34ba8fb99ab302045520260d14119381cccc267700e88c44caef7440f9c67524a73cb194ef8d8d9b71e58b62d7091b8f471cf679db7851fe8d4cf1fb3e443d6134f81335ade4f9a51db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc24882b2afb068012cdb6f365306fee9be54b36378ee04e1f8ab2ce9737a0283580149d31684dd78ec491467ddfb82bb2bc94a0b706bd4b3fe30a5a5d6ac9ac96bc851e0e4933eed61faaf260ad931ff3f6e623c6cdc71e77eb44416ee2ddb0e801182b00277655efcd205e7a2a485290;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha61e622dec16ccc2c2909b89ea99d080f71c8c4dd250899fd67edbbb26cb2c93155d12e7f1395830e1101ca0a76e9015d583415b47afbf885b620fd05b05b83eeeca05512b12bebecf56b8487fb8e98785405d58e5c27c9d38c1d18a02ab6a5acbb52c9e2b4af07e479d34837d53f28b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c803c3e61afc4e5c4bfa1d54e14d88326fd2fcef9faee829888285e309e33fc9bee56002eced52620f680a40e37815f3a5bbe642e5d878e29f3d28ebf831eb96acf90f494fe87033abe546b7d30d87cab1ae3bc26434dfa1c87395008dea9dcc742b2584cfa81350fe4d02c07d165489;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd740e88c242091e288ae94dfa68e44867f18d716c8094de42ed88432820125fc9acdd54e157e9a10b04b168249e34e6b7154d2a7b86591f7ab3e863be589705e3fbe25f1ce0cecd9f07fa77d5329c3b83501a6c6eb37426add6a7c35df457672a5e28ee7f2442c25d6c178dd3bcf66466;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h337566baafc8f25190bbc8e21a45b0932890c3762f7dcab2fe0e14f9320c165e8cbe74ba89adefd7809475f79def44bf5d39fc75632a5dc569a92d30408d012171400da9970a6e67e5aa0254115ba8cbd5a21d581d3b57737b14d80deeaeeef22935b7b519fa0b1b9ec065475fb0847a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5017d38bb7bfdb895cd5d229c6b2edc9c650f105e933fce60687527591d10851af050e6c62ce778b26055dc2474058f7b39f57058ed9728ff32f88f3989c7a68aaff2a8310bc9b743e099f1f0a5591f11df43f5932f94d4888621358caef012598d18b59f9bb63e09d4b3163be0440f6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21a8072df73fd6dd50cb911981634981873c9c622d75857e8b64b910b02ed2003631bf928ee60d253213c3c540f0fd3fe31a7092ce17a0a60d79397396460a31507c8e9c14452fef220415dc32bd1c5da627554614df7584655edfb5d5a69c31d57681434cc85a26fd273179f5466ca86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2659815bb19c99464c5c109200d7a45f0a5c6e78d6978e74d3ebb87e2603c7805c25a6458b8515b65cf5926f3024af05bcbb684ff70e83eb750bad75f2a3395cb09639bbac366f9d5be7ca63122319340ae5c00457038597575cd6d87485b5754ea605068eae3773a787e6939ac38b99d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90cf5966c7227d9bf64eb311b824de239e50e535b35103b2d84f6fe058dc1bcd369f6b13c328c68afc9700f69148794e33fd9c7118fcfe5dd8a87556a0f6d4333038ceb647a850ab7eb94b43de8a97aebb358465a800617af0af72c9d8f6de55fbf5f8c42eeeaa3cba0b9ee89e11b9eb6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f2fd79421a1c5d3d4d8321306c7136aa15239253ea382d15c0842ec890f01004491c4f0b6a9900405c4dec742497a221b1873a89efbf131db329462ad30c753b0f4c503d168070e2ccb2466fc11ba9eb6326029930ec7a86c8b6c3181ac83741cc80162cdb6e442917f51c8fe2cb53b2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81f3176e0d7909625fbc835972da961afa447aa1cbb2809a09d99651e9f38af672462029a04610cdb4d3ab376814838045ebca34d17f84648cd748e7be945e765928ae1eaa6c74e53ae00aae6f7c0b18ac8d22dd71779caaac16e073185ee84786cf8fec4f9b9201a6dc6849efbcbded3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h377a05ac66e34270f8904837600fef72a0c497349c43d82aeb86f73864148f7cc1255e2cb4396836308079d6edd43b5392af0c6fb37d628bc5bdf9459e5f684cc5bf177e9404473c6005f0463556a6e22b800ec4bdbd83c8a7d3a601e714f919fd527a2cce61a3cb99126ca16135e0314;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h792a1057b544003fffcecb126ef5a2d529ce633f8afb92c0bba044e8a784824d653a9cd15e8d5448bbdff7227eae4614fc298ee2b4c3897f4f788abd3d931675290d43a106f8b4f08f16b11d775b386218854565a53c580c5ef4fe435c5631685f74d7c102721c4bc145e60ce67e8e534;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d39c92b8667581553719a499d905247255233e3e57f6078db447972c2e5ee22a6a83364cecca9be965fbe5b773a753eea2d1876d20f35306bc3a7f104109fa213345393547ec67172808f3b0828861f96b07242a96fb2c8dbe7d1d731c00b490c0220a2b0ef503486fa8a33064aacb56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h109fedc8f8b50384f41f4bb7269d50794468c950decbe7fbccd6f2725be73c61e5caa84518570b0d90a2686a81884b3fa7f0a8f5c989edef6e8410f2524a9dbbc198a3cd3cbe8586456dcb3743c524e7a849ba20e2b8bf1a5403c4685db13753b9dcb650f7e21a62c0b20a5c8d933021f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h967c0f8d74f373bd85e76b030ddb02379cfbad87ded7e18e1d79067583e741dc0ffe0460e673ccf540fb4d0745d8494b6ca7991952f488474547f62acc5f325fb1a5fa42241c704a9f678de389647e1da946b8679d993536f03a833ef0879d06d2d0f71b160b5fe456b07ca22ab9d7cd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e0a59f3e9e8c27be76d99c556c0f648298d0c28032b6992eb571994875e89656f855d6b77ef9b3b508f1b92d153d522a9e88146c7ce5ca5e98cb6ce6c6039d7641387eb7c2b3eb9233618089fea32244d30c66c8d8e100badca48d2c34a777a240df34e549f6fdf704024e5cdfa98fbd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40588ee0bfc4d34122b4f77e6b7ddbc5a04b320fc360db6e3a9f58e35b19007fe4f8d292c8aa7fcb701339120a6a8a1dde728ed7e2143518e7b04b9c07610b24c7c63015a0990acf21b55838e57d193688598f68b595f1000e829b8a841a494a29483b45fea440ef4cecd02fef59fe32c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h210480a5bf643df32e00f8c6dad93de748ab9a10176fbc83b35ef3042a52f4ea8834fb9dce34b004de3d88e1a234a07c1c1a47d4f6910f5826a493eb21de98b88a4a678d21680a715f216e41def2a8a1a7bdadd4b317cf619c60913c1b3f959ecd09459329a01d633e29de429541364f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84561a31b5a574e9e78fbafe52b9d7952700ee909e464bf4e57a4e55ffd3eb58a503082a36e9e9d6668c73676405f06990d50ce460911066af7d8adef336b22576c27b5f9b6d9562e0ff83e570bb971857e376a070c722267f837759ae1f24689615184172fd9590abc1b1d8392f231f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467b69ac1e34b4320f1b4fb46369122eb601b959919a4576eb227c593581316b746419a951f052e10e5cb5b0f03c4f77c2e71f352636e5b1c6db9a946dbc8230c399a9473bd9f0444f81cbb76658ce1e7e4b6e2aa353eaf952f892fbfcabccaee6c6319ab01de40c633b1d48aaf9f476b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfbbcc6bf012b8ff59d63b3cfbeb940641344b2dcc27c55a174d7c61e465532f71f144d1fe7796c991d8367a7775e6a05bb3f33890b92e2740f4fbd1d4725f2830dfa5bd92c3b3a7a333b93be3ce7eefe2a877953cdf83d5eef3c97394fb02fea970d532c14e758e88cfcd6eeb943ca92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9c618eba74cb7b0d39cd1158e6b1ebda69edb61b5170ad9fc0626fff84eeec6c363e8432c1cd124258fcecf6063a11e536476de745a06564d8ee31a88acb4bd9788e3398ac66da9c1d66bcdcabccc38f89cc42aab606457d7b5f2e5c797316c6ed26aac5f8cd5519b075240c47fc6d93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc247d5b5dc17b33a169ea1aed88075f0a7fb4f07a990da20f7ea98f2d1d5f2535849d834b4064dc0b9e1396b1b8416f57bc4bbbf25b76ecddd53acfdd5da0c2c242db1efd9d7198af000d49ca7c3706c75b9c09150ff58258bc2aee8a1071fa9c69621620037ac038da5c934859792429;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2c3e7e2fdf4ae59a8b3f321839e6e49829829d2273c64805fbc08b6304840ff501736330b7be9c01b3c3f708beab55e03e0f7e57f2027ddf3d37f06f218fab5a74b311ff6d962851f8c16f7f7cc212c5adac4e0e5da9d352a50b4ed90e5d4c4c1f3e498070b5776a6a5b72b3b808ff6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c86f468f73ac5c8fffe6d8b6bb328ae489a76a454d2ad437a40a67ba296058467668251c3628188a677fe3ba3395e25fa722dc3c578870f82ed9c9b89cf2eb4e9a8caa5a55faa406ac36e31255bf820147706e53139269815942eb0df3edaeb1792994965a786b8dca8acbfd40dde60d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95262d0668d2293962e120d4efff19c82b556de5b33d4333fa120585df5ece80381624c2d1b98989e67e56d96e217bf6c981f95515f6106732376b1d141e2523a4a55d347cb32811f2efa4a3360cb7e6865d8bef275536b0456962e8b24f80acf5c49f6304b4af03eaa7cdc5f3cbae259;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e8c38d974926df9388d225ffcac399ef408860152bd6e3002b62a500bfe633dc76983ed6e016bc7c1adccb35a34c7aa18bce5424e9113cf777405e6ce6bf9d41ea808a8c2ae9a0fb3886c4f3b0035da7ecd802ce722f81a02bbbc2b18c27d80fa9758c0c1be68fa7787a950cb4fc3a86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49954a2c5d430fbcca405bdbad39feaa928c4c81adefe1f392e3d3f4cbff90dc5fbbe4cefe1667cb8f8b3b23e30a21bbc6164bde31dd6faf6d25d423bd87f519e6d5879a9e9f89dbe36eb7010bb1cd8cb21b7436f06c6c681b2a19f3f10d2e821dedfccadf8236cdc723ad9b9fbd9117f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4635fe3756dfcc21bb1a84de4de7dc06e5d609a09e8255c7dc4423733410cddf5364eabd2c1ce0b0c1adf817acb8b9a891b12003ee1b70422b71ca6947d72aa9505cb52355eab5eec3dee0cd4663398d0fbc56f66065e32b8947da267bec77bb2000fa137e21c35584fd779329c3ebcc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b1f0405c2b42da0ab4420ec132845ce6e3e94b7c6361c3b1adb1c6295218a3f5c449308bff84afe6522e47b26721c733843c8d285c299ba7c399c65f7af6fd8b9a99795618073c2a83dabfef9a4500df80b8900348f64fd316dd88a15e364ba06475e1fea4b67b2ec61548cbc7067dd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b016431925b7fd9a4a381118862fcf10bbddcbc479852b3735d2b211ccaa6240c90ea80514c43e215f597ec6b5c96f0600f278295f162412a98e509f19c13ce21e98a26634478dbb36510ee538830f82aa296974e6c3722cdb867c4298f1f2fc4211c5b2e61ef81f013dab57f7ad0af8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5d813e97202f2d779d67365d7513ac0d9628a76b2ab0ff62eae8e0298663613000c43a40dbca9800e3bfc7fa0c4381789e9d1086f6d0ed98e486bd04d56f09b7c9d4355e59f9b17f8395e583bb30e6ad9591196f7977634e5043ed5e80982a0dae1d4a583be96f9babb16fbb52d975e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4859aa6730cdf0e1760b9bb541519ed146a18256360cd0079e77af93447bc3d2e974d1e6ff5e58435aa96537b9b7c31321de54bebcc28f072e3109a87835c7b789dfdedb4b4115f3fe73a5304f9cc9e8c7ffa60c202eb3a0ea4e29f8a2b56e447997e15f0b1d810250992b045ad39bef6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha768c081f525125d7cf1afb0329b74ca64581f9efac1fb15400461ac0f5206a24aaaca9f833b202a0d6b937e90d0802c84a4a31346a82a7802f5fe5ac89b2d257b326000fa6ce6930c4ec401e15aa49cfd8dcfff71e70de05e4188e3b8116002e611535f136278788c74bfbf51b5f2411;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h105877bea09d459018792e32b612571f1382d850c4472a4cb0469bdce4e98e340f4020dd0201174c6369666736cc6e8453af1bebfef60a18a178ba10e69020d655caede0785731c628c8b6a5c2d3b88274cf243fce91cd4d9c32bcf1b58c977587e6b3a1ec4e766d2a37c8c2edff31301;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5329bb5ecf8c5bd31fef1df0c31c53fa10a9a5456527148fa57258eb9573ae967e85762ec2c96d8f1442d5b2d583fc09d6a67537d76f80e26549e847fa0c3de6ad5064e075fe86d888d274a8a005102b73a6effbe4a3bbc121f357ea1fe81d45b479f5ac5e1aa6aafb64fbdd254058d11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb736e32f2a76ef160d3f412b5b86cb68a70bc51a792af7fb83cd2188a5dcd7c164d04235614e70f299273bc0a5ac4845482552b5da9761b57bff5cc471abbda0fa4960f46acf7c1a4584aa829bfe00459c5929e697f761ac6afc3335f2521e37affcef4fea6e42107021f17e81ee5b2ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5daa1a7b61f075fe1525124804038f78426b56ab12db4b868e8fe738fe1fa1a4e6d1e8f0ec521ac6148a8a455201946faa8515ed4bd6d5a93a881521eddf33cb165428a7d4376f795084443dc34c9099dc4a573554223e8a1f274b7af1451e28e3c6a7c6d81b3dd533bced7a67e0698a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6f47a7efcfbb88799625663091d409b087a57da1cf6f84cdd06b2b248eed85e8296a6fb7d15bda883b7e9bc55856f7e549feb6077cd42898b369d797afe0b305cdac84ad5f554b488bb7536b1fe698c5bb71f00a068eb658de7b9557b4af69a74d31e5f74ad13ea110e84d1ab5d2c968;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7025addfdebc986add01ca0190d3a6176b43a4038a16c9d0abd238e02821cd08a309102a533a0e674ff8b164140dbe23325de0f0613c3243b7fe722a162bd791afc3c2275d8df9d8b188f8f5ff6aa80fd9a649ccb04821f0417c84247b4e730a7328bbef8011b09f5c9fbdea6554e15d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h944f1fd7c77877b921c8d46be76232d3ca548e3dff41395691a4a38af0270384d0216beecb0f7a207586e0b0a47f69339cf28e4628c133f6e73794053bd597e0ee108b7a4ed58dd4105592351e1e54527a9ee7c257513728d19a2bbdd84e4125db88d4f47b15ba93c6045d17620c0e501;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h646545935194a5878c25212e1671e4e1b57cc740612e39ac9ef31c2870ae6bf0791d7f39d3b38848b6eeb55e8b0b033c49532a320c9526aa8788a152e72018e710c07f556127f888c1fc3b022c15742ddb716c10dec7b8eec7c93f110550a9078a27f44a7f40102b87a3cd5559ed88340;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58d1229c5abbf2f48dcc64afcae8b6d890f7ef79e2f732f14dcd9fe3fe0701eb6cd796942b657f75d17a637a1e146d8cfb80b2c4874750b65b85098e05e469ef9eecc15fd8a5b9a255f7a5dde6075ba60e36e7e082f86d5ae4bc4c63867549c624b4a335eb409691e6198a3e044b2957c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h319f6bfece1bb296155f798539b542b1566595bf2d4e578abe0b13ffeed498d8bf2ffedb7c256e5b9de39130bf3cf9bdab55414c307adcccaf11fadcc400d123089dea11e5562b9dedd5b34adb78d09325ffba37e2cc7182638db89888a2a912fc7b489953631fbe3f22b012334bde83f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he931ee46aeae07134f77c4283d272c46ac8fb7130054381adcf564dc665440a030abf4cfa52e3e349a59772caba5e36d6ae5d8837d6d5d1ab3304ff590e5439c88f00cfd0903af11c12a91197eb77a6767d8a160825cfe0b83f088efadd3941ecc630b8dc8e46502cb31d9581e342300f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a8fc96eec45946538e94669b89575709ba2d78ccb68e389397304d200b3546f5f41cef4ca6b56488743852f007a304359bafbc6b915fa9dd4fef5eafadd33c4a076d4afa324e56a7b48498350ff4cac0d26211da332cbe6d0de72c37b45e2af9400eab28ffc4aae33d37a03f0994e4ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3789fb7974ce14fb91f5579874b5535e9acecaa954b0111063ecf9aa47922f9958b9c0408238bc7d418f0ba092a71624e72941ff13022c1b02b909d3464e21acc49c2533daa7edea125b50d5fd9bb7f8d49ae5cab233f5a20e2f7b97de1843faa75962333af9333c5a0458f70237a97ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef6b0d02ac81c951cf005a591dcd6c907b182ba3ce711e33010a18f9619170e8a2761c0cde9d7ba22681b3ccb55ee95c0b19aef54e2b6379d3b1f6b6e60fe939e6d09eaa9e559aaa7314dbc0ec386642eef6c6f5f54dc77ff4963f3d4f0d27b4b9eba7812d724cd9f53c672dc3c41bb3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haba32b06be3bc83ab200ee3841ee13689bc0913e63694b5049d3122937b5e8eb5c9a9ab203c1244090ba463d3962f3cc3a218fdaad32c4556122bb7b59d4ab35f8e8d850b362deed2b5bf0af93e36aed436b755240415c3cb86b644213f24dcf45516b0c85e67d35ff770c649852d5a42;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2dc19a65620b439e9ad92b2761dbbce9170c7ed8d81e260251258b2ea64935a562ff3c2a43c0bcaf3e3742a9823b76340ed51e9e3f6e330ef8ee6f4987e94901a2cc167283f95d0945ad0fe1595c45a8df5b5966f123c7aa80eebc60c256659e0ab242286783bf971a9cb444a8af4f9f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51d3b2ccdecf3aa750f93750d60a95a7db395f061fd7c5c77c993faaa8d1ed44c7e18cea8b70466d5f03a31484e8c8836e3e15c242eba64f5e7629d52ffba65fb3ae93cd8d8efd0e12f11a66fab27d91f5c58f994a2e78ee32a68f68ca1044b07d02eb675ad90da25cd5d11da5cf44060;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dd40548333de249e56dc602e11f964f6054daba6c515088511e37c0625f9fa10a5695df18f3a247554a9210a61025fa65bc52cb17bfefd24df2d3afe1ae3205da133a2d0c622a177fbcacba273f4d8d99cce5ce3487fe623a01811bb1a44a6e8289535c7db7562c4cd94f9b5eb295900;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbf036c36ff5676dfa4cb8d95c640350003d4e5eb651eb75101c2073912361ac523857f9a3ca4b0d4b9b024e2fe1e67acc93a5ec13d4c9495f7f5fdca4c1272fb21b9f727d7523f5ab4caba738061470d9940c3f573d9690d3ff104468d47ceee7406d2521805494c88809815547a2ed1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77aa13a80bdbb341e2379bf06fb8dc2a8b2753b357a45710d3ed6f4834e4d3c2f2a3a72dd45f63f3c14cf73b3da7d7d5bb7dbbf07f0823394fa400201cf2fddd69686b5cdbfc27d21886782f8cbe4dced4dc14d9031d156058453f731f1429e02666a89a26a084bbabec30d1389ebcb59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7df3a03b531c4525bdced9664212c09b750f0352b4fc906264e714de2246596d3acf090da8e85648feacc92bd4eca40606320eae35589303ca39d7b4392c6a1bb140264a3f4801a0d14e1ef35a5187504e0941e06b1be6242d9e65dd36c132718e55a2b2d5f7eaa11dc54802905e61d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h227f92f6f97afdd9dbd5482f69e3e382f8cda2bb66d05f3949a05a01766515c3951439efef93ab6a4e314963e6de3ec98a22e4ffd3a9559c744d49266276598fa3cae1e04a8c35d04f1f7ec64d42d7964a9ffe361abdbd6648e725ad4f7db6e053e7762aee57232993ba873638a89f838;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e96daebf9abb2718355ce3add67f6d4af49bae77159b1ae95b2c06f91f37b171a6b5442027d9402115b7282fffa4783d2d2f3ea157e56a766e2e7c529216eadd6f3ffe0bfc270651d7b2318f486707df2841c127fe1c00a020ce7c4c5dc8bd2413419596e011c0f70d180c97d214b60a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb54eae80277f2568cdeed098040211cfe3a0f3ec4bacb6050b16a04f5c912c1ffd777634de22ff70d66feb764161ddb8320e1614e055bdb2c5b306c0d9829e97f9829e61c3153b1091e87e46630229ccc2f85532f0588b1dfa5c93ec030d9b4ddfea6f36d39b6669ba30c12781843ecd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99348f75204712c305f6565ebd11b9a62ff8858c1dd39a859c6a6499875079c1c788953a6f0a37eaa7b4b9f529707310a43b5df08373b88f587f1486f3a7d8701c156787d75940c576bd32f11bcb17b5baefa3b51a3dfd5099d0a2695c1e9359e2b508d26ac87e6032d03921d70a04bd6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50de82d2faeb6a2dacd04b40486a0d54341107dd1eb66a8e77d46e4eb15cdbbb520636f9d890bebe6d1133ea448dddae8f315b13779189bcd42ee0f354642c3051a99f9f64a04e5c9c377f00efe9b48dfc42d52e53209c973da0b7eb0d9fdfa1b852f22a4da17d61b744bdb7a75784846;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58f96605785be0cd09c4fa44a786f1d665186c57f5a5be154f4800f1106e1ec640391d8253c4f680afe69f44b0f372161a02238834fcce3f7c22b11baf14f52d94addedf5164ef6c758b5c33cc309ad737c267dff3f3a078134fcf82c48077ab0a64ba4ba2bca8d495e048fce0f26f830;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf078cf36e276c3028250c9a30b79e867ba27b19f99bf9fa6900d21f5a78fda42283608a001512a2fb817c3da911c1c4063b52be3b6f423e1d9fb5236e950ed4702559222def1f5a2384d05d4ada48e514f69983cd27fd22f03e72efc23229a4ff400d823e80c449266f45c86c8a715d18;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ae843a0d5f9a53d50b22ff13076ef3896d7d42e2bd7d2a15cc57f0e2a96a6b1c9402b73000fcdc0399d4aa0bf3a7923ebe78de99325f0d34fb65b44390c9053fc0fdb4f34434b13c738984571ee90d0f995712c7d256ec2660270b8b33a5b66beac0b01c2fdd066b3ac3b66663cb323c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f0b9ad136cbfe07c697cdcd9e92605864566aea78320ec94d7ea2bc41c0125ebeb72dc6b269dc613aab0f30ee28b666c242f550554826bc7f19850f24931fff1c7a87e6b2ef566b8d30f0e219f9294310b0e19aef226336d3e2a92f3c137fe502157b58f4bb8be6faef88bde12ce21dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c5052f598c8a4c571b24e5a0c2f1d814e4d93814ae1171e5f51f7c4f8af4bf65b386725e62ca34c0cbbbb80612d6e458d6905a35033b63d3c6898919dcd129c4670df244f7dcb7a903bbc8bc451c14511f33653b7efd29735ca6896c69a6d7982bed75766be55cc6fc3c480924e9bed7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25d1bb0126606d0c7ed5c5cf48a127ed3536ccc4351e1af821bea4bc605b7a1f677c8e0956584c3c0df292ad2e215d7575776288b902ca344054fcd1a6dd3310def5a3ef8bb74822c8e293852c47095d3935c5d9c47689b33fffa6047b23751b73629fc6d626cafffe5c47540a223df53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ca28fd0723d4350e4c8f332c9946f5c927415dcefacd235d40465a7f388e990c6b57ca6cec2614a56193a37ccf9f3d21f69201c8cab598fbe3fca577643b46b93476f999cfba9d10d2e776a4a0f5ddb79b0ce3930599199f91997b5d543550ed3a07a1f228c22aaf6584b19e18b8884b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80cb7dbc72e97cc6c43bf54feb4033705c3d34bd2491463904372b4f804ba71226df92c3b0cfa2efa1ec56636f505586d890298f36361e969cbadb8dd2a4b251ae05f3da7f53aadc8f8365af4936a39bd888868a9aa29084e7d138334279615cbd5ba06a1195b7c33952169b2fa30d573;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd70d7bcec58f736f9090c7d77ca44c983af214d79fe7ee2a75f3437087b9f8050190aa80a478cbacf84bbe4f71d1f4daff18c85314c687866d923496c555c866607728563eb9b839f91d42e9b442463e910c09e0a0c0f0547771fb783732db9da2c34a7e5ba2f4d157ed926c4b890c079;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h198d5978e2bb0b8d3d51642dd2484c641726b1f394d7c8985a14a44e4ea6fcf7be072acd55ee6aec16ef67daa4bb83856ae81d1384eb729c303a2861bcf116888ccbd26ef40092a4f794eeaef232c930114f0ea32800e4eab87238f282206d022666bdae99a3ddaf9fc0886a9d6fd2d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aeddf366cfbe9f8fa425d66ba74ebcc3c85e72f76d65c3e09569ca8b0e60394f9d4db4373896f9056f0086c1c4ad682256dfe2ef81747cbb2279655275b73c592300d72b8993a225d3e4b8f6717f1184b55aca2c59ba680ce0fd2f1a0438d29691a72191bede00a05701b618baca4607;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf61e99f78c62d460557b4e7b60f471936a5fa68e4815c620ec4b3396321ee626276b9cd7cc93b56f8bccaca8a5b27d33059783dd6c1030f52073af0987f20580177cd66ca6b4dced86e9cedf9feab63357c2f7d5522cd7301708963b2bfa9a5929c8bac939696aed12110ad76106f1e81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac225f44a7b1c368af86cdd311f159a96229d1ada86fca84be1cd45d879081efec6d1be7eca414d8fb5eeda06151f1d961d3a8eb35e2cf864a1c0155aed0c83f2a973bf1268e2178787d8546594f4fcc969e7fb0fc1054a0b8affa412701dd532995f16646e7874c020b7260e4f1b0bbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5dd7a8d74c3f1e4684a0aa93fd7ed38980bb66eac0feffef47658227c9195a4b5b18c4d59eb6f8f3b0b4680bb2ba664b0a80276013279879ddabd3e779efc2e569ccd95901c04b50816f447b6e47f18938ec1d8f7b4f47e5c9fccb930330c9c0fd1d1e0831b5d7e0470c13572280ddb5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26166e44132b0fd5d31f06a96a809a6d39d8f9471c004c1a7057523ab6cd056bfac3ca91baa7d194aaa862e788336c25bcecae67a5aad172b996cda57e7458c9f99aee5ea9673de0d318ffc71e6d0b1a6706c294d3c488932f6fb0d720627a0b5f16dc461e0daa65d35a995c90a4cd219;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2851e0b5a51821605ef20323cb1d5ff8dba253e4c2d41e603779d7d6376cddfd7a7a3e34fa5e8289a5ad715d524d9a54d41c6dbaea0d2f2ab3e79b635330768afcc6e70bab2f63866a9dd8d3593e97fc1f0895635f5849764e60817e787ea97c6fef49b11f727def6bd85b42b3360e52d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4323520a51f6061f04bfe80dc4b0f08a64f9f905e4e0f8369df85ef8216e19a72a01a3cf1f467b6781a0d2defab07fe09e1972575ed4fc8c5d98bcd903b12b0a346c0a6040e06e93a7da578806e000ffb349862cb591c4c8e5deaac4f82e2af780f6ba15e609adc0d554ea7e91aa731;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ac4ba860f28f5674bbae57fa3b68ad0f3be72a5d33076fe30a670e6f0c0b4ca13d8166a9c1cd51634f6906f24f0a7e1c14e5bd192e04ba2a8d97f1e77213dfc075670eaa13f22f19809175dfdeca4726bbb59aa9af1714aa1b68693e7347670897d42297c81d280938dfcc2a5a14a761;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16b9d128938cf16b8b58eb6538ef78a5b87859e9abc0f3eef905ecab5f802916fc004497ab9a048a6fc11dc6ebc3bf0ba699daf6fc27c4f606316ca68c4bce6ffc4977cc1e311cff1dc97b5029577805f3178c5f07ef89a508206b3b3cbfe4a1d177e8c22a072ee321783d0b9d426b4cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h798a66bc3760f87608e222096f09e2980f2dd15a4dd5ab0801dbc96d1b7189336355d0bcffa801d726c3c23eea7982a9b6bdeca4320fe70d7273c6d7b4fa773d59f16210de223ac2dc3a446eab600cb035f9d3da81893cc4462fb54d3443bd6d3d816193ebe562b8c49d9f9e5f00a6df9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a529413a1f68a8135ec6b49b3dc12e8d2e1187524def9b5ca923d8e11292787b7e6dcb1212bac6b57675b8e9822c1134f03b6497007337cd9eed3f2dc2fe3ac5b8c6796321951dddaf16519081943be76902f8cfc407ba5a00da56b1c323a4798fde09e955adda26ce52cb4e7c0683a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cb0a73f594f7fb2dcecb4d9545e02deb02d80bf36d56d37809b0804489d8cc4fcddcd623367d27cc9e438ca0d5db71801226968e623715c0a8710a2b145d19dad2222aa46393457fa1e9d8c4b9bc74d73afd6d6b692d013844f9dc2057839ba328ff08e99c98a06a88e370a7a92d7d60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d7f76ac741c6d21a418a0edea42a1a08172c79c17cb3022a2eb35fbeb70061cb8e6a79d7ecd4eec33ac156bfc63c73287e8e29eac01243de2a1233949d2ce81f168ee32625ea2520d261374f8ea705eb3bfc33d7b970e11307fa8cedff73429ba9818f064c5be26ab3dbeb2aa585d81d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4925e1c2602fb12690d1719e30ae0bb37880f4567718b58de8610c6d8bab8d09b4705f535482e8a98114a244fc00f483a6ab862721c25fc5258bcda3199e1fcd9d8aeeb37ed82b006ce6fa665b9ca3398e6d1b043124e4914be276ebad085aa1992d962f42f02e4f3d317efefa22938ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ebdfd7b2f136dace390b12e517e6c2fbb36229b5f96e5f49a0812d48b238d8abb4e23a5a04bcd5d9e9ab1ed1e1099dc405b787fef97b82419760f266917e2970ebcccc62847f2b5af2ee6d23c8b9dd95fb29ec787ef225eb60c31a6967f8eeaf1904027b346548d1a3c6f061a3d3b695;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf1db0726b40438ffc70494f4ba3036f2ca265376af6285eef8859890dcf2c89bcd40d0edd810bac15ef33e946fe536243b24b3c1d590b5aafcafdafc5283be0ef8a959eb9057fe00e3e6f14a8dd67b520ada2151dd1a27d634c4d97c63c4790af9571711c5a60abfd7ceb7ddcd7f72bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7c5dee22d1134609aae93fb7be53b1dd1d68d7abd2cff0c3a1693a537449d534a01d754f7b07b636db41d9ca890b996fdf82c17beccc101fef96171f76bd8ba20496917ff7e4439d3b4c2fe2091d547f722b366735008eb7aa8564d623d9a4fedb88aca0e3f44be188e60527b440235d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6421fe077e1889be4a7ebb96d837c97f3aa6998e89d15c4663989a0713a51478d25cfc2aec25df186a23810aee9044a4de0ebc3eac0b34a90bd2218d17db8f9e4f8623a863d784781cf0e74b34183e6be552b35a36555e84b5ed35ea7c89ee02481072cdd18074469e9c0368649c1d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b873b9c3007d8cbab8cc69ab2641b7c8d958793ff5c93b7f4052e2943ea6e8ef1c6b1c7d6f0a252f9dddaf12989ac7561c3b44d5bc243b2270bbcfc4de8cf7e054e610d6669638abdb4bcafaa24544db8e6d71279055f3a6ad6d51fd2246922064bc530140f6a74a015a20174269930f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9dbfb0264b80052edf89b79c9d9cc56a38e5183a2239e2d1cdc08eef73b4ff20248e0300c841aafcebfbee52b9dca99e0a27a12e5a589392d210f89567cd2363f5ccc5750c6518c81ecc658e7d66b0245a048fabb3548aecba4f3725cdf955118be4a4f5dc7930c0fd08337e483e2de25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb9ac7e3a18bac82ce14af96195d8e829a03ab16ce28370719c99963faa68a7d63d515d1545a6c638aabfffc431328cb185486ffc1cb990aee1533936ca26035ceb94ba59268952daf4a05aa37511e92fc757ea54b5b99463809ba7776e1f8d4619cb3c834fe8587ba48229e4c8b4d38f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9acd6e072f0c750ea732d4993c4907e103350d1d52bbd96c263f38e9bc2e07cc95806807af8af000489bd0b46187b2d3a0693193bc441f0a9998200d22c8fda6b524cb9db72fa24cbd762381bce40f381617fd5c89e7d682d5bfea874ef2d0d9446bedd4beed27f4e926b8e5e9513db7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d3796675ee1bbcd8443af04c0f6e2c63f0fc80356401a95693a254276211e079253fa28fafd813906670906af85902b590aa2747b8b3d176b2f5dee0c7c7c8e61ee50b4afe2652f4852ff40195d9ca614cbc6520fb01b94a4e834727976d28d1faf35d04aeeb5aa427d15d6e5fcdcdec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d4ae24ce46bc58bc94d77fe07600e803a90afe02b7e95144722ceeced0062788952a5d488f2a4b0bbcbbd8c4377716aefb3534e5f5ea9df2113f16135c9b573fac0ab2cd4ce864b82ab8e0123d2cb12286af988998ea793c7eb05c367ea06d4a2f3e47572a2f82df3140e783ead7ecf3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbf88b1543ee7feb42def43af234312b64c8f03767e0e3c381eccaa27651a053e5b4b7dc6998035617b30543828508379f8fd29d9ddb6b31c1f267f0597c7e64a88269adbe5adeea6043dc36f451a5c31c1146c3b3c595d06ae5d6c156da7e7fc1505e72dde9e9c5c830a3523cf2c9461;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ef7a16b0a02eca55b3f5992daaf54923f2eb138107ebf44db93af06fe6f7c4c4c66b84d9ff3255c23a38363074d2c43c66306237999b6e894fb02db6a91b6a1866b18739e48ad0dc11733ff0731b83a48d9980eafba3ed036d84400fe005049c5e457aed5947bcca6fdc5fd3c6acaee1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39ea210a2fc5d8dd9a627aed800eb0a98c25e88ef0fe097cd8ceddb7e42afdad20fa3254135f80f48a9e49eb7498c50337294aabce6d693135d109228f2ca6b34e72ae29e315f28d0fc25ccbe7f6e76707e0674595e20ab0b75e2db82c026d556a866ad2bd996ea891d57360af66b526e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65628e14b3c412389f31e5d675d43dc126b84499286f7ba0f1057481900a6fbf3117e24f42c92afbb57008a6a681c88597db8429fce3a8276c45ca01814e3fd71cdc3ef06bd87c1964fed3b959f66067658fe72406ec8d88fed20c2ba39abd8bdc242e76ec0afa460fcc7a6c3e6e5daac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ddf5acc1dd0674b40471e5a95d656f2cb9deae78475e4b53a7095f10bfd839e8061148990fcbfd620f30c76f8d3bf9c918241922329eceec792bfef8bb1b8faf5665fd9cbf962d68f4f2c3b544188ae2f4f5be2722b29f3faacc6ea4b5b27e013a45310b4237cf33968e20077aec071;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbef8f9488801de96eb43b33e0d93e1c09b590c6011dc24d940202942477240165de927d3113e0ad89c8bf9fc1ab1587260da396f22415b364253e1d7600c0624f83c8c660cc2fb8fba9a85babdd7d966296e994b04f35e4744ffab820262926675885e37140ee59a58da94856b7dca8ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a2ea72c70c0897e403a7144f1451f6d7036e2cdc863d9e2d8fe2caa2532080c794e958d44eef6f0b7a7bf0c14df843ae7c8c12c67b8ce940e5df8e3974face37d769b378b90a6e31f940888da3c1eb04fa7189954342e63b6ad224d26c577c14b4602353ae71589f66acca8b4f92b5e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467becb16a93f69a77dc1e4248858cfaf74e7308d88b84b1c86e11f5b9404e5b8b3c9e5d43e15ab23579700e410e8d56bd3b3822b38d11eadee56a1355407958b44de078069a857f37a60e0191be0bfeda3b5edb4d777db7a39e8d6e48469c21240ba676941662a8f48514925ee4434d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16755557923829dce351e1251110108977815b32335c95409d4af4001312e338c9b9f856097328092fc474f5233d051280f91d806b87038eaaabd025c1ad4ccf659e001da7697acf47c84ea4d1e52cad5caf1ead3ca854501b4606f97a8d64e54d2b8826e75d24a51756b9d13d3da92c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aac4abbd81ccb2a7f0611f80648147b06d146b5b9f1839e4a5c6f1f65525e9baf7bec80d42c60008a15b325d86867958981292edb1707414c2dbb6345adf8e68da4806f1b78adedc1f4a7993230f9946e51f2b83a90c7a942b2518afa67ac94e7b5b2f9638bf684da7954e466188d869;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha21cdd3eef6d199bae2357facc0bc377e13abfdfb91e833ac73f5bc38cf4bcd4551e1d3a3bec08d425d41aae4a1ab4a35dbd459dea58bafd33d3fbb3d02a68acf9110e889669450d184a5d3e616547b61c779e92c8682d15f034a10ff6a193d2ed048e59a87d2ace7945b73c7ef378ae0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf04aa7fdc70081491ffbcce3179c328b6ce210f904a58310cb4804f046ecb3a7631040eab9b9a44102dac946ff01b0fcade9cb9e84a7c950b36bf43c08f50f59659760aad7b1b50256b48f308ba36dbfa62209061910c233a18cd082dde826163258d4e973c2aca06eb96f1a6ff949;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h104893d98cd7d993ab2954aaafb4fc5d6bfd7cf653b011e3043f0d33c123b010bf6e190fc673b843234956a296cd8edc551b9ba623163952684a402385618739aa897a55492007ecc7bbeeb5f412161ffab86080121d4307596637df7a144ca398f56206fa7b0dd679b096ab8b65269ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f055b9296f4990842f243db96c7826553702b7c387350bb038d4cf46d80eceadd8edaa3a6effaa4d2544bd850d1057bbe2e8a02af9e760b5f0862e4aedebd8be1a79108ade03c9ee70f73787e372987db06957802c5c561f4e41bbe2b7662fbe05217df5020e4fa16029f5c401eb432;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc358bdc67cbf2781b9278b5978fa1f081bb0389877b1cdea8bdbebea241d7a4d0ebef752051a52213a68db2cf75dfb12fdcef21cf106c20e8f39180b9b0dab0790c0cfb78a373937db641bd6c5579c4856c9a53b552bfcf3d505d86abf59f9fcd764857c7954bf4c1a5e015e3c3bb933b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had79e05e2407455bf4633ad6ee2bf36a1fbe4410404ca7e66708f89f54a623b60815912955356da9e70a9325895d53a8dbc0582caa591a49f82f9858a8f56a18bf47d7d1cc8f78b7337f5b641a5de38cdeeee7b2c867cd7828e592a374a0facae392ed6be39d791f6517ccb2b26dad009;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbf55951e11178f4d88ffa1b0178ba3e019d7e22eb9630ef01ac98d6a15cf542d035a4b4c7f3132872abd416fc7f8cda3fef598f1b9bf0401cbd23ffdb7469f78cd0d4d87feb9c538e123457c757b5ce5172c8631c479371a533d358bb2a4bd614da57f3b93ad22c13e1f37b5ad1bacc5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7632705760d8aa2bb1754dfad7c7f39e75dcdc29fa3d1df8361d06020f036d7c71dac3ac670ca0e153b27d5a932f9a6a46450a94926e267ae7fe423c0f309ed302d1722e68311c00afc4ddb268b7b8b1c35940da29851df1d0d73fe803adaec22b1d2b163ae55ac072c466e8f8ac655c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cbf6df9ce0ec4d86e77b8de681cad46fd0f65eebb4e5102b1a94410b2cf77d3d6ae73dd947ce4f7be9a2a5e7497d122fb70a01a15964ce3fe5f678b34ad01dbe88c5f7133f7cd1476ef93a60da90ed812a2cc0479c1153a725d109c36d8f127879c7c57e11934f990320fc63b6e782e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b08e9274bdb72979ab6007228f4b8f84911cdfb1dd21511b28c9e4479fbe1bfb85ee4efd387095784328f274827bcf0fed17f19c1dbfecda748a11238ac1b83a28a4358a6d63b2e9e9cab6acaa81528d0c69e0229ab49ea534682f76ece8b3a42d8c5adabd2165865fb43eefd0293e57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd8c9b7c971584b609e66ef0532a7df1fb3de10fd62614aa23ea013abd229f393965ba8bf9364cb7b8b7fa202b5be52c32c364fbb6d411a8011acc8bd0232b5ef6e2609cefbe1277df53838fac395ec674a2f210082d279633c3d786c60a434692be914a1697227a87cbb3af3d6ef7e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3acfa037fef6b57a86c0224394e3925a39adeef8f98cf4bcb517a9ae64c63f52885b7a639eb7cf019e047107d504968caffc904cd22e727bca5a1e6d8f169a35508038237a9f178fc4ad9b390210d38c545177134cd3d2008a8eae75cc3a39ae4ec2babe42dccf005361beef74abc71df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa6a8ec7daf6f9b2cb22c2db1e1cb7f0158355e65bcd7b7f5d83c782bbf9d5240aaaaac7b99d95b55d96278726a956ba5a64e28dbe533fc637a5216372f3c125475e59569378777a8f220f1d2c287ee8e49e0b206c96beb5bc5d277a96e54c053fe8b1c3bddddf7369a2b98dd9f162a21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h116412b331c4498f9465b96ac45e715ff3d0a6b8a4e276aeb3f61855ff835310b19c28d432daf641964351ce62df42d675f30578ce3ef484417691962057f4aeb689337ff2d96a8c76375010913edec3a73b338497bdd69a28d838cbfec2af02514ebe7c8eb974da9dadcd16329dba1a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h400c3d6cbc21b68a09aeca42e6ece7fe8541b1d5cbb1e8be6738e1481fcdb1a7aa1bbab8b6b2d25f88bb58f740e4d347454b6478a9563b27f64050e94e476011bbc018aab8008aeb83ed76066cfdf9d8431d9798a8be715ff14ae91062508e1f1f6efcadf752fac83136607f16614919f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb1474c7d5078accf89ff9790760305d0acef7d1c29990695e6ac920127fedb2d3d81b53a7e02e867e621a12959a122e79b514c946c4113545553164146f72aa7eb57e64698f6bb7375d854088b74e8e84e4dc172ffd98fdc8e308eb458c8fdadad9250cdcea3ba32b1de335b584f0d6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h332ea56f30c7cd9e92b006e2aedf2a353d2000adcca857cc056fe1cd275244d9449b98f32de6260a1ec6a4bc230b570cb642e7d4d58ecf90332732afdee3ca31518a9fd3c2b5f3085b32c89fef359e694219e305cb4be2072d686a9dc295e7cab2ae2996866c0f89cd7b6cfda4f636a92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7181a863c35f99d7703024ac6930a83e7aef2192311d3d6120ee1090082a9ac52ebee8d8e82bd66a3a6d9d0e025a01726d3f0fe596d1ec519833a6e4564c7bca73b3774db777c3285c74e22d95c82501d250965282aa0ab2ab4cc54e4743aa8940b15ce12527319863997999e4803b9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16835b5f0df77459159ba3ace74432691d1e3ffbc2ef04cfad299b15110e831fdc5a0a643e4e60f6ec4eef04a71fb2deeffb71f7e40862c290ea690fb4a686c450704c07e2532d50a2d42f382e205a9b3d4f5d502636c9361efaf5d1eb9203e6ff94c90ac587bb1c0a65c8e96dd326c62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23125059193275e30b9d46ca05f3fb584a63fd029009ca47f6a2ce2cbd8655436b39a3e3f883c44f743414428ea1377f96ac6a65543e7930e274d329f17bca1a37f74a82527ab44f047b4c7cb11f38fb74a3e83f35298362a3f2ea60d71575dfa5fdc5a02ecacf354c9a08bbdc95cf30;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf801dbc3a147aaf8a6832ef67974711c8ffac076c34880c2c7a6a6492fa2ba277d11f4e7d27270c8ed6d37e28a8a7519c9cf07cbfb2c50e4f29b6291185acb34b5727ef7574311a84d7dc65bec3b79168ca2ab55c67dac95fa5cc41ba6511dbe71ab3a2a77817466a0554271c03ed764;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc809ba89921de9725b0f309650205c337735554343cc22e6510c8c5e70cdfb2da189a692b7653963b43ef4541b61da1cb752504cecebd60b66159cf20df40f5e72926d1896bfcaf34f97809121f90f653bd5d2aa6c7a627bcc0822b652cfec0b4a7fe3178c8363b7e6c0af6d9a7386df9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde93ad9a703afa2473fdb586daf69bb1ef27eaf936196a835270f955a6189e34c865daa2dc8d024db142e41ffab3f6917c8b8fb870281e797cadb048a5e56bc0faca59cb374e6829e12c4fb12a267bbb00c2b2f75aed0f5389afd34ba6fc160280716844500b36985dfc70fc3ac256999;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c8b2eef37c4dd610ba3a9104be37a1c02432f4b65de52633c5f1eb4d2e482dab9a6f41788314e8240a0bcb47438865bd9645992c50e6a94d5e4d9b91c75f51770f609d28feca2803ff06155c044c90d194ea18dc8ec292015ceef878aeedbb0bfceb2224fd395220f3a672e46b44f52d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc23c3cb3e7cfdc42d6ac08b0363b2526e2519f451ee6313fb910b48e6009ba046eb815502f067263537f5ef21c88a5c14e72124aeb22bf50e0c302c84b45756bf6e321d04627eb25a6f9b91a695da6d82f367dab8c07a8f3f7c28c7b1366e52d2b36c6bbbec3706c55eaf8858b2e8d76f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6726f30f0ad75d932f7f46a79ffc3cc8d74b5faeb22ae5a2fefa53586aab007759aa44051643de5c0b0f8453095f74ad2fc59a999c9ed4367b40d86d5d9aca91fd6cb85ad59338ebe9a9ceffbbc6c38f2920b5b0bcd47ea6e58853b99f938ec42ff606f0a14df0853e379a6f5e381bb2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ca6249fba87264a63d10432e259e4af0d1315e3ca8f4a29e0b0f1b8ba91f3d5caa90c6677046b7c93447b78ca5482824dc3632f275a63defc4904abc0e119e9547bdf593c03840b6bea4b75ff040774fa94d54745d5bc91b82c180fe15392b04ce48803479e1af3956521295d50c02f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ffccec67d1c1449d12eed0a3b91eaa66c0706592a6bcf4f66a667fcbbf76770c9910009f51332a9083cfe7585397f5d1a4254efa8cae3d55386fea2cd4e543d68b281e4e5940a6fe0d13bb3c01b9947b14f1966ac4261d31df7e7ca2f1074201cc89cedb424455fe7b2678b684999df4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6eb250da24d41e4a956df90815124f262b50cd5ee2f479391c0332b5c37bdc8f2371125887b788095b47a0b958287495dfad4fa9fa192a96c82a8ac39b50a857a7b00ff2ff8874fa7a338a69d98e9b38816a1400a43612d02a45fdbd8fa2b54c8a0a4845afeadcc2b3cb0854b09a51bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he71e2a04f6af00b4b12db0fbbc27c349c3a871a28fe0f0a85731aaac41e6a319a9e5942939fcd730f1718880db4a66516f106a116579f54102b8b56e45d52650deaca4c750098dfef859819c25cb63ea1e8990e6400242a347113edc2651122b4b28f8b527cdfff953dc8649291baa7d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h263931fca21e2038adf85fc8d4ad05d28ece132da677ea497c008510d39bdc5bcc0a4b29da5cc54ef276db2790ea142e2f92d0e7ceb22f3a7c03c4423fb08392ac93df8ce5760351ae11a2e48283446d670db5d2a1af46eaa63ebc29537479051b9d9170c9807b4b58c40abf40fad7e3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf529dce657074d668e2e0e08e2881205b0ef33baba0a527ab8562260e875e9485743ccca676c6c5611c92d610d519741f7f46f765032b9da7e0b44e7f003dbfb2aad01c54c996c96b734d13e8634a27838988f7a9aba65d3c9413961a772f7201016a4a63422a40aa8f3d2d2d26d673fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h430f0e89ac2b5340b6d511ab04f0a966aee93eeec3991cef17351cfccec7fd2c16646d195f56de8a25a5434500b6d82cc013f11c24c71e6547d63bac12f02e114d9ab639192857b4a356f4855280dc6542c6362c6a01b45479ab63aca9b290cb7a3517327a9e903501f6b0505b9d1bd03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6104e62f5e3aaab11e4093c4ca59bffb95267b43cc46f80c9ff9e77c3a9d27528e05d9c9e4cbba7ded4f28e2c5a9be8154bb988daacf80adf4af3cfd35741819ec722b5e1cea0848fd8a006bf8e3584959250ccd167cdb0f5b50094ae74211a61d33e2ee64d238c332e2fe89a3ce2182;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ed3f39708fd7a017aa88c7436e7e49fd3ef20cb67e6d407f940eacecba79fd87c61f0f1278b274d7add014a5cbaa9d5c58efc0a9185975ab3e92148f36172091b392bf8d0237a15e908ed251ee410c9497f7d3a90f28cc6226e81e19eebaf0ac477711faac0054d5cc3c7c47eae3e863;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b9fe5492072d7372533fa46dfc2a073c7a64ff935e7f60fa62114391a4c7848e1de6ffcb037f673244bf18981e9665f6acf26100e176749ec4c3de8232a54259d60b5847344fa75081c4799cae4b1b2a25673dffc28849356e8968f0738019424a7b29eb7b61256c198afe320df49cc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3728062ec1ec2f166e7ecee5a3804b59f7d8f986c8ccd7e868b8a90b132a2da92fff5823795466d656cf8a6a3507b5bd89d5595763e6ed866c41eafeb449b4512a28254e198ee17e2e3f5af3f171ad7324d1ff2306ffc9572f15645f71a339d8798abe1818ae331304b4c75ab69c016f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41846304fb81f152517f5b6736e9b922a5d1350a92834f7ce504aceb24fa86bd19dd13c7a7c228e4894cbd7c22d64a585bfece42618a34e1945af7cf2575c68a0fbaa1ab591d87fe19a8493cb20a6b8cb662da5d294f7ffb0b165b248749b35762d245c263e41c9cdf131907f55151038;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c733b948307c4c68dc593700adef6c58ce005af8889c458ca1344ae55eb25f8a16e153838446cee971047124f09634928b888a9e6004036222535400097c4bf4e23a9aa8a36835611613863cece69ac16247848fd014c08922c953531adacc578f5b96c16492b7ba8aac39c55d768f6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb071c96a1d51c134cfa4bd8deeb539ae3060ed92d13a95810e5dc625d71bfa65793f8106c5e68df62650ad35bd682693eb606f1c98a087dc1cbce5bf5fed8ce6a513ecb83d00bba7c046b0a1b030057e7aa2d98c88cb9fd59faac940f9b39130a134dd35e26db885d4bcf350aea5790e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e5d941c6ef6f40051ca30945935b991ec8e822dd6a7553a69dcaa2398e2a40f774b73dd48d317c962b08b40e93733f0c638e166a1a20b6eb740cb9f983537fb7753091653e1758ff4726c9efd3bc4883652fbcb51d71ce58accc36718f1ba1aad6207e069f4477159668dab8843e8fe8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ae3cbeaf07460e5f5808ffac55bbdba68f8d99996e3f71c6972df40ab9e01fd223aebf1fc4735e4ef206f5141fe51f945d3d8bbcd84a2b04ec5d0942028e52c7562a09437063afd6c9fc8121483a4718ac7880e4f40828028d28dd2f765c2178927677d0b3fbcd339243b8cc5abfac7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf0780421ec9f210efb39dc4a4ee4302a956348c0b0386f85cf1af67eb6c837cae19a81d0588f8e9d6c4b6d3043b5b79cd9e7a0cadcc286487c864cd74bad53e56a8e8720967e64213b232c46a279bfcbe84792e1221eec194026576df02bb10d29320ac94fb1bf64b4f6bdcc5465d050;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ee6d6e9d53dac09264fdce0d25841fd4525d409b2f10cffd474c84b1d1a16ab5c618e408a556c6322bdd60c76feeffee6ce7007d4837a09298cc34cb27040b2dc53d486ab6a89be4e78926db0ea60fa5a9bfc142d3f513e1ef90a8896dbca28ec00faf8f4a571d4a3b87559dcc0c19b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h362ef743cb7d08371d36413e063367e31afc74ac8d2b32efa3fa3b1f0ce18b91f32fd2f9ede1f3f97a244de972c437a255db0161fe8838e75d2a0e7c5f492b7d365855444063694d788ac4fc262814c13983095d087d5c07b4edef8c55379c33aa85ee6393162c5e6709c28a321cd89b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae868a7add0cda1886391d7f3391398756c45056dc5f6902d183ed208dc3f2581a48744b45dc4be971899e535687997c08e497c34d2a8c20977b9b7d689486e1a9ca9ef0934c9bae565fcd9af2ca5ce775ccdf60c1b92cdcf5dd44fa336711f0d190aec8483655dda84e649ce9073db4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42021c4fd94dd25cdaede5d628093ba8f07dd129b5b702730e62a6109a720bda5c20696c45bfc21a56d0bee46e16d543a55e5dd9c2a10b036c8b02b6470f7bfd5027d8b566ff8fc71eb07e162e4116c410785f908c855b0e3b3ed19ff6dd8b81799872f6d0ebfc16a0b2733a5c9c6e8b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e4d51e329f30a2cdfb0cccd6b95cd30be3939bc53c7ed7c4689a077027c88289e226b35c5ae8c89bfc8610c493bbbf65ebfc0d07ac87ff93e43baa0a0d548c3b1ca412a3336b9a2792dc5be765ef0d8d0acaf2ff79ed34b51946983530fae7dbfc2ad475eec769acfdc49af29efecffd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6679e4ee83b7ba00eb6d3444bb81cb6dcd73ef7363e8fbee8b4017334bf056ed9d745565038b26d60f8a62032f0a89ae20cb590dd1cda2a3a974191447ee8274f642b948cabe2cd19577646b8b2897c2cc19f874799917e5ecf5394ded9573a82bc1cf2f9c62c15ccf4a041247b3576b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f06a564e0156446e0a26fe28f88a7b2bcfc8242f3f6c575d1c9037bb93399b02f4166e6ac3e6017e110918164fb7522befcce10fdd454bd2b41d323fa8c3d10d046bfd3a40e348a4ec05d114b216b4f4fc190162ebe0811ecc68298e51ad94aedab17f61fb600fed7c10dd4bc66a29d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eaef6a70bc3b7f2b016ecb8c3f2110b7d6623e8b55244fa62bc515e6b39a541aae999fd6b7e5f09d0dfdade083d482dc67d307544ea3e7d4ac848c1f9aa2684c6976f914779edbcb19a7a38905ea7417711af42fd53be509b5adfcb314250d18bddfa77d2f79427815f7e8509f549223;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18a1a362f8e2791aad7d7cea0f002fb6565e6d90b721d548b15cd7c466500a1d5eceb80145bdeb261dbccb6ce786177a1764e4dc61de664c64920408e69db7082a974acf02b3e8341bb2781d6f4b16ad263bf8a952db92c817d6410137c2bec66cf19fc5dcf55adfea7752fb241bc5c46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ee07943ba5f4e618b00d1d67661ccd060cad701d7cc68e1e9df3671e53daf27005b0f9e37184510e5c15461b30953daa8b04d01045a3980fc29b81f4a252d219457d12c3c5b7a7966a5bb7da19c9b563018c59931ebd51bc2c80fdfd1e6c65a58b19939707f5d00563e03a735efba264;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbaa25bd7ee57b4ec31aa6f5f50336298b8046cc744aa5a8e3e687efc9cf6bee799212a2a0d5a2fb612ae0fa437f45180f8383bf76bfa7ceff0731f626d105c6289064eeb0e7bf13238b33c96b2da597adde84d7fc8acb60e0b10495c8dba58b73ad493525d0a0a5e8bdea4fb52aeb33fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3345f81656671a55b78d113a92d950d07976751ffa140c9dfc937107d81e571fc8d18e8cf17a849b4d2e54132f9ae1dbb4c8688eb5f74ba175635cec848ee964be3a2ad10fa6c9754ed91da6c430dfd4aef27d1499333d62dc1e2530522112e5bcdd454a4af5a5f3031f77b81f062bb14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1740ac1493770e1844b00b8ea660c3139b04653ba5174d8f5e50f907ecdd13dab2110f039c213f060f4a5f569c3bf1a4a3759fa7bb126651628592e47e8db474995c3193fe6a9aba16e4a20d8b7ae13ab2c29a6f2d83f905097ece864c6b00df6308d5f2d8d5a79bd34c5aef347bbeba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73bf63172ad50d71bcc46b9278a381d5644cab4ab3c98bf7fa4e23638b19270587fe9c05e64c8759a9165cfb3a7c6d44d33caf86149619ae489e36201b155d42e0c322be682e8a35cad37ae9f9f561e2c7c1c628368bed157c424c40346f4a4381e4049a23bbb48f873b90f435e72072a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfe1b594e96dd3d153be42206d22e8046df6e110b824bc77b9b0875a5f1b0555b312571348a051a00d3b9ce24d7c408b92577435d9566568ad82541ef358d7c8a1b1203e278f96ebe062e93572b2ba49c21a24802edef84ba3ae31395c1ebc53bd5e6e6a29374ed214b3773bf9bfcc9a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef03a981dcb3948f731b04e3acffbf8b2a40f1af75e7f8e48ed9eb278adaf3eab9a741264ff938bb435c242e077767a499ab41c215af8afd0cea5045cc77095b56998e3f2e56275a9ff30821641f45cce1d404c6433ec4be9170d89fed786637c5d93b825f97e3e4c1565635d060ed333;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h326dd1cdfb2bd7cf0824fc8e5928a2e2720ee07cc3532e38a45b4ed719909425db6663be1c03668a0b84542d71eab2631f1f8f53054bca0bec7f2d42d7ad0c7fbdc7afc5e2d2a76e26816e83eb9f3406739916f31db6b7a78b074e413c5c641767f50a50be8b9eb7d03214f0ddeee9bbf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eeec32d9d9c27a740aaac37f19685caa02422573f7c748c566471a4c99d46218ac8cdbb99f79ab1a4523f26d686679e615c30bc9991cb28a2a7eaccbb9dc14b69e41474ef552542f88b7f1ba787c4f4871a3ba968bce916d5cf0d7851c93695d9e60a72eab6c54681061d0d2eec7dd9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1c0cbe97792f5bcf1ce2972c8c47ada65e5580226ac9a6a7cdf8f68034a2ef643085020f82e8ca3909ee061b6d74259ea6a699a3fabcc6d8c09bc1a9bc8731060b276895292bda3ffb6ae9678d34762657cd9ea9914876c0cb4935bed357171be17f4bd1bd2e6ea84560bc335376921c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he99c245254f2c9e4ee6afbf9dc047eb3923f5da8307712ddd46d0cc105e6470646e24d31c2868c21fbd171f55832ee0af1e4200edebff2f8c4aa4c15f0ff77ccbd4681a59706228033001973deecfc3c794fbfbb6517231ec2e51b9aecc1dc42be751a8c384bf9f0bbc474e2b1dcd530d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37c2d82a93cb89e0b63db3ae1755364ff197f886eee40b218836cc1aeaf8ae8be2eef6d300c6c4176e1822f5924628523d3f023765a91bafff9a4654bd35052950fcbe7b91ced21c08d6396f774fc84ce3ed837ac7f658a3b853e9092af3bac8e10249b1ed04768d4ce8f8674d74250c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf046d37d386ac48831ba42b0090381a6005bb5421eef6d14e6dba0f207ab210f5c14010b80278345988ee1f6230b08ec738a9e719f8300b572d655e2af745ec31bf94ec6e82d181c86db2511566929f5a1730a7171b28f862535c627871fb842420f06900d18144c5e19527768ee70c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44800269b11ca544726de306dfa79f84d8139f688a1388928db1ce8a5a415ac2a916ed8c0aa5eb0cbd2ec777f01cb64db921bfcd44421aff4f54366694d27cd909d07d621bce15cbc63367b0b3866994cabe9d093e638ceca6077f4a3256b2e2ae0208b85fa509a82e2b4da9e12d03ebd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h834bafec5c4c533162a51b2e1bef2c1c83a2de897ae0c9792ea29964e41fa776718440e8f84ccdec31b38cab26a168a43b3a6a283a8728d2e45c9b6ed0356ad2cf8c62b16c1424adebde1497fd8a4b87ce494013343670a191eef13588ec3dd50ce37d7519ea3814009f7f0fa81ac9008;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b1992597a95b8c49727561cab54a904e1b3db5e5aa9a057d31a814c9f72366fc194cffd0bf3182d9b9f0b2e619afb382ddfde3aa2538939d67bb2ba7000813c8c4a66cbac6e4bfe63b633b30f1723d63dd450a68a9299fafa07178ad03320e00c3565b7b344a645a5e68424666aa4ea8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7739798e0105f4c4606c4470072126b6a3cd93beed2c8bef2f7b1947c75a6b0dee62e72bf59221299c6f8505209462f93fbc51194c76675794ce9d734f3fe1263f9437c7a4cdb0086a76618e6b8140b83e293acb3ea79fedab4f429686c98d87d3264110d777cb6a5183f40545329ea9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb81cc6088338f4ef73caf725218097e269c9f169ae749ce1cea42989e5596d376ee7b338934a15c48b5303b476452942e0f366f93bd7079093a8ff30121f0f8d2534024e43156555ac2e3705a9a81cefa1be3579acbcbdcbef0c77b87ff3871d1024802afd71f133832c542f0f35ae83b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he01ace0365fbd7b3ce9563e02b0ffd0a16fc2d5c307eeabc55bc07bec8a9ebada696b4e333283087513a3e6d7db13843a4cdd239f5d832c685528648e56f871eb9e91b6d6f50f8b7b16c59642abfb521a6e84f7940cc16a473dd502cb7752ca06ed04c90672aba80635acc84b7354eff9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d78e65a84502664ccebfaef32105042b1538db196b0afcb1d6134a4f2f58af62ded16cc306d841232a1028c4256674e25474f0a4b7a90cb8c172e82678f962667540a038154caa9a9f871f676231ccf068a198f707009216802b3400782c666f37de7a7901f65fa8c1b879d6d6287b06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc248bf2da55c53101a74a34024a545887af60042c8189e7a5a10ffb7a666f692b3a33795755cdc4a9eb17154c1925dc767fcb22ddf0d7b24b555367953a0c44b9c9209870a2f67149167d97fb23d16a2e8f11f1b930593dc573bd5e962476c07be4b1f35df94c22aa319a5b5cfa88f208;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd2dca21c444ea48cd46699d9611fc42c3f69ec5557a7292da22281e1be7047e7df3385b3b13346fba5fa714b7ce73d2cdbc0118423659673c8c76c33402bd06a58609ce58d802f3ea7780f5b1bffd62f355196fa73147298af9ad2e9ca9af86156f81ccdaeefbda7479f515212358615;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61cc416aee8cf862f916508d531f4fe8f69999ad29be1eadc1bbc7ca9babf0fe8045ec7955ae1609d59e149c64efca0a50d5263c0747558b2d889b486205e726d8d23ea3a9d78981e311593bdc519c3fd65f416a2dac3f587f7a62d60e3d8c4d8f457cebeae0f8a31f591704affdb8cc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha81c9e7a4685646a001bd8b32a4ad3d53befb30d325dd5e7a6b1bfdc906c1571c9153a993180faf330cae89b2d84526a775402a65e89ffec1ad658d3616882b8294064f973bdaf037c2f2974c5db0a5aec4fe7250ae28a103b601afb9582646bb5db126cde21e3a0d1130181bbf574741;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf275c5670b8d5ba54ecc5257f0738f9f404c032d2eeaa34b5caf0463868825ccba921631123a603b38ca4c1eadd34cc4edecf19e30a69c40e2716b36a254ac84239c81c7fd446e2375f2c83b21e4ee12515c998213dbb464fb3ca5a8a897746fe806f60bc56b0110bf500396caa34de7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75372f3cc0e5dea27d884db78122459ccb19e0f752a9e1cb76a7701c5a4c6259685c3e687bbfd26775086391efe569322d9aecf478b940fa3ddc111926d42c72d4a642d19bdd86e53684e59f625c4da1806b5fef36ef18d7b4a97bff6b4b7aceae6574ec7af1b92d9a4c58d4b50b98ca8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h299226b9620022d00baf77f09068cfaca4a2750ac8505e4533c843b6c646f2e695d3f53cb71c629740e98dce7f8dd6fcc70c6e41117d69a23128250c2748f1c1c6a41542fabf9053e3410ee405d4c3f71e880cc8d03ee3761758acda47e3e876c4763f3a42ac3ee67a01590415eb4105d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e3c672c44ec28f108e2d006d96e86eacd0c54d28d79f0eba74fceb454bb87b03be9557928edc77c40ee61bbe1fb6b756ddc245053fc33e49c9d4dcc294fceed4a5fd595a1d51893b6e9e54566b836885218b757174ec4df9e2f2313c2204ebce9084311009cb7fd84cbaedf229908368;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23c8d80a56de416e74dabe104f9492acb9ddab46e9bb8dd1a6f6d89d1b6fb02ccd9849b5b624bcd7b7770a8065a9ddb6a2e693c0f5cb6ce53ed89ce9a187f7f1f89d4a8b367400a977dabebfa4decbb771d13bd6cfe6f5204c4f16aaed2b2e6af530012a1586d23c22359ca218334533e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3379cf7234bbcc5a2fab66e330c72998bfa74d14b5a2d7757a3754eea042fac3de1ca1b600f44dc986647f01fa3c3c6c2a8853e29d127866c219eee209702d4b2c9ce0c90efa50f2bb0a57a0bc6dc9155655dd36a149900dcf356fc58aff48270c5d1fc0652af9c346cb05c38e1200eb8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8526257df88dc2297bf1afcce1d9185c6f5a8a92f90d2e5c15ccf4cc4568e5ba1c048194019f6d31576e8b715740a1a82fe558aa9e6a3a646296f114bf48bf9e9320c043eb277174da61c649aeb2bc9b6aba77cf35c33ad427e68cc3f343b3a690384233821ea09a8283e96d5a44c72a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87741630785bac2d305312d312c97dbc9e90480f4b14332381351e931a3c0cbe43c5e9c2995c971f8a4c1577a58a8a3bcfaf03bbe2bd1cc8e8d5bf979da172036320c82171676564f557f9fb12cfd4da4405a33c8a44023d422e8b6c82bd31bf9a9dc58abf424f0e85f4425d82e5c5b65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bdf0605617b97467b86c45b830fa9133e176493600162c1db5d129d3037f8c931eb0b686ed8dba78d2585b4bcf4f7a96dc831726c9cd935f1c2e98d160f4575b69ea3c61dfb8f8256ef98aee5a1adc74e8976385a9b6175c6301467e0f2572f95ea8a8a2c623ceb3432516e519d466e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2ed6285229128c668d729e1d2286abdbd5c3f35f610cd594ecade599b285b3492ce974b6e83829b4e02ce77b63d54595355398063ca03d4a2e7beefeb82b8dfe10395bdf852d507efc76f9f9d026f87386487c00ea1fffe93c99a49660d5fa99de8118a79a84a516c65462daa2a49f5d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4934bb9296f94315dfd7bf8ca6a21c17c8ecd66718c2723017c878c6cb03d22ce7b76f7090664b3d1b3d5b165eb141dc065cebbbaa1dd0d79c872ed33842b0a59317b50aff8d124a945d7af12217facfcde1e416f2cb0530498e489b15ef1b58cff8150f19d19739187c65b6085c9d0c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92fd21195b9f86cbc3ff6811ae77f3f02c82e679596289f3d4e24302f31e8eb825989836b5ae910467c7a575a27956452b1739a4edca0325daac96a5f03e1f9f9b932ad4f4cb58002a2a85f738654db01199ce6631a490c7dbe513deb780abee4f1eb9b5a017a8dedcc58ba6d4073d551;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h852e9361de87cb1691a34b5e36c31db3a2e697729496b6863b906279c692fa1b58293299974abbacb4dced807cf1bb71b82033d6def066bba48d0e91ac41706dd75bdd6d51de0d038eee106f85af2a0b3f978afd8b438388c11a45684d24882bb5a9497c4a380214c6361504649f32e6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7721198729c15228577cbe4345849e83410dab075d700dd519237c1022352cb1b34811ef796bb3203d665fa7a52494dd6c9e8428d2083b10ceb8cbeb47fcde00bf27bc85bf610f32234d675bcc07624b7198150222cfbca4c8290af207e306e67bf052c243a013b20da8596c05dec6aa5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3ace6e687fcb322a83aba94ab7d7515c0394b898cc94fbe50097f0d4de6de8ee847d4b62153995a29de694e0b81fbe5610e740967502245bfd5a47ac51abda95d7954060cb1855d511b92494807fa22b35dd802d93b7863345b519801276ecf1e205e7e0e4785016d6354cd12835d195;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h161243c3f5a6f63f20bf3f01e505dc909f95cfa0dcd5639e5ecb20a6191098e7055c1d224574d18b8cfe400fffbb2f1a706da864f1f896257285550471467eb1e888ff992805f76b2d9bf685fe917a26d6f3ae235a47bb6d1a0067017dd938fe9f27ea1f60770cfb5668b71a2b9d737c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9632d0e009af50b2805644e7693ce67497c13d361fd6e94d41d5fba9deb9505eb11485d4b4e09b684c4f83554aee30e2afba52250821f7437e4e59a4295b86736ba9a2ebf1b841a340ad1f330d6eea036e9f39cfd3dcea0a15fd8a32d5f139a5c153707da1a5debafcd8c5fff008f7419;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6b16b89a864c52a980c4c01158d80bfbf78635a4ee369649c84268f793b4263e1c7840b88da31bd880eb92e230751a58a34aab38022f6cd8aeb1a2c0160b8294ec73706e812ae521a8f832ce3d3a234233b32b93e94a6f330b879bf3985f9b17cced4f998d07f2c96c2ff510c7e6e910;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58e8fc1b6aa5b1121b182fd30db64085845a77dd8ff7f1ee536ca43e3cf91aa60a632c286bbd03e349f0a927c0178cee238bcdd2b7cda91d2dc497c2f9e87236811d29b346b2cff78741ac85cc914064e13ddd1b576f2fd76e9355f3b9edb0a1f41a447fd5dd7e71eaeae1b5f6a3526fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d7c4d1fdbe5938adbb1c6056932c1d3ff09538d64cd3176deff593ec5cd4b5e3fa7f7f5287001822ce07ba6db18b302ff687d8752a1a4de31ecf88436112ef7650fbf3bd8711ef98c4afd718b69de7ea818eb1d8df57a0fa158a126d5726e90662781847b07813cb3537e65ad9a29879;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8abe29f2134da517f22482cbec4d0db93ed7b2065807d13b74430bf7c0869b9750d37136336fcc48c395889ab5f49fe154cbff851cc8175ead41cce5a2144d4dd5afb7e6b30ab35946753da40292932c5a0b12196758b363d91049474f7810d0f685ae926ecced4c7a40c8b76233d91a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1eb4e955a2b2ce2c5147f41796ee0dd3a76c3d4e7867a0d4093265cb2ece24804e1c6e8443cd39796e345fcf1e5d1483468277ccabedcc34aff5a6e50f7607af352f0d15de99d8f8488350f8c6fc11fcdc8877f47f65cedbb8a776f35c2c7f0763c6371045d2498ad19779eaacaaf863;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f224a1e09fb44c1cf70c602fb5c8111d7854b10521113f23d14523e3abef8ca7fe731050836c3b323aced6b4e8195effaae324908594712a0edea73e8efe0c1d621c45536cd6637637806c8e43b15357b4454c655e639f33a57a5bc13c381c71c2c5aca94104d1cff0ba9fffd75de7a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13fe98b70fa142f87efadb927d27280e3bbd006afb5ac564c25710b09d590869b4987872290011f59b2ffdf3f19e313debafbf79e2adc601e1dd006e121cde696e64cc23fa17118f9c477391a7634a1142d2edf1e7916ff135701b18710b9e111962506ce65c0d6344dbae3b54706dce0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9da90a9ebf883985da2fa7ec31b89ea92424edb8c367e64906da67d50fe53edb2d351b9df62d6a0fcf21176048c868129fa19716473e7ced2e20c49b787232020f28f96e2884b3906304ed0058732fcce6e46b03c4d4b6009da91cb311db29a0345442373404e594db8863f96da13d245;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc84a4f25e9080a67c60bcd75f5068c8c268012873a1133ab787c2f1d0f768502c7e9a388443b4dd7fea8d52982d8a68b130c5a5fa5799336ac9b580bf8db444a95dddef515d87a2ac0d0406ecec795a45cd806a3ebc07eace9f5311961038b817cf60b529d11708dd34a908272bceb006;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3988761c4db06f87a895d88b48bb467ffa164911a1a2ec1d09880814b7cf3c518c459deb852d494b85232e1a5d002d37259b86830cb89c79710f4e86f54cc58cd81431ddba211f86020fc4e236eed4043502967e96c5b08ce8f0a31bf5d6b5473cb558fb640fc5c379693fe6a339ad5e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h491214e605eb50082258fe69b673961ac5f1b1abc31c501c95266908ce0120154c25f77abf51eadf8b86db863a5d243c8dc89499a6609883df9a1cf8fdf525054e63598aa61f470471cc08ab383f831c89536be98b2826829e4fa8023b3464a9f441a5b612facdfff393cdce58925defe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb46e05c166678ce992954f4b2477cdeaf9ea7d6bc4f4f8ea93c816121560cbf68a30aea06d635a72b7cf038f4b4c56b921522d3781cee321d4234f9f99c03de4c64bba890889133c6f3a2befa30be62464d7218d66f73f6718900113769bc950a978e21c126877031526447ca7beac0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc52d8087e98fd57bace46bb12ac53ac4994818c1364912fa037e324cffc011d452dcf452c4f76a738e61bc12afee7e940b10fb7bdf75fd10637e0770a1f493a29c1f372fbac2284fbd2280db1128a15bf9ea7d0f304cbf32c7828595d979da160e3bbaa29627f8798f5af4fb920b42ab9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h270fd8a00758f14a3b95e21870b32fbfd14c64fd14e47d3f681746983cb31794e49e82a3303bdf76719721a5e90bd8405c72eccef04bfa6e4fcea38505900cc68f22179fffe3f3876920508f05ffd20003d328a608bb04de27cd6dc01202935d9f03e48acb7509dc1c8521335a917caed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1567ca012f9c2e8772a51707017302d9712c2f9cec42d0417ac054669ce1f6f2b39badd66817df3bbf4ea403223eb5466a598233f157eb921348316d4a5c063e8572f8447d6254cd041326d39f158fbbfff283cf6c993f1aa77f149b0257d6210b180a6f0c3262a0ab2066bc38fcc0694;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30d1a607e14d3e2aa5a5f6540866f25914e2aeb402ca96c2e83b02ef5ef00ec6b1e01da7faafe73b3cd67bbb21a19655b0b5ceabd9133074fca5268c458d838fa7c7a33416b02aac136ba84486c08c3447acaa29898e285c2aac18b6a62a6df22696a9cb2dd178f5134acbbd064357606;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8b628d3ee23c39ebf645bce3c6158eced45612162ecd3f21f3b4c812206636d54badba840dc872048b73302209d80e47319af57affb39193ed0b03660430c0c2fde55574bbdea9724c6fa6b39bfd17f42aeaf116ffc53ba3d4aed4f13e1641b17e65b7fe61659d5e1de7e2d0ec5eecb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9a08698d077ad85fce0f295ce9806629fa6b16087231ef4ab50d555a785a72b4af2085ce619a5ca23d25e2449846166ecb85af7bd45cf14680a0476ad690176e263de31c21df0d4003ef1c2ca6e4aa88de379b4a3f858a3015199be13d8f154ca0a832f1bb009d5cf7369c73a2b608e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b1e12e7c628a6997031db38a02b26663d5cfb0db2ce5aca655c20a23dde379bd3511ff19704c15141420f9f58c132746b0618e1b1f11853835922e72e3ef20735e3fef14f5f74fe833e63d15562f7c941386284f099d6e25f74c3faa8e2f20050997993707c4a1c395c7ad979f6baff9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbd9bd06c4190271a8df3815efc66d2f4cfc04a587e0172f7e92f2f1d383fccb271f28b8eb2e4512e8f3a2771cc8c0bd2a09726bce479e3774ed2f53c4655e2747807c0bab0c7d51e979a02cb1666e4eff08953c65f036464358560938256abfea226de4552b4cb0c60a72ef95d6ae774;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde27b86d6407b3fa1d0317764b87fcab23c7f410c450460a19dca5d13988befe130ce7a80d4e8b2081506ba2cdd30e06849cd7850ecdaa8043c7704d733d14f9b20886f89b960327ff51bbe494edcdd45afabe17cc3e76b60936a6859a67f27e66d1e6583470297bc07789314239783d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cd7363ca52f98a23a14a30823cdaa1e2c020403803eacd6e64df9740cbbd8026ef485bbfe1cde91ce4041da6be52904c42c75524009c2698df530884cec77a68d97c01ac7fab1971dd969b4302912a44d6b58ed8c5bca8691d462962e137eaba6b9cc0e8d4ca11c56edbdd65d7e11007;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeffb257bdf01cdce27c9690ae90e389b197ab509310975ecf1eeb97246d359f0cfca032e5d98f3649856a0bc9b12674d3b3314760fd8f51ba6d0b6364075d194217a2eced46e64982675c47ea3f6c6c793ecde66a4d11ce813d565647570ae9f80f2242c605632144f51d878023050f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed839b657148d3058aa698c395cfa30231d46245b23ce65c7d877acbb3b02c89fefca4296225027f0b7eb57a28a9136db70ecd77b06785c21cbbad2980d3600b9ea56c8f6c9cb31dbcbd1026bf4fc611af8e964886162b583780af6a9eac5b495bcb800e8d6cd4901abd200493560b380;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h271d4c7150653fdadc131f8a74a35ced516529a741bc910c4c34560b564a45dbe266c0b36eceec585376b7d77ef667471ea0517005b1db4caff0b07e268c0e43d9a4ea0b6e073fb34d2f788dd928d3b030d3132892da82bedcb0d2ffe736270eb6f3d9bffdaaf9ed203fe5c62f199ae72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf365b1fa1a92f99a5a279b9e4cf6fae87b14831fadd165631e82a964598d875c4b01440bb8f15f353ed0c5cdfe8942c22e2e667104dbdbd63aaf6ee008114efe8fc6ab37378ec38a5ec540f6e4870905cd84452de3fa684754b38e5660b38fdd68d3754ba830930c756d494afb2483a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h541e991051f8d1d39fc0e3daccf0ab16252a1efe8324af2715357b87868e48cc93614a251563dc37e8bee947807f7af2f6ea98a20d0a7bfd12b2121b6364000bdd734a2f7faa445f02eeb894b310ae3ec79c509213dc106136933a3619367214f4157c731d846e75a8907f2832ba4e083;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3729238fea303238ff947ce524f0fa626a4a7660ea71a47620c1c7ae25dfef4f2568c5cd1562c27af2c10077859994428dbd1838a597d04489613fe789be0ba7f4eecf324ba6243793c4f4274e5e41136a5f4f37aab145c804939d4a641a8d9d867b50b45e7926dd725547c1bdfb93d9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5478aa8fa0a6f59cd538bbed9303733104faef7407dca23fd5ea510abe341fd780cc05348f030299930af3b8a8844793e1788482b5d784faab15a5bddcbbb0a7fb19e6203685ebf7f74f43062ad28f96955edfbab5455eda4998dcb781e3a741caaf1df718e285dcb8b401f319bf7a875;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb11b03f6de39e8acf20f030e1dafcd8c91b0a83a1c4721239133a39685f089cc97a3113f0e7515967c81f1c8bc286c386ee5010de1d4df2253ebac1388a722fad1ec2de578e483771347df8de98d452f0448d1dacd9809309f6abdd97893ff85922697abca048c5620199c44f0bd9737e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf421a9888daf1628831c3301347277dce8be7ba00a97488ef0bccb5094b3d8060e942bcf0686bdc329f202c96fd7c0440c4f6e7882c6fa5917dc7dbe4a637bfa405364d94001b142984e4de3d7510dd7f9d0bb803ef55d047e30c642124402dcb1db46b9369737b0cc5ca600ccc66661d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f15f88129ce102dfacd0df36cc9e36164ccd5f635523b5b39bd5cb213ee11407aba6d0e62608308f597494aec4887661205c713ea4158a62674fd700facd0fc730b22006d3549b0eab64eb1c05b9286168c7ccc230134147d24928a6cd5291fc9c0aeafe514d9cc994d5f8bb3306986b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b5034baab2841889c0345850cc2bf371d21e874fd33164fc0dbd2662900555462ab8b5725dd8d93864f8abbd734e39aed64b8bd892c4b2fd0d6798cd30a1fcec71d09e2668d6c6593a6d9b07e17d76a1d38664e6d6bc3ad921fcb8be0a8f039835f124f95e7c9709673f35537da70c09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a7a7fc08bc898914767c5b6b688b6630fb0f2815b12586a33119c7c2e90223cfd140a734969904b4113e648922382f55931abeaea6f8c812495a84f6f4b05b1c1e1c13f6bd5796f3d4dd0896f34e66b215a7529595b61ad9a4e0a8c72e6a718444e9427ef184e9f963e3bbccb04bbcbf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habd40b3cc63cdafebe4ce60ada40f3894b0c92a11fee5d85c7e791553d050fe16b6f8cd7d08b4ff20a25f30c35359fe32e64d6b28209d871f3d3167e3fe439cd769fd2356cbd4f49e3c284d5f40b6eaa3409fcb950ccdf5663f96d22202d8fc014653f4262dee1c67d8a06de45ee2c546;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbf54fc58b0c1d96b7b3605195cffb9175d05fa8e6d5ad48eca006f69db8d2d0fc0df14c7aaaaba92b9495de8cdf33ea1d5d577554f64296045321cec87cd053d1ab323fe4ef83af3063e4250bb411113859b42ca58853a88d69d69aee7bd355118613d500cb70f26791d93122c5263b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58374d538fe14b04a92a921cc92abcc8da23027b733e1b809210968fa96434fe0866b483d7557608ffa1e08d4c02a52970d4b6a0b4e811259d7b48ffc56ae292afc2a33b912833696c0604671772faa34864e04003b97ae73862448c7da3d8e7d15c9390d67bad7b4fe8d50512e9b1aba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdf5203cffef656af40b3766e42a214bd2e7111920539faf2e1fee6abd051cdfb97a199dcdce0c337504214cb13945a61f8088514c633c5a1b00ce37110acdd820b750de3deeb4a9986c7bb54dee81add261de1d7ecd7f3b1f929ce5452e0b04b1e2955e1a087190c9a8a587b827d16c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h515a55d6e79faf3d52eb16b901d3e206aa16d260f47e98b5dabc32fd181dc88746d933e1e40ccf5c7d6f8a3307af73af37f234e2e5dfe80cc6022ef0105e6540f552035864347a345204bc6db11767044d3860103c83042068878bc333d5defa9a661f46f2f3c386ceb309fe5175f87e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b3539ccae188b583ed0fc0259887abab133f1a25c384187dcc4e04e9e80a9d0e9fc0958139d65b2cfbc135aec6af03ced21bc8bf4434e7f79ffb641ac16565c6259e02ccdd6dc07e75ae8154fdaadcf67edc74bf39483e0559621edade0998f550ede1c758be3c079f3d9eae596f5c7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f673370a9ef3268f7e263fc552e77892f12b89614d06918a5cb4aad47beb6e5cb8258a489a8fc7cbc960b246f8ba2c86e184ffcb8ecf7b8cc999ad1f5308778ede783a2cada1da987071b28e79ed4cb9157bf19b37275282bdf0990156d0ec4473ce3eb9294e5dd4fe0cfa2fcf6fa461;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd65a6f39c0eda1a2ed7323c1fbcafe8a3d48b83a761dc599e4256120f1cba6c72ddbba3125dc85b96ebe2ac095fdf0d3bb37df4a7694b7a9ce2658dddd2bc87456d9dbaed47d515662c3c8238632c2ca83d945015d2eccd2e8920be0254096a3da8d845e4728e9c0f27c1d8df16a4ae22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe861413844df1127fa2d7ff93df4f948ead420356131b8cfba99519574878b7bb302ba98b11fbe4919c78322f7e0ec4cb4d3926be55fb76ea0ba99cdeecf3dc5eac690520f436007d2354312149c04064e8ad45951dfabb2341a95eaed400cc5beff12cac68d1784194a7671dd3b9526;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf430cd77c718200552c8f5527202434b1466c25af84dee0a41ac554fa1dc2234c22da3962ceb6ee1d0854934d8779151e3473056912ae9f1ad9d89d56f53ad6000198753caf747315f2f7c1b53fc017c15d4e3af7674e4e4eceb1a57d4bcbd2cc40350dc4283a89aaaa0d9f934b12c9cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdcb7e6cedfb2709856081bf2858bb5f5b79c35821bd443ac70a0b339c8cc1f3460ac16bbfe06583f670e2aa11f2105b66bbce7edec043eeca7805984e2b0a33c935564e365bf96ee3f6c6ee29186b7b9dc8b1f6404242ddfaeb21c1e0397f78a76b0c06da59cc709423e8dde5613ae55;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6ca848ad746c24d29e791af7afedd5ac79800a4d675e17bc57b269c43a7c09933184e219b57bbf85ee577d225247372921ffbec21e04a8d05aa28011839cbdfb1fec0944e3fa5a446ce822b8f019306255bd00ed9b76a9a9adcd4bbd8de208716e0e68896f7eeff0f96e3d70f177affb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e417e87e3ea1b3d5b768250649099d9d49f6688d763f623e58d340818c158402b03a5643ec85cd1f4504f3ba007bf9fc8695827738eac7bfb9d6e9e8eb10844eded034536be5fc7522e3fbd3cf493de3fee9093618c1effc797961365fef869a342e293b37b7ad3ac4f94a0ed741fd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c5958306c05d511bb7db6ccf27b50e08c8d54297291505245cb64d8daa36c5006998846f9ed792b51860e1328f62100c143646d91b62f42fd6fa6223a87405427224628ccf6ca7a837445b6b11e4048887ceb546708ffd5fc2260dc0c54479b104b906d996e69137a17666fbd37cd2da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h253d155200b8ddd31fa2921c0d7b3b2a3f2d6cc50a27d365d0a4948795fff52d2ffc725225335a77765ee91867321151cdc75a9f057b8d2675b8b3fd1df534882aa22353a8f3463f4cf6666215de5bd252934149517358ae35ee55470e369307f4ae3442f07e7e3c44f2632942801bb4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28dea2938261c36e12e0ad77936fb0a837eb3f17d83ce674adc61d9030bfffe2fde04f9364b81d6c2831913508bd259a95c8073670d463f9db1e3bf2c2df9a1f88fdb75a9d0ef8f391cabadcfcf96749cd0ca99eb9991894b95feb9eb565058427718748b8d9d59cb53549c6a07db4c40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h902b21b09acd29a1774d11172459cb53cc982eb07dcf577544265be9ede8f9c34f94c4f3ea5a43a3ede72860b9c230b004f6d50834f819aa8fb482bfeda9db249f998d92d8abf0c02880b3a7fc1e90d49462ad68e238537982f1917d9e1bc4c9ff99626b729ec6279a34adcc68f410f09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7501e06b659237a03b5f50a92eceb8d6c55b6b3df7eb14717cf2c2cf8a9897e94e1fe6f4f675b64910a4f5b4113e70769b79e6742d01cd9e85c1e835b90a1b19181a78cdc4545aa8d708037e2a773ddd08333d3bc44b8f4d1b0c32c9d675636116f34ce764b2a938e866459569e59d835;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa07796ae3534867464e4e5107d2e29726de8965937fc740aa3c8ec4d1eca65a113af0dcfc51ec00089bdd24c12c46fe0317db4423c6d196c310e4cc05e398526f0c7e3bcabac6819034cb9b83b083e43123f7a7515e7ac892c700ebc50f175af281ba2438e8c27d065f50c1cae3bc8db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4f9c2441ec0cb593e155d5e6ddca2904e6bcf3bd9f80918c55c66c52e9401c90e3de3454a0950a9ff9e8b6981d00f1b4697ede25f348e64de9c080086237643e83f9a3fa4c0609519070d1b283af379df4cbdca1a1b9009fb5baa7e1852afc2dd28dcb3ceb8d2deb7d1f43b563339fef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h297b4c2452046c521781fd1a73c54c2236bd7b3aff014af0c8fd86f209bcb855f8c62ac014882ec3bd96fe9555d4b7460c0630daba739e322a4bbfba697db8b2b2b8644817360af7e8f6356f807841aa77092de0d14920ad9c89383cc771e18c837f5ab28a52f2b19ae36fdb311a32065;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9518f3fd116a1e4e06fcdf64248e9c1893174183fb983802cb2282d16c0f4d06270e99e7f1504193d1ce40b7b2fd624ff50674dd322afcd51c1d648b64640b6a50985342f861a402cbf15d46a06e81b137191270230f6dd047d32d5c3a634396e565ec571cf9e9c59a0c4add208f93234;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cd2ae4449f204b0568993dae42fb8a1374e04c50703e9fa53a5351046fa4a3976385ee6256c461b01729bfbebddf2181ef9f647e77cc1880fa3b1f3c85588670ed00f7dba3cc666d7c68d868358234b6a965065c44307ea396289cc7ae7f1e0ac0895cb8e40b6295ede3f8841a21ad2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60dba7ddfdc933c48cc73b6119dd19a11be4ce4f4f978971e6fcd7f70271bc3d5f0a92a1e8927107ed10a0f17d86a03a28cc2e7314444c980327d06506fcdfb12061cbbd7aac7dd76dc4ef22e6a8e56c436d59bbaca2d52d21dae8af4a713621fec41248228829061a426fc24d75fbc0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c13a4a7eb78dabcd6bb8df61f15237827b342cca533a7ef647acf31b190f9b7bd555ffa37079ce206f1de3e6f38737c11d75e0f362596d3d094a1966e11c2d16914c2041f7e1914a222d4f225983bb9dfde9a186bd5d80efcbd2ef61f674bf148229d97cddd5664f159f65d1991e7d49;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c414eb015a086e8cf87a556de57768dda8297cad37621cabbe1166b3f8edaff919fb53f9cced9d0eac60e284edb487b7037f88c1e0f0aede0a31d6fed78315a6226889f503b1f09699a7c79510644890886cb67a64396da0b0e00c89e0971bcf5c1d7eb05f100c44da7134343477d97c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47a15067b916f36b08bdde979a5038a5ad7ca30b4ae806958925bf46ab269d14ec1a1d315a3b87c998e116fd124659f7eedb2f9be88dd5fa1b1604d2b8f3071833ec0c693dbc6014fbeaaa4d509f773a82688eff23e80357419e0b173fad6f70de1d393f5d62db82e17bbb4d530dcf211;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d0c923bf6f992a25e1e713c2dde98e424f5b95d21224f7d3a2fb328d63c152889e1459ee98f5a2343152750f98f7516418e1fd9fae8287591abdb641b0b9f3b6d58b36a2e204d7f5133aee277acbbc5cd079a340bdc89850d147ac5a9d75f5d8311d986263116049626fcaef5c512da6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e951f8ceadbeaf0bbfc567b3db082bbf587d59df3e4f675564b1810bdc920d67d62b1331b1e498d2135a1fe4fd37021c44f5625d741d8338bd18de6bb5bdfd3eacb996d4c366c51b791f1d0bd8e00f8117e8a4239239e3e8d0314a95b7de925d0725cb6e940d8732a23ec192be469137;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedc1588d736c1babd14492a56fd76b996bea07cd26234c4635097c9a55d3d41c9c8ae611ad1d71ac5b6d62cad55917a8b6165317c0a56861d092e1e55c6ea4740357e3bce5d8865809429a9584ab6fde011de5a260a5045d476cdfe8340a8a145cd15713b894a374d9f134683a178ac5f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3426e7bd1c55742b9cfabf42f98d41dd9b33c73b9e71f3c4df2f2ea8eda30935719d42ff03006a4fbdd27bd191ff08388c49317a03b7a9ddf07ceb70c4f6443d9e216e18394f19ed37c26b32c4f835183aafa05ebd0e181c2b38012539d1a528a37fefdee5dfd12951caf3f4b12740e2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d636e38b9ab8c416b7c9501e9a5441a05ca47b48c59f2d1aea99e14b397736e0ac693c505cae5ca13f5462e933fd40f792f7816c590a6896949cdc570169ce65c69fca01c10f5f62940ee8dc17d0243b23673e8f18f94f9d643ea1f08d5892755bab5e5b3da49067a07ab3c52ddf4316;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h108a26bd2f5d3643bf9f34000b04b7dc4a81c138d179902eb5c7cef33c458abbda4845c7d1022252a83495c2a49a0bff4ee4410da7d0f999bc2fbcf07d77b250aa74f0a93b36f2936f493304d3e67ec380a4b9ab92161e26ad3fda18129b8fa37200606837cb6904c99630f38866297f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d6f2a96923f4f1a92cf4c3984f18af30673a3d66c12ce9ad4d89b79121024a028ef0e19cb1034c9e454e47a9d901869e3aa1c494ec5357c1fd34d58ae48794eafb34268705208d1834ca903a39465a79500f71f587afeead8dd6a944226374a855e035cf811f6505af604983b20f1856;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h106ff4e2c429591de2cc3d5f61bd2832247759c3d7d5eedd02268a03837770a9d41cdf209972da330c2203c3ad738b9c8e69a95bdce25caf11f4e06c8815919087a8c83f169eff6e2ae4ba9862ff5312d24b508d95d5cbd8474736f346a7613aabd8ea256f48bd63da4de063dda190048;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c0f55b3efa2e26833507ccdc4cd6f9a76c4a13533e93b4d0583eeb244ff63c9a69a36f59c92eca1e1680f7d91141bff9be5ac3785b85e00e08ddc31997e3f263bce464bc834bd418e87535c0211bb4874e8047f3604e7c3ac9457192e7d94814bc3f8877e49bdfbb9e1f51173f94b24e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c8167e3134a6b3c115d84386bf388671edf5a7a77e8f666c8a38f05a7ebe7035186f391baacfc5f5dce2d5f5e70bb4113c97d0a6aafa639781ce51b684d5b99c920f43883cc1077cd0c617cb4aaf00981ae7fa38b90a953364d94b0ebce92fe139b1dc1ba7e7658284bfd3c4e70636e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eac82e9d675acc9fc7e3e198eb229fe06d8fef0af3d6972defb0aee776a1deace8bca90f3441ee2a1e7150eece0f67affaabd193f1f18e2c23e1dae979a88af9f1e03d4880ec7088fc91650b2e1bb7cca5f464df4d6ec916bba6f8b576cdb582cae9ba3731d782ac40d1cc43abfd1947;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbbad0d5f2201e03db9fa90397368e1529e4efda2dbf75f6add9bc46deb29a292f51171c37f51ae0843b8ce3bfadafbd4d9779849525e249d3743a72bd1f8998b5b40363ceee993d49d795c13ff5dbee16dc8b5a157ca86233582fa39a2a80074fc270a3f2b1a842387f9383e36350718;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc80c3cb3106d52a869c8288a83882c5d46fab7ee6cbd76aecca004eb51f8b58e75855bc881a1b12bdd0e0b9e7ba646ef03d41dfcc2a8c068cabd26776199346a760b9a41bec0c3d520fc0e22da301e0ed016453404e12de07f55c694b465c83fed507431eb74f57e231564c8bc384ce76;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d5db79648ab2a554e6db47bc798627b818845e158a483e3a64c1763da4bdd5eca581ee9aa757571381d160617195e6a0d2064ad5f500a1da61bf07176b30e7ce64a75cdba18a2efcb820f7bd4a55741b39b3bbe86c3b0895c53f803fca8616ae96e5d5ce5c1776a091f550e091fac255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc5e0da88dd83be786c75c89ce00ee62e4cb5b632be383d47dba42d811044729885e7ec805435155a0d0114271cc8fd76737ecbf12e38faee09349b36799d8cd811790b406d1b40de746adcb44f62c3604efbd78742c3f4532977770f0868c7a8003e3b999d972bde136b347f465bf333;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7eeaac8641ff21caa99a7d6c1681eb4e1c83471db3c3b6002f874610332de148d8f59188ecffd7761cba407361f150ebbdd63fe79bc446b0d77972889ddec42c75a836904a45041a29ab2904ad34feb1569a9e0681189aa4e3b89f906b23dc7536197f742bab011baa1e680d645bccead;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38bfeef10738766b2f5bdbf5c0446cc8d779c9cf31af78165ef9d2148c544674057869c6392c4d898cb264d11dae9757fa0b8bb9b8fdcea1a2ce32546e80add5ec6a3f9d46a11d8a78ea3715d57825612f2c3cf0dc571ec96fb10a98b1a2be93b2eb486c5b3d1047350f67fbae5343eb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h969ae7034ba43affdf01086ae3e9ea02d955c8c10e7ee6ff5a9b510d98d304d8171c3858666dd1b79fd01a82e228543ea89c2512bd9eb4513485e595b3258af8a4634827ca53b5cb0d6349e7cd2804061b2d17c7c065eedfdf92e3e3c2425e8485b8fafd04dd58c283e5b8ec77e8cdc1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ce7e90211b6d8a543fd3a4cd2d63843bd7042cf311e2b907a46ead484c86b0ea8da99ea3de1bf77626dd8fddcf3f66d401c3b7d4c397d6b37edc695cea3db3123a1b3a6ab735eb28a17b710b4e0f17727eff20dbc1070e738af2956331d6a0561bae6546b042d0ae59a467f653b49275;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h391e48bc12856e249ebfb4eb389ef1d31e367290b1cd73c63692d908cb13959cfac7aadcb36a41dabd0fdde2d21bbe4150cb584581c6cca8c02a83d266575a7a0c505565dba53e66566c2a154fd48e00fa55c7b402f86d41ca016509e1750dcefcc35ea22e285c70a695419474b32c0b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h185c3f4349ef33b01c233735b40331f5f1560d45e3073de9042c1bf45b289769be18e168244e1b3566ff3c9e427650bb8efccf626c4d449a1595ad53444939177749cded65e46dcdc42fad443249dbf014a058a680173e909175a4fbf630069a6b0e7aa09c3afb801cf3dd52924e404b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28b810d55e73f7dec909973f28ce91064d56ca25e2a3a420605eea49741c1cfa4bc27687691a63f2d5e7ce0f4418d3fe50a2eb75f67091cda78d5ec46edef6e031b5d04277771ef86631fd8156bdf88cb71fbae7a5470651a742aa320e7663140cc35ae0fc8a122a2cd474987c92d4772;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb725910194617bfc1ce4cf9027d130e522fdcf1a204d814c157f816ccbe949e7a0934d3862e3b391ab521f1aade2d9991835e055dc2658a08c73c7a5a49b0f03a0a3f4d8df186fe790236d3ce3b08daa603fe3b934fc22c923d932d1d8b1af093a11059dcde46d854a75817a04ec89d81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfa061b648564864680c0d2d639c5d31e7dcada0ad545a36c87838d93965c193812fa30aec0868dd48e85bd9ffc7089037b283d014dd0fa162071e257588efe784046a81458acd16436c7f4631a2b4d1c23fd8848fe544cd4b261219e8fae9b9ba7e04ff3443f026dff7429d646b0fa9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc781d844523fc5c211596b38c4c2563ff3901215ccbe33e3d1f58637dba59e4f267a9097d3ea005172049da1e6f8b41d99bbf4b2b70b0a87a0ecd6b34fd22dedc163ec15dc74fe2fe8bbaaa8b7d7c02dc16df528cca57eab3b1804bfeb120eb59e878bc30ae83f034c288b486a7dc3f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he830d31fe4a4c55fe223b53abe85be0b2ee247614b9277e93ed218ef2b745244170d92f6b7406e48b55f8617893e15a714a3db887c693614b9bb42f757b64e95da31dbeb72e7ccb9e879413b87e971dfc605eb2a1d5b087c68f4522e48eb6874d52c0366b261229b7bc708a7f950fd604;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54dcbd0b534b68aef188abca36788ad23dc5077678afab0094beb7a0c5a9e9ae6a730e3bcd75a641be1be550e2b898f463a3bc25ecc6d50d54927ff69a7699d208ab4b37c369563b5ae0866495493c8609883110eea68f0caa898329be801f59819a58e1d85a6ead3875fe4a35e044d03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb72e5815b3fa95048b852e0548f863a56217eb72bcee07fe1c9648f55ae7b53be23d64b7f39cead209ee79a708b5bde7e9dad758ee3dccb150d3ccbc55d5014c5bdf0b415dbb9a1868cd6288d1295dda134e1fca45abec0bbe72dbfcc3aec5159cafe8f252e52dfac562b873119872b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdccc84a57a9cf2d7297e4ae7d0e7e09fa0234c9a5864a0757fd2a94c983418684dd3c3c9d936084adaecb707c2520bb98da07322fca173d4470bdc1105d58eddf61f2f6c5c1ef9218c3173978237d61b55d773f0127c3eed9760178f357af5e977c8c249128da10ccb5c18f26f2ba4f51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6cede3d139ca20a41082e12a70949b536c53807f707271d610b6f87d317f6131c7ef174fae126826fe1eb6d6b2ba5df3b81286fe7637c7d0f64abf9ab79b6c4d2423644fab3829c0233061c21a2454eff69681c5f7d134cbcb840f2f3d7d4dbf70e482389a0e3542f283c86e53b83df6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb164542ad42f8f60749568850a8bf02c238611fd2502eac63778e19bae0efd6ddedce31e0d865bd0731c0129a5f40603dded1e4eef4c5ce9bbede4d8ea5ab6a1013166fc3ec8cc85ff399c61bc7e8d1ea7ac6bbb25ae52f0b4559fba1671829eadaf21ea1d36a12fc48417541e32c3cdd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78affa9c8260b06375b12f8b6e966a19e80e395e8f35eb56d39afffd17bd470c698c2e1560ae6798601520d952117149634dbadc0386fa3c4211e3d472d932892b3d2b84502bba7971226e7c0bfcdef56c4303de0bf559b7e37ace1938f0d75df22cc863f045cd38373b31d800d04ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85405b5ebaa47e68679db243c73c6dff99f92f7a045ef558900e7c745a92f305e4a3c7a5f186bd345de575db2f7ac7089cc4f9bf556c27aceea9ebb2da4494c1b91c873eec7b7fa3b0f6db85e925bfba2915dd60a186fa84cb4012327fd5c24df1c18e3d8053864b9957c6ac12e3e4fd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4c91e95286b62546264605432bca49c93e4eabbba206618021bc6d80626b370192624f376b1dd65384dfef02de24ee5bd0fc1106e3265caad22ef8b4ca8fabcec277541b69e1a82aee8105011588fa78713ddd477039ef588783dfb3d95bf48eb0d7a526ed1448b7820a1ff4ae0eb331;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6571a16a2e21d8957c36e1224d4695c419155d662399f257f4f4b81afcccaf59b88928f641e9795b657d513cabd1e8cc46456d0451ec2d6d0d120d667ed37877b5ad48230f4a4612bca1aef99f186a7f0259336d3c3e6456f7843f539bbfae30f2ee3abb79ccbdd822d780f755a46f68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ecc14a733ee4b2aed7f6ac138e492f6425d2b60e616cbab4221d99d374a1ba8bf5b3ba286b3cac90c09553718948de1916e701e278f3a9c6c2cf105de237c71138d2855637b8e1b50a9586f7af7a3faf8687c8c3df23dbdfd5e53a97bc62d5855ee08c7dd204b31cf971ff07aeb8d74c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he455e911ad29a054d21d4ce272a02d510bc675bceccc2ad5e4841868dfa448523c45e97d6b4dc563bfc688b77cc7b6e3f7d33d5130769afb718ac68268ec2cdefbe005173fac32ea70f980e0c5650e4d0815c469b16b6ef5572834b940a0af82c9c3d1d138cee0e27f2895f07c7f88bb5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4144d7e0dce958e94770d052beb0432a6fecba54dac57bba00bf369af180ac5771a1508998a826d19842ef9710089eebaa664eeb5a0b7cc2dc792cb0487205bd00d01899345e77c1453a33b435e53dc15c2532d2d4ab39cf001fa3af24ac8e8fbbaf3c504d6d525b2905e5e5c3234e100;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha13add59f35969f9cfa72ac5741f517254053b2f9b30d92a8bdf20aeef9e975800ddf65d6e9f6613104ae3f35c89e53d85ee61dcb707013abf10758350f1f2a5cd38aa0346121f35ebc299e2382ed797e5c0cf6ffef41f0dfd4098913e7880999416ff49940e44d42b0ad9e08e51f283a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95469f7d0fbfcabf03a5c2d4955c5eb8209cd483b0ca9f41fc04fa089f9111a7573afa9a63285c740d532b2e728ab6917542cddc3fc3ecd8d833c31cce658a8876dcd9590c67e3850b31862cc0263cee3da38f8daa537774a97d7c8ffad8ab134c42a0f845bf62a7c8275f64890cc4cb6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf69222a9853224bb95589b062e013ff37c46c6844d2b39f40210b8ea773197ee4edce7f5c5c3476e7f58303244034dc748bfc4a89cdb6232ebae50b42274a3c203383f34ffac929b80ea0e79f44aedd4b5a025d78af21a888e1ce7b59ab0b47c3d0b5cb7356882a26b739711531838fd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bd9858a54cba3ec8f3bfe10bc3ed735ac97bd6e700406b6b143ce407bba2dd255d9c7906b14f06e7ac1b6f68d6ad64773c72618881862480a0ab07d1fb65cd36ea3725068799d43619c058b18a70fbaf1d2c2fbc07124aee5aa2e9905c7de224f2f745b6939ec4ab23385cf850806550;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8937554527ad1abda577f609fd3c2658af2a9d44b040e4aae8fe30db0822d04753dbd686ffd553cdab880049c3b5c3c24d81debdc2550828d4de58d32cbfea4a3ca6f0b050055101c3c0664a468d171c56cc391d39505166009bb6c16fede3589e21911c42e3fcc3be3318cf01f49d6aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9cd13c6f88955119bf2361b060d912e7e0cc794b1953c3bcc1f28dc4fd7f714c09298db4bc2e4e11fd74362c75c9b59838f5706869b0b70924e193b4fd81a1137d38eaa0e61e7bb3fe7d68055dddab90d6aaba817e37fbec36707183fb9b454fc6013dc1a06d666a5b9a89ecdabac407;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a064970cb37d83515dd0ca9b9b35436ee4a7b37a87296ea12f285653a3d34c4d0c3e3103d142b82702ee1e8c9dd47ebfd42ca1fbd90e69375fb5e40d322a0d81d5c6152e5e33565e63f65b727296a3c5878d1668799aa1d1fa627d9dc263d605a29a083e1c95a8a71fdbf902c39716a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65a5fbb45cdec0578314d14724379687ef02ec03e28785b4266a8af16aef9b379742299d4c7297bbb592619a943597a6f494b12846e8412784fde423192ce8ccfd3108e6db167cb39593d3a6dd5867a3ed6b7453b846a30a0a9bfefac87d3e5f88a67d10428d2d30dea3fe5be415d7670;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e5f555ac90cf70a39d3b6605913c0ccb3fc23a754bfcb671924247d854ba1aba70f8ee7f8a43670e493b01ef2fcb7a16b4f6b78f39f19cc279130bdaf6dc0134ac7a99411fb79e181b91e6dc5df102addc00edb30d979dbc3bcd9fca0dbf28e2e85445b8acf5bb05b963d250e0123ac7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b1604481cd1679244cd4b01000f240c508c2d971b12f4dc20019938621a3d27d06ad50cfe8e40292e8099a56c9f5b52a2de1a55e80d5b1e484f1e47cddf91b06117f28445abab536a229723e4d339523f56f8d1a545f58413f7a863f5cd9282d94404f7fd813b8c4a9d299dae4bba214;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8648b8f0b12f218afc3473734beae9e9a130136235edd5e067c76c7a9007574baf93692148dcc43889c9fed8b9910bdb5add8baff8a23241c06b3a9a3afe150eb55c16329e28017f687f0b585034dcd69a0bbebd03cffa018d1073eaab02fb33ed54919b0051dab7403823ba43d1d439;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d6b1a6642b18af1de2752882ef8974d8f9380b30631a48b6fb70d0689c116e2ba243aa78fc29328b5f0f847e530325484740ad8f94af814040a4f7cfbc57d8fa0a2ddaeae9f78edf1555317fb874af643df7b7520fb8ad673d50218729a7710c8eeed231b7c1f8920828c0fca22b1296;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74d89cfb86d45c7819e0b95eafa02e4ade852018113b09605e99d2a940df343cfb5da8f3635c801b61be5bc902fa41cb5c0cef10b76bce8cd169a2d08b79e8387af82ffcf1465d99f61f1196b5db9e0d5ff36951f66a2ba1ea288f030434a633498635c22c3823f84a9353f1fcecbae9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb48446d53702779178c81bc554375cdef4e6f45229e1d39fa5ab931ffbdb632be14c381e007fa44b99a7c2b291c7c2c132703b831beb6c2e7d3563f076b84de3193f33f3360e75cff0b6b6e59f090d2205cb8e0f72e2378429c5cdb916d1b2587433d4d6ee771f9cef38a5b517ef05b3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd7a33fbf4de910911d72bb3d0138a34776d94734cdbafbbaa474d4bd3daf7d70544f12de9bc39c7e469b27b44eb9e7812398686cc40d4199d888899550e1695fd5bf1bb06d74cac79232c58233af30ffceb6b7f1178e274219d28759c3106f140c527d03f8005f081efaf38dde434c2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95625fb0ff130486a465013c750b9e1618e4bef15bdb629550c0bdf6823270a8b99894b5854847c454e0cc92a368902ede3723b42e5d91cbd60441fc63375bb566e3f514309890888d2f3040c01d521a0e40fbe86c1723bbd24680749d2bb2a99f8bb9be615df26fffc2bcd5fb611ba29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacdf9e858720442847c7ff1efb011be5c001f9fd0ed726409f060d4d5d46bca52d6663774278ecd43b9b60cada1530b10b02a8ee191a6ee6cd7cb05677b2e7033386e24c4d0608fb868c49a7dff5dd130f806aaf38c0cd7661a0895aa5d2aff871f3931e4fd082fb00dfd45e9bce2a1db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d8fe197b07edc2a2b9a3493d328dd574e126d2f7103c8e53e727adc53ea5cfe36bbe8c4724c07ddea4add4c8b9361da5ba1cb5a12add53544984dedf25bc3e5219d6f9133f08f4a68051f1e0675df022574476d9d567810800bee16b093eb8ed828a23db980ae1169ed6402049f4090;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca0824cd70e448d8bb62d587a20013a80a2d318cdb01940199f1598a88700c84b33a4f614b3b5a93486d01fadb66506d1c20311e3b350047ab492496e8f2c67a4375ae96b28f2ed3ccfe56bab965a035ea16d13321df71aa17413657652e127c3ace15fab92f63315db2777632bfccd25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3d80ed04420a76633a8b4874e207be6dafe163567358332096367fd70b9f4d9ed9450f3aebf64a364e00f1a355ad53adb4baeaf7d9f963edd729db304cc3693e3c69ed6a7a0d8b54cc26a2a7ce55c41c46f563df4b91c8cebca3c60bb92d3411bb7bc379b8ea2a9b70e0b03c451ce6a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c02d72544d4f125bfa8b56731b71478511abe36765e9706bfe09cbf496e3a5dfef2917af53d7e68c533f8d38a4bee18ea27a1974236b9198536347af0a6d421512dd67ab38551f48a858ad29452822da79436b65da7aabf0086b006e1cc66012b01560242595d579cb3f6ffa34076522;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ebacb0a500188e9bdb1efd47af4a3cb670284ee3b3756794a1434e2a70dd9aed123e2abfcc7e2d62c6ed841aae8663acba38f7525f80b9498b2e5623261495b4e9ae9f6b8dc1073f61f505917b45f45064832e88a174780df318b90cf3b92ddce09ed9a07350e62db8b3f2021221c86a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf76885619d8cff4f9e2aa7e31b747a6f1e8396e0e05b7f968bf8a5c0d53d6729df7965ac90bc58b83a3e90d7c34c8f182d21e5a29f2b38ce7913334a448ed32ceda460df69e1e573beab934c867d07ccbeeca531f6eaa3433f735241f4695d06b74dcecff2dc8bff10166844f5380afe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he179d0fa09336360eb1ee08e32ee9af6f9702d84b952efdf684150a2bf9ceee86da5fbcf3978e1570eae17a65ca3edd5f95cad49f974d2224ca02185da5caae4cd13ebef55edfa2d40d4cd7f2f69b855202198568883b4e9249e58b4dd9af113c7c014a5551ed3e7ffb265851871ffddd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h704cb66a5e24bb799e5d45ff8311b452f883dfe0102b3c0fb76805788147ff55aea4bd06f8e726775dfcbc962220b88a5ab51eec3868441abd7b9bf9f8c8fb51beed76a449c8c862ab1920ad7cddabb0d12530b98c2b6d30c908f23de91695188223161022187f6bbb8e95440543c47d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf542edadd8dab01c5f021faba2d3b32593dacaaddf87dfb4abbf8c5ff7f6c07605870c6ac072f7ba05c653b05847cc35a7bc247fc40d2f0ae9fb1bfef3e48c7fe0b6258599b3ed95c9ffafdac1ee89950147b9caf97079e5caf129414ff61a27ef3557b91edc1a082d24ff0c55afe7f50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40b0a2417c0fcd8fcf91cb58f54dfd5983da4e9ca32c50c67c8046c06888816775f6fbd2450e4a4b7ea4ec493b8c1aabd74bb58d44cbb253a27f8534eae4d294d9ee53266b753cc7b78c7b922a2b1b7f9f4a26d909c652230dd6334e38390c0bc1a82cc6b41892772bec4c86004166f19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda7fc8557cf95fe271f73d8b8635b5d62d518aa6bd2aeb9b330efa828ff6bd2fc1a3678a70923805ad44547d4dcebd4235b10b0b4cff1341a5a5f22131a4c5c10cd02bd257d77c57bd3a089ce97eee0e8e92e23d046fc2568d6033b2dea97d169a50a3e2061a7e34c1809f0485d52591c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h409eae069bd90493429325c236baf93ac5d92f92871f751e12fb74eabd105f7c3ed9d7503cf18c9732e2896cc82ae0a3f02638deda2691b210f83faf666bf8f9d1d7ca8e29b8420b9d9b62f46dcf435138e099e6e76b7e496091238179fa8b1c53b256c70b755f1f5474d5350aeaa1fbd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4db707bd3b3755839229d230845414720a71695ebd8420b951ed1aa3cfef08f16c87c9b958c43d9da4e489654fa22b935b12c16f6cbd51d90c249102c4c2f6a49fd80b3dde351ae721fb26e5208c880d496cb8706cbff4c542ebf279b3ca956c02e41fa6f5f62278df3b96a1e0c635210;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46457d7d6ca9381d1dddf30216ef950a70302ade31012438db6a8424ceb8617df449925077422412b914530bd3b22f38f7df7159328ba76c93e0fb43f19e2f96c6c3df9124157b44e41a9d013fa077da14665eff88361907fdcc56f7758f267ed7adb202b8fedc5a0306a1b4cebeac01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbddf121ca03cc1eeafcf7497845b3d10b4db4f89241c3145959b10c7408a5ca7ac77c3d18f4b3f95058ae1563cd85a935aa7b0462deffd5445ab00291a055f83d9ae03f773482a7150710f25bd47c353072c37a5f1581fea4dcd5f91b6a14a9ed5ed64cfe649ea066b9fb36ee5abcd54b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe797ab5c189792b5c0615a3a1a3012407d152bf1e53d0c507fe1060b3ca9a4eabfe3c0da90c052d75ffee3678aa86ff025f885566386a573bfbcfc4764d859687391cd04605f61fbe46fc6eddf5904117a93e86901d656dc9aae62e7a594f4f5f29aeb6b40e31a626555130334c0d74f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h155f875897d6c56f593f026248aaf5cb0ab01162b2132ae930b8839f9aba0a674ad5b31ef5d73edf6a05c1825ce3ece5b40333fe9caa6017c213b320dfb85e108ccd9558c1abb2091a5ae46f30dea6ab30641744e4af4ee72cbc2dcdb331e743017f98b13f4aba31de0b5c8b9b0676a6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h423702c4400fdeb3c4cf02c1190fcd7464b03bb8ae7383aa7bf5a27b8a188ed43bd7227816e0fc6edc9657566dd4ae61698ad27ac877b507e37426949dddafaade1c4a2baba590ede4b22e6e36a627b2e24325cfe157a71b56a43ac7bc4c948e92042e4fca22f1b02365bfb88ddc0c2d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f4fcce7ed1490366522f979bd5f496984457b583bdfce12f8312836b1146bde3b0f89767104c40db1b25095a7c4bc9dc50fd640e28c5c8442f4fd90dbd1b714aeef252646793b2059684529b781afb7394b5367ed506233d2f83b0c303a84cd31db690225e9a4241a75d2e476e09b5cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56c402be03d91ed3839e2e7926119bdc1116d42083eae6dc07f4a1ced9614998a17bdf108c637f531369681181fde910718fd079715586f320705201fd61a0d38b06ef9ab3a53894994d5c847a6e1530f7ab7b5ab11848573a2a89d724c1efe52badbcff4365e0386eb81584de21a899a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98ad721695bb8a85b3cd50f056e27ada8fe48898b9c92f6261ea0c48955b88781036c3fc6acdc1692721863d8ca17e6d7c1c273adc9fc38a98f6bab3e088491359b6abcb8aee1cd8d39c95da5a7ac06639c540102e0e68ed5a993a8e4f3967514d1c2d71f0e8df320f6ff62403a06ae3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc70ff2cc18f59655db243a798aa8dd6234257efcc52f7466e3440258670f57697e35b9c76ed6cc8c8cd66ad8558764826b02b5a4a6a160f359eb5e67e03920555b69d3bea473eaa6adf1683594a1cb004a11a79a1cd469c50d259c6c6bbd83b4a0db5c24fa52231b77b4a8340594ef690;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c25dd1de765eb4192dd570447364ffb23944dc69c4e16ad6e22647820eaa7f47de4afd7f7f393aabfca3015e738c05233cbca895838f10775636db95bf5e8b5973c35c5f36ffcb3c6fcd165c23f0fcf4cb7dbb16eb71a5cd31d51887f8d2abd2be6f0f6793394af612df8707422fe490;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbf2b3c7205f8b3cd3490e5f6c60038ffe388f7d99ea9ebbff7ee1609d5908bd1b66dd242f766201dd47e02e8eb54976cc6a1c7250a23d2939df09574b2f7f0964c5295881d20556835b98befae954d0401ea90c3d7ed55e4d44cc00c9856632b52dc4edfb72407168a4372c3446a5066;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7151ed7160b7ab4243e17eaeef01e34972c98364d8c5286c038e82c583b9069671191ca6ff9d0f549ae835f40a28c35b1f7759503049a93dd18c269497e2e83b0e1c1bdfeb70d057bac5491bf80fc651effe1f402dcb538672b7dbab0e57b9d5d7914d0cf7fbe0a27b8a4f30c1b7fe764;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h979d3383631b54239c7996b9e764645c5804d07dc8c7bfd1caeaf32e83c689f77ef78a416cc72329b0d3c6f510138257f1bf9e0d9a073fd8334364c6dc56ed65711de856704fa107ae7bfa6624c064fd35e8a2445590571ff218c6e9d2aa0c0dd5b065982d74c9d07794ed848f3a9f255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc523bcecb396b3cf3441ab49081b537d5912495bab80ec404929ed3d6e90ff88d4cf03bc1b3330f56773b4e2243fde55d517890a4164ae530766de3f13d5fc64ef6d4cbe550c93ec70a487d83565cb0305fdddeec87aa581291ea7df64980690948d7ddb6739fb1e1d40e1a610d71106;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7eebde94439b4550871c4c2e615d18935a4fca37a874f240913c10368a7a4dce97950ba1f459bd9106762e92c110e809eca1615e269aaf6ad2793f16ca896e9c674dd7f7e76f64cb0f1e9a2b6b7ed8113ffde45751f2585cca2b215e301227dae0e82103d62491aba5f426a548e54af26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57e5d05803e18faa8d7f3ad60e26cc99f18a0053a0a710c4e3f20575d9e5c3918d5ce0f2a5144d1a2ca7dc42c0951b80b3d7d2141dcfd4d50ee9a27836dbd342569af668168aefc7b4d7f75e998492dd7723bc3fc5f50b56c9d14e0fbde54039ccffcbe1d4cba83d3a0ea87e927a13292;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h184b8cf01601415f7a3909a282e3bb39f0c3eb38eb4075618f7d7f0916043b5947c3051a4d057fbf7f446792cc710f103d6278e22bdd1a3ef32fdb2ca4f2a87263072b1339d3df4043ae240ea8f43314c463ab02dfa4cc6cec33d42c531bc12fe04ea5d74ed7fc968589d7a7308a97f2f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf03de07a0569c86f183dd4b66b16e816450fb3073416cf5dfe2831afd8966eee487cc2dc9d84248465e818e31e825aaa1cd8ba47acfa6be1383ae999a143f8af5c4e20fee3e4e33132588833a9215921c2b2ec6e7bd6c7067781bb706e599c3aa5c1064607fea35902a0d3cb06a063646;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68f25e350ffdc705d1ddc21d0e353ccfc51b952a41b88b622b819e8bb8598044ed386a1a5ab404393c0314743db5b328d903fea55c677085e36d71ca7382daad5ce01e70999ac1fac76087e73ae900389c51dbafe55257a3b0de660c6a4714e48e36bece48096eaf46b96579d0c6c3adb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10b7439cdba58c72496b0b10610f32c1ed5fa3255a2b24adc569b0f891a62dc06cd0644a57654943a0245702322e7f9209d5d6a41e7f8803b97a80e3a07494dc2dabb824802dd7eda9767f545cc311c7735f7dfc47c8b705972acd5448c14c3d0de2cc3918f4eb414f594765528bd5305;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2281b01ee5031d463ea9f0ffd05150791b31c232b24f86b758279b763aeea613e73697df9e2a4051691520f8679b386167fbecdda8f8fb74f038a805c65a31b3507153cc9c884456edcc96b44ca8251c9950c22086e48bbe19d3391ab0d49ca63a00c745443f770e9e3af64fa7cdf796e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e0e4d05e5812aaab75551e2e6b2aa61433d7202d300fbf20037fbbc520c0b37f1a399bc6bd529e46d0fb2ada4fdeae94ecda4efae46a0efed499acb53663775d4d7a6b8a562f6e9901551b6a3223da912471f949474bf31bd58687399766387976dbae8bf9e4c6e86957e0ba63fef1bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3be297e1367050a59aeb83c2d313a919858d065586b98702134535470b83703865b2ac04d81b2a911725fe05a1b6c8a092ef780d60a369d61ab4ff9258cccc2f16d5bad5dbfa411c6a4957bfe4ceff3eb8132dc405bb24f4104ba9af983df94f53c3ef5d313810a642f262500cfb8eac4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4c6451dd84ae7de6e248aadf57ca98f3f5cadeb67d4b35db1dbc4b9fdd2138ab5c5b567d7b8959951202be4d2d712c48ef7b9358b82860715b3beba69a704cd30c4515de10d665d114e2502f958411436c7787b51c4081222d44fe1ffe13f6bdc279feff4e5e276ccccd2bbd745294f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc756b650ded40bf0b54203876763565b7bdbd5174d35f4f5e843afff17e67acf1a710c2a347d0ed68b9fcab8b0a7b11c5cc758adc20b1359f16d627d50337f766f130d8191244ce5a59ad26ddd2d695f25ca1b2c840d09bf866d5d20d81b63faacb8224768214fcce94d136a613738d77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2605dafdb8295d2f57648d547c03576efac40bdb2aa025b40c371955aef3fad09573cdc1abdbfda851f7a226b2f63be5a761bc0ca44fa0f8ebb3cd03992fb6499d2c045f9845b2ce9aca7eb93d00a148fdd32b8163925069f8d85da5ffb4745e123a68d3944b250e7642f6cec9ae51550;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4587358631668b82a473a4ccb8b4c49f3081864491a09b587479c15a48cde34710c83aa4da59bffea4bb8d5f77ca76e6e0abb154e8594047e9a8f2d5cc09efd739a358047a549cbc4f903951763591e6c1ddaa538abb46bc4f3fc7477df865271df3da8d0850113c9a0c3259874d476a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8039e0dbcdba2fa1b5c72cd600a95c1d1a4bbaf0a94705661b7edd46bd7d7f9301c2ba8105feb06cd68f0e08779545710a6d24ac4609d28f9e29b369dffdae568c4ce3a8b46ec483a56fcdd435abe2a8835d11ae88940bbc38727cf4459a30f3f74893bf93cc16e4faad67e6a87acd770;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ad706284651b5552732678b0e8f1043212d4c93cb0820e6c8c0929f9712e1b188f666a2df0c2e9a4c36e86d3c57669104f7ccbb482c2bf218cba39c5a717301b6c026dd2cecece981dc224ac456fffaaaf8bd0c9ef424d2d1237cbb986e89c9451c84abaa61bc3b619c4261955196d94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3892be3f5ef36c1bedc9a75ebb72e5ed548f67063dba3212aedfdcdb9080fbbf7ba596c585ae5285c2c6879040136c7844a9f1c01b5fd7ea37e0d194e738fab03986ad4f8ac92d37b28266d95e54e2222a4618deed0b1748719ded2bc800982d07324c12198c2c4b21741b51ee5c77f14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93d2e403cd5f5006c14b3d637c216b246dcfbcc3a1acd36be34b59d0b7821fa04ce0c59a16e01ae475ea75602c7af6c1aa11d4b77c4b0279f1b85873095f6380d9c5cb2149f01dc90dd7ed1e49b2f24311001cc1d8235e506ba35a3790b04e68c7e2ddc53a676a301ae5e1d8cfbf2d67e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d3ec4790981ceaaa45732ee362e8ec258bdebbc2ff2601f675f8e8f5b242b37b21569e2700313a17dc258017c7c5b39951cdce199c8e0363a7e998f98155e30129eca7087e6f9f2285c031ba37826804bca3e03ebcbb62994a4652a2c54e36a4a0a500f12be4c4a900324d10b6f266e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54c950390df5dea68f1bafbe43b9571bd123183c1e02bb9e808efe4963bfe3ca24157f0571f69bed8135b695168f3441e874480b4701d8244f3fbc1edcf1b023b858fd8da25ffebdbfb7037eeecd48e44caeac368ca3e1f8401c680880b6553b11a24290c0e9cb4d0a1f567b8f2235272;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1acb1bf22f860de2b8172df765de8357311f91d181eb9bc80746e72d50f4d10483eaf2fc9f1c956d14d0f71903720060081dc0ee7e3393513bc2d051c3ab56efb3cd774a9671c6bbe958ef0f0aca00bf2f3ec4ed2106222063b324e91a86fcdf8151723c7395db06278fd767b548e1f61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha76eefdea194ee6e90c1dc57c4dbd9f6da14e959030d940b5a6b633a7588de52359a398e2cafd316e892c8f25eed72af13b04b91229057260754ed67a6d0727ec4b2552c5d2fd8974c8924fbdce1d8bffdc3432885ae344e941a3e022784ce15ba284d1f112ddf0902ec1368dae6b27df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fd5cbc4528bd252cd42cc17dcb514faee2006f6d15865433080fcdef1536d3ae3b02fe1e5c77d6edaa8c9ce8a87ed536f2aabc3380a6272c0bb086977ab952a8fecfdf1de43c9dc7f520ff80f2434c7b0d298b2b6385bd3182eeda5638b7cf28111e8421417458cbeea7f1c224a9323;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33ebb86fc9f68f18c14885ebc188cd654726f0488fcca4172d23938a35df2547e87d9720bfa6e0e0b59c095a56d513bd6e4f68af85e4085677ab7660a7262c1d3d7f7fe4aedbbc60f8160e00565f35089f3a678d4e3b9b19403ef9a9c1cc55914661c91246fe2531711c4fa90c5d4c182;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea35642832da01c7c83d0227a0654cdf0fa8234895a65e9a2a0d67550a5860624059969b3dfbf53477701d60a7f92e8bc8c31362b4c9701fa02124d4e53b56d8ee39b14c3103bd0413c5e6b4a4873cb57975c4316770ab111ad3b4318edb0d45d2cb62dbd58102f781e6a782fe967c47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h316207b7f211bf5c16e3d48fd5d8efa5b01be1df67cb4e4a0f67275762b393e33b8ae2ea0af2ebb91ae7a6051fec3f54cdb8bd9c26cbd73c4a145aca367a995e867d1464280862126ac3aa0e87a3439a0e6313d845cb740bf613b2d80d7b28124fcc9d5d84a67a4c17b14b2d812309ec1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c14aa77ecd588cb848fb3c70009b0a01cbf235778497554ef189c8c0ff446e08b98f84df67d02b635fa4817164ebf46a9a1b924ef7cd0bd04b02a7eabc77940ad64b65caeaf30d3f42aedc425ea5a752f1a52c852d74aa03bce58a49108cff12eb682802749df3f991361caae9764c72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfca61ef0f2a05fd3ff98615357e8b9304a5ad1c12d30a27040fbe6d8f2f1815328f694b3453fd34008549408657c4759c672095306bede49042c5700b4249d5895e9967cc844caf83a557d04a33ccb6c1e29a704ce1348056851c7af4d4a09b1c4ff9085f2fe5444264f871ea5791deb5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76005dac0a1fc4d503ab0a316febf00ac933afba39747c437454f064b31caf5e9fd8954ef19538868d54f0bb6f80a8728900158cf5975c428a0419319e24d5314445dfbb53fbdc238746adadf90eec0729ca70bf20548119b7bf57862ba0c1a3860f2ef5912cb158010b2f13d325b3e59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb40e4baa021958758c921f59f6e5274eebda0ac18fb3357ab1151f7b84e0edab1952b1851cdcabe2386f40b5f11d651c1720cb859dd848bb7d3c3d9e1757b90297b4960edbc5ae7d1299d7cf348c24194343f13d089a0302207907c0eb9e1d045b90e07cc004c853b6c1720188077e537;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1557aa8786730e81f49f9caf6025c8e9cfd2c54b06322bcb1caead53d9e5f33e88ec6a1b66364d78e7067ebafd422547070a8e145a902710916a2127fd412e2e9d76962d5164d6344a77bb53b40c55188cc3bbac6eb7885ca1f102772b77e63c616e30c8eb7daa3156a29b7a9df79671b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9087eba7ac4e3e5b4457481997925f4d44e26a1616f5eab859440e67d49b2fdb10b686b11d5213c1f3b0b5ea3cf72405b9cb7894b10b9973c25a264a804bd34845d33e6e5adc1f1203f2095f5c9df210d8fc1d19c381668702a4696b9be5b255158f3df15d8f917a27e43d560fc61dc93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde89902b8c7d5e8413b385398f010b11938689bb8a1c909b580a7707f7f1c7063808abc107dd9ec4c4e87a04459569513c3115cfe6dbc04c01307334eb4a07346492c375655e24ef721754966cf00455f0c66af3d6f80984333cf9b9f705cfc32084dda17595660d90585be33de2368;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha350fd1546a4305ef7203e27f4be7acfd63aa9db3fe691ab5ba6c91d472bdf765f877395a0be4c29d61bf2a35c8e418ec03b5226faae576508a378f16b83991b182d217ebd2d6252943cd7feb8d8c74c34553cc59e6c04d10b10add76d3d8ad3b61047f6fb17191363242f75dff3d4a6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf16dc7ff04783e23796051a9086494bbbd26193c7697dcaea574402274336b3b4a0c18b153eec502ea051a11099756de325cc50b187d7b39397df2363139915e1f2a69cab52152161680efae4869a125744e70467622d40ee2d82e08a26c828645479e858b9846d91032245aa33457e0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f5930e532d415612501b01ff4cc151a8cc43224777cbb10732e8e219074cdadc6310db80977b1364779e7d0a480b014ba480494d1607975cf864d1f971c975a3ed81fc463ce266ba733953cd1b94832e4ff641cdbdb7fce4f53a10b34189fc77e784b9ea3dd17dec3f55c71f9a3fadef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7142dda697111119d78b56ce5049b1330e73c5b232ba01aa1534e277c9ebf572475f921fad81254fe44110f6d3363e7ade28cea3ff8fd819bf4bc374d4906f180932b74589fd4e6d26afd78488934abdfa5b2b16da23e1a94dba69982a9303fabb4a57cab3467161d8b6ef85388fb2b31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e8e66b380e1d784bf6da914e4eac4a627a41016bb64fc83fd3ba16aafe593447c6f77dc15231fb703748272b24dd3146e6b66599e2a27b9a91c79d5434b732a0928e478af93d44090d8cb3804292a362bc2e63440850f100d0fc958a4520c464f1705c8858521fd725e1ed1fcc8199df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9d328d254f3c251718f0fa64e3df5c948a191d980f59617782ad8c14310a62bb72844729925e568fdd5da579d9b304e64ed0b75306f1b51e545586b59d4b5f76a1ca389b04ca62ad145a6831e0e1285aebfba28a5c12adc3b42620e00266c1b15a9cef48a8ebb9564a5d8bae9d66b65d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f71e5471fda4de41f2e751066f929751a8641a5ca6fd8cf0bd1631404e6458390d836073a7e44beea5cf56b0f34615359df06b96f08c51258950dd3a15d311ce841bffdb88bcd58d50e28c7d9f287fd99e4cf816212eed1ae1fb8c616897ad429a48d149d54200c87a467ffbc7b25882;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29257cf9fc1ead0b280ede26d079444c8ba777720e73c137158838bc87ecf8dc1e82a606b25a6b50f0ee43985dc0f072978117d55f91e7b94733c292813c70ed5fafd9ea6688a28f305f082690e0c5c996393b87fee5bec97c86d2bce16cfb565c799091b1bb0e9f8591b74baeed6e1c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e162cd30f2237a927224f0a3eef2ba500a42a57417df82a64c372a611ade74f346336ce57c4eef5c60457f0fd884321f125a6de1a6507fe9a986888882a2b74e8ca24671117c5d76d73e4a21508e014265ac044d8f2ab76b83d68815103db45535806f45e72e9751b7f02fba38fecc72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2366b9f50b2eac5f12122007f351a5ce7dc5cbe1be0013a9260e27613d9bdb9b9db5ea2faa366c6570345fc270de311e7fff8bcbcfe4eae4b4ebc184b6330a9d5af2b5f7caa06368d4224c3deaf60aa267e553be372ee871188f4d233c030be4bb3c6e02dbf135551a3c14dd6c6271753;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c9b302c115c5aec92de03a445f623fe899d92718ffb875a5c9bfd9a63856945cfc9253dc85d37f475efc85a4925759f328e1e645d9f99ef52d503790a56d8555dbcf44facc93d2ac13d85620002964525f402b0a808ddf5e0d54477d52e58346a2015c30956560289df4cac6a2da2a53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9e02971f4b86602f0efa0cbb0e6c073b87c4eb41806ac33c536ccb7d9f6e732e3128fc4304e1f3a674887ded2ebfc6e08dea559da79233c885b2964832551f30d8e83d35fd46d2cd34ac07be5b9d108364d6a978cdccb48244cb5f520071ddcf6dc364f03c2ce858bf11f49f5230ad59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c9cbacc588b2f13269a02815cc72dfd75454d93a80ff0c31dd8ddc2dd9faceb39f99a6269f7572f3a9b22000766f8b2ff1250dd8444cfeef196825d86dafaf6346271f5b58b16d308bdc91f3abae362097beca02d2c9114116a0776f91004e666b7ceeb72857583dc773d4a7c3c6e066;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17f42a4bab13c5fc81213b0109e7bb3232e7f3d48ff3300ead42541ec1030efbbc317c334be47b95c3e8f4fb284579fe431fb538bf23670482fe2fafbbf5ecc415f138bc55b0d8e5accaf3ee5ed79a8d64cfb29493e2ad9e89732efa8eba9012de7450c41c29815bfa911e053187696e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2006783265bebce87b381fcd166528bdb39102d92f3cb397270483b48ac35c51e8949637fab369583beb71fa3f5b754e75af3f61d695f037170a74f5a42ca20f94369a4de038bc120e57b7db2b0a1c466b63203f22f34f9f04ee780abd8eea674a70f1b2cda72108855ba1cae53cf807;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22cc61f1ace0a7d3c16ac648df088472d43b47e371b6c693b3336f26173a0fd1c4cfe8a4d8ff589670a94055da5291340892c666e93cead284a6bdb519accdb314f37730ffa806fe6c01b1ae2a335990e8fc063c7449e662af71533221e48a0eb4ccea42c3e318ed9e070783a001cac99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e5a8918154fbd56920b9a4deb6ea5d00537e4dcd7e40116f2cd1e06c6244b4096073807132114e18f47ddf5dad7bb54d0ba77f08a4a84405606306e4b6ac00ce4f62570cbdbd1ab60611c7b07a3ee0cada5db9583f9d9d30fba1580416cf45b9505d6fda0aa32d01779ca709888476bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d699709ac8932f8e2e0d03157febe6533194706b805abbcc31fdf5783fcea6c7ab0ff7562053428b404944f0b473a82dce2d0e5729b5aed60b0b2c348c863f7e93f5d850ca1db0ffa455a2cca8f9a2fd9e71f287aa3d586e3ffa4a5abdbdcd4d7618f6145f03a61d06aa857d65a869b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3e64f48c652a5275de8d47146340d051dfcc41f294d22ad277f157b3e4acff283480f88cc692d33b4a323b82c94b34e822f5ac8b6d440b695f0451e68736d5b19f3425aae3af111cc5205e1aabdc86d1fe981f70af42a54e716e69af5d37aa08df4f63630385d7662e10ff28875b5e43;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5d7d913031e04b150565be585ab09ae405716cf031850847aa6f13b060e36b83bf9b30de735d8499bcdd6c0e9a3457a10844eb315565ec8e2bdccb48083c56550554fde7f188166a05e03a68264a98242c0072bc2c6294da000acbd3ab902b8222a1f39ae0dee0ce5114ded5709ce7bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3569c78ba94d4eb4c434201004f30507389c3fe7cff5869a973b4af7c4e884722516cb3b672b506ac3e053f6bfe5cd6ccaefba29e6e85ee7c90eac84e6573610aa2456e3418607aee137dc0423ee7588808d37fc1e4459321650ceefdd5c78957128e245fbf4855f9ed09bb2a1648c256;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c69118906b70fe4c95165bb7acb26d0ed7d71def47479c567c0a2232aa2019960abf4a4848bcaa0b2c052b5564c838cd7bdec6d1673e9ea75457f30fdbeb1d77e20b31be6f8a3d66c0fc54c206e3edb22b48783a68dfce0c6451dadaab47a48701ef80be574a242c7ae2bf780da34c46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5fd1168d02fb0dfc30357a59f322a27c7804066f13d3d5527683bf749d2c59a5d0468c05de4478683230c62ef8c86d3a511de18f298d0bf6b6ffc1293b29d7ca9c1fecd373f2400c0817c56fa7a0fa9dae14a466accbb50faf2548267e73b45318ec10758a8b8af8a1890af6d75d0072;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7344ba3890e5003940b7f6f37f60d079b5314a9d4ec61156779c8f80cd3815e9769d34eb30eb10b1a5db6d1c120a139403058fc9819eb2ad8abca29aee2e978118a47cbeecdacfd6dcea61572b9b58104d023354d6d1bb6105c207d44855326bf7c60341ab09d13c48320b2209cfc7f0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c0f15f55dbabc60a61ec07e984f126fc15df6120deab568d01f02225e9f880384cb7649c22aac48263061dae221490ea474a4ebcd6081ccd96a1a7ff7342a4c854287f25759f39865f7b1ffe14364f5462a8f933a2ee5a319aa1a772bbcf4bdd5064eeaf479a5cfdc2b259019bae4d28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h840659a6adea13555e8f143455e44c1ca43ee96929f4f24ae5f047f05fbf080a7caa76e69f77186cb790db5dc5f1303a54b5d2e2d5121284ae322d5410d4fcb586d9e46a95cb5f82e256d02077688affedabb2b13218f4ba7fa1fb2c3e43d1bd072f8e76f88f9923ecdeb3de296ae4b3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36b9f225a592a782a053a6f66165fdf1689fda9e20ad12d1fbcd51deac088fc92700d3930ff594b102b1bf0281ca89d84a3049bb143b28fa3ab4a74435dff96ddeb9067c741160852278e9691fc0a64239780e63d2276854189e665570aa35c11773eba27ccc583f216c87c2a45bc0636;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42993f66bed30e159691f2bbdff537b6656ff2cb5f78c8a09f43a55b4d739ea2b9939b37c5433b5bbaad77c3c4ad32892a46047b894201f405eb873fc2f454b0f0179522bc780fb3a709ea7e80c70a79064db7b096fdcf626439bc9cc6bf39a2243bd872a648b4b3275c00469afd5722d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h791cb1b1b43c253f699fc581d6cb4d08589cd9224422366579f47df9605b9b3ed163980307ad5e0e493c4e7fcf9b9066ce8159242ceb5cc18a2f9283af817cb82c51416679daf4b2ebef1b1a74d834aa383b168609172a4247a2f96975be222d8b8de116f458020856c97cde1cd76e6df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf48db506d06298bc91298109fdd64aa15d4cc00d778067f9c81224e2fc76c584bc4f69e6bcb5192e9056c78b6941486368fb39dec32c24def2b15db9076ab520b973375961c602e91ebd648a11fa472dba0a04af21211e291683d6d55b5edbe730c7887fe0b3a88383442d71d2793bc79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42c7bf3dc59700956237510a887ae8f677e2f2b24d3bfa88e1c1a27b700a056576e8c8fc5a713e647e57f4041ee86bff6e2fecee8b0771fc68b0a9a3344ddbe1a662a70037245a7a7b731a6ad69b0123e2d873c6c47b9d4d9ec2c6cd9972d7e052ab097874e11bb768c6baaa5f842fb93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74d92c635b0ee8a44cfbb1c51e83a0b7246dc79e791641f8e5ee62e164713f9265f0f9067a4ffc7a6d2e97b67db439ef6a8952df46c149cd550eee3389c108b7a3d226f98a6772db40bc5bbd49cbc49e230c6c77cd5034629b69ac7283542a04a2cbd720418b9a9cd5edf8bf02d8beed8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3c6d5e863b94dff6e50c9d0bbf951608cc3cfcd088063b8945144700d1a4d5d6ca5e6cd3362e63f4374cce6f88d170bba70503776c0c80681419c26f40beec6b7d4acbb091e99bf66ead96f8fa52ec49777c37e7a3c15c2c5b58db8b675fe07d76d04602185364a59c06ab38f74a6659;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda5983eeadbfb83ebb5ce150d5c014df9c921d0cb1412b1e8ba152758a28c357d0e95af42d85486155dd5a2bcfad1134c9c7c076593f357d9715de784d99255c77b4c8fbdcae17aef5e37d7b640282f1069d6b94275ce519693dad363bed6534c52c0a7bf8c42ba235fc8a732e15a19b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7eea6698ad79e32551a5ddc814dd7df04b4a0c2ad131e2e849e1c7f94d7804dce7b313807c93e0f949d303a3f55ca38bb9ab6106d3525d16aec5afcb7c2232806750d1eadb008518b814acd7953fe933ff1e3502200e2250affc905527fd6325e35a64141842fb6c53acbef2202d5a61f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h929c89fd4c58d3dbfd779116408dc723f2961ed9f9e2be84556b6798c39ccb9b37a85204e454d4b5ad8fff678a73f664cad139e616cc210ef77005c9e58bc5811a2e5653da2118c4f2dc8bfe0bef912165578da07cac64afca2a1c1b5f44d45fd790267e216062770707abaae71e0d04f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93b7d8a4bf4688907c04ceaa1bf31b6db3798df9f4217452609fd8ef38492a298c60ae1a50ab4402addd7312566ee628c8c297aefddad99ebb37c415d93f74ef3196663eba69038ea78bee3d367e03e2e2e939e3b8bb7ab5eb0f90792f6cf7b9132f4ee3c509ac95c8d6cfb2de0570599;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha60345c617452a9adc4ce7d9c98604e4ccff19e05d90a4d09d26db66f31d75f164bf8cac8bf46070d38f76fd208f51b9c90d553302e4a2718de7ebf3a4d9e975e75e2095008d69d08f2db8a143085ed2dfbd6e26746aad3305ac6d9971a3d196a9b1b70300f0f5b4d371d7d03ef7b8783;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h748ed93eba22df83f79e6658053d0e43ad09a729f85a9e2f8b559b2c6e3a6611ec2067735e288bf92f199753d963e218444f8d48839f2aff56f1ca9fc17be352ae9bd1df0d5d98ea1216214e30888ca7fa4f28c192f044134569921ab75770d9b32cc651f9ad9551b92bb5450b14c87c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd875d8b2f9677e63ea9c0dda1af3271b04b0ac2098200a537e3cc2c80305d57ecff539e0ab22fb06f09488c751a75de8cc5121db01d8fe32beeb06edfae88165af0242155b5361d6886c681769aa8f4c6cd2557f6dc7335aedeb8df5ce2171031673f544ae44000ebb2162a708f4a553e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bb2d109fc7ae85d611271e681e6dbb4f697871733f7075f7aea9ff92a38d72fed21dc8a002367bffcf1a22eadd205583ba8b6007536b792251c69dec3d2dc2bae8642fd16f844d52c835d933100c49a93b2a2cefdff6075882d3fd0bd837b46a2c01dfdabbd849c739fd5a5f1f97fbe1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60af1e165401471c75474170ff5b07be8a1f9be8add621b709244086aa28e28b5c1ce85cb031b1b465b2f3005fdf5b2da79ea409e5925ac312b8005bf180b0c23e87a29ce25fa3fb2f92c8bc591a48c00f06cdb6a7b896e914b62d2364ee43e69e5374a30238faa98f56c71ca9eccf24a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffc7bdcb403e4ee1ea0519ce796ea0f0465a9eadf12c62c06069dc80fb92bdadd6cc42d5866601e3d33395a4e9f53d015e81309afc95118e54073bbf36073d0c7448c277eb8cd4672c924f8761eb153bd30acf703d64f5e7a5c0a752fbdbb3293a21366e17b010b3d60e3ecdc78fea3f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac53ffb7b130ae6f0f16feae5116d11c28a47893b1d2b494cde4438c7243472d5df56d2ac9b0bed8c12d7234c0746f7e7c197d76ff4cf301ac95154a50826365208c217603d2f02bd86503ea1e32ae1b17a69bb614a3fb230cfa9382da73b77e0738751b65d806f75d0b6c598e4a37958;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h829c7eedd667159760b4ec0581be234b6592cdad0ff7f9f4110ed32b99f7ad1ea7be0d30db6effd4d6cba85d9c5858decab0742ae52d53af9e95de965c8cad365c911770f63992cb4a8dc1c6305e2fd3e77493b2554e299ae3acbd900f5d4bb7c46d54d54e60fc78166199da18e09fe4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d248664a6330b8846093a3f6086ff9d5fa5d30cf013a9956a8504b1a6fe26779a17b123bdb0bb81c35de739de39543b855b4da5ef46967111073d7fa902a15a2493d7594ca3a1fc5832ea0f68278846c8b87a9266c96029e1f074c8bed58816b57354ae8ff5004863fba32e93c553e13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac1e2ceb00e2901fe5c55dfda369666677fbc3a04c35d339110b4d39d144b88179d682bfa20bf7d33d06c3c8c0f68a5f438838d315bacdd762b2fcbff2b3bc5cc339b80afff9e4a062dc971b85c2a323b490bd1a4bf24d39d23d34742bd607be109b54d59d0f8dd5790099f7227fc2ab6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ee60a609637e81087a718d35ccf08202aff27f80353c4ad774bac69f65ed3f612fd7abe18a3b4a2e478c3facb832697cbe9bd34dbf1e34feab3c7a9461409428c87907816f71c6c7a6bf7147464ee2a37572f637c2baa27501f059a64a6707478925e5961eb1f1d404c83174e3eedeb3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f974f2ab755ee1240be886fd78a191f288f1f41038ab61eb1051784d906638a3878d5afacada6f67aae23e776354845f0263911ef5f97e11c9c31b488644cb1feb93c5bdf0b59be7e2a26a9cde20bff0c2f66c36555161d68a8b71dc6f12117e4fa7c207fe2dacce68e3644431073533;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98843c6339f76d2260cbe00068626f012df52cf8a7fd871854d9ef6e46ce30f6547bdca36e75dd15a47bb3b50d6d88a530774f77ed1ea88ac2b5951330869cf4fccc4ad5acb96fad64dbe0f7db89d7db7f843361cda7994b8bd4ad0faca0203f7a9052d848d2cfcb5fe8552be1679b2b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38a76feb03f7080090ee560e7045c69369eb7dc35f84abcd504f5ced884c4beea11321f9d1d04b502c18a34b5bac1ff4611b383e31aefe1c15e5730295e0faa27fa7c317ccbcfe441a034eb0c372ba992139b86df78c845299a6f3929fe625a329cd9837d54dfe2231b18b8187e6caeb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd37a8955797d76c17d7b834eaaccd454c204cb2f535097c88624ba7aa0a4c7743df13031c148b1b3b953b3eb8f20481853bee6f58f4b857b9e713756cf9be616865e044044a3c62848f9798d199e4cdfe37fd41413329d703578e7b2ee304a6b7f9baf9f7794e3b595ad1606718f87e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb436309a38c557e2df3ea5148ba300631703c34aadb2292f40dffa9bbb0212644cdfee99f2ddfa034f0bca3e2914140f4dfc4d31afd2142d4842e311129dd643ff7a7f117ba284f591d564578ec8bff4e5b7f9396a602de6fcea79460e0281e79d0088dc7d5b3b990c99203abe24b16de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f09e9f099b7d20078b54d06ef0f00f43075c8981eaa6f4d7d51336eb3c54582117b64ad55bd234c7130b3516604cf60b5d8ff1adf3a83681cf8cb95c157cfe63278b6ea5a185251293611b73e072b809ce5c1e22c8161dc35b9dbfea98f8fa5558e6b0713285f9680d01fc60137c6374;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7319eb7e6f0c00fb1e00fd311483e63c7d02ae122eea8030fa04e5909362c32980a721f9be8f8235c1e595addb26b87c5373379feb9aab92509963dd688e5e022abd5a61c246b4ff69de8e71887574480b9eb46cf4535b8bf1156f39cc956deec1b300a4de7ff307551794c09a37eec1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9a03e5346feb6ca20fe8b9d44623c4bf61dcfd9c9e098a749d92148ec6a970250ce4fcb479dd96071054546275e39fc1e762e31fd73cb6ba6066bbffc993eaf105c8307ad398c843adceb5fabe742d620974cf1593759fe99c605736599befdc6c77ba740a7772210e24b6442b3032f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbdd9b26c843e1de53fca480f1aff0804e3318293c66147408f0b2508e0d3e3041391ab009ae66d58a0723a1018958629fdc30ba69c3e978171c374c93e0bad1c823039b133b62ed9e9245c1054486d144a0c0f0122c29665c91c1a7892596847a1628d5a4c278cb510c3500dd6942169;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46bcdcc1d030e19ff192bd1100391ebd35d0ecc7852f0449be8cad2df7b96b41f00382181e7bc3212ca5c0debf3f23854c85d2ee9cdcaae0568c7d8ff8cfe74f3773d3e7ba96b7fd4f1dae9ceb0c6f7abeacbc1154579cb26a4b5e94cd676da3ae8147b3f53a92748557dcb6ce2a46e94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38757f5c8430198c4d41ee6bc91e39690ed23a516a937041629f422203f9c679d4860d558202ba981df23bd887da3716c8ab2d7a613645e910c581db2453d2a13ff3cc8fc7b20acdb942aef372977629551517ded02df9321b1a063dfe5b80686e8c526742ec100e2a89b7a58789584d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h106e8546199f310630fab149b1e157763a40ace04b46b8e1a9c62919f6fcdfd3bd28e87f6ed615e428703cbc7cf975080f629d1d680f17be6af6b7123c43be2f772bd2040a0b63fdc7fac3bc9f240347c499de295996cf597d5398436652000e65d84089c19eca020c95a2028b2b67227;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9ec6ee4256ac091c40cb5d1df69d9e4e4ef50193dce92e44dc77710f0bdbbc33917797df31bc52fb159a9a5ba062d176ac0b60a4fa8f174159fc18511a9d8c01361b7c4bbb3a4894f4fb9246cf30f9850fa605cc4cd7103c7c7c5cd49f99d58a92c9d34bb45658821b1abb407c15c9f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20a37eee151a2c30c4c9739bee85519cfe70ff6ac63e843cc70d818c9db77ed240da93bc163e8f8f01b7592e0f44650187b08af1dd697aa95942dd930f3094ba9edfb9bd147b9c76ea55c4eec1922576622ee96b18a52ac226e87efd44447d5ea1c2a12cf6beceadbe1e1eb536bf945c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb79ec792cc7390a868a7d3910e60d37b0d55b39bf0aa13785494e287c6e9c059f952d44759b1871943a223df28f1f01af711ae0cd9a4f99d69d93e1a0eab15d9e4b123c1b790fa6c8d5cd129854d7925024eea4269e9c0bbae6c6db4a82e8d2ae539f255dbe843350804e2345027173a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6995f35278e1822f9ff4ef6520bd6385612c9382a28ab250190061ee1e2c6c93d463820c2a5fc4d918aa7d419dbb2e5cf6cb43a702fc64a97211a49b81e5493d026e5233ba7a916e8d05908ed40111af7a52fc3d0f8f70d7e5c55a7e8065ef0059f4c82e2eb3fd069e661ebe6c283029a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52e132851f54c38ad4d60fcb3bd7e629db4349f3a465602e347db854b7c453b9bf5a10474356681f652c844debc0c104d6ab7484ded4e99c61681486d22fbc78d6aa39b518aad41e73b59995bf1c1aed2a00fa4e4cc463ed58e3275123946aa4aacca53f6b25f178acfe57b6712140a01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d9819a0c59053a2e5fd50389faedb7fd95c70dbbe876c65579fede370f2344db72a2415de23d76c95554455b7897d54e9009501128116c6e4191a96c476514407038a30212fc68b17bdd33cb54e768434ab706eb06c17ee47ced1254ab89c6ae0535855aa7dbbb21fbdc2c19512f50c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcfa84427fdac8c70959cb14a15f3c6a081fda766de74d761ee315fc734cb35007ffc81c77471e753fb0e19a1be71edb448f2df81ec4bf581176634dcac2f4270a727d15b6be6f67bb8368bfed9c7532d826370646bf99dea246fdf35060e80f3e19e9dff37ce31b1c28c3192075f616f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf264c08f61cb6a7b36f155c14957c294611146ce22c659ce99ee06d7dc029f42a60a170ff4cb48cbf06bfa7eb77f5a11ae2c59a6fac921b930803fc81697950f33310512748934f37caf770ee7aa5702c110052f55b4f5143799ad6df35ee4ebb02a4c431418ddce1fdc54ce6195269cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9e626e3f1e478fc89fe9bafbff24621c6bdc9d48e60fc4c20d93d797bd6f976c7dd5296151215b767c98894595d8341746bbe302aa7173185c02ca5dc52eafb3d886a2b9d108362bb2fb0a0ad16641b044cf88379b9eb4d88b6042d672f97050e39503b5f48378187079c75fc72131dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40a6d76d1879f82a2e4a012414918f61bf1cfcd85dc7bcae67383bfb633ccb4dfe6f08622307f287b2b00be658f9f3811f4e75d3b810d11fa2e6f5abef8a12c87de80412b92359cf5672c6b4082d969d7dc997f2b3e74dda627cb93467fd242c298f0d09e426f1a40baf8768440e205e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ad2e1f754efa2f9c8cae4a0a188fbb9d833fc6483f027a88e50cc5c6a217752ae1650dbbf2a73a17d4112c2c7045bdf0608bd7e3dec972751e78cc711f0ce7ec4af4b6b7c2905e7dddcaac1c6e0c7b367fa773dbb2f390c18044ab577a34a1c1497503f16fd5087d1c40c9b4f3525fa1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca870a5407435aec22e30ee87c0070b14bbf5085a599313333f91a379504a6072ad9c66c557378e3bd695f63cf4c735113fbd962e1358a75f03011a640951bb2e4a366a14a6f66a56cd5b0e2ad716634f28e38b98482ff63ba5eced4eb27a6babc06155493a8f7ee091a0a95d082eec53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce7319015d613f49a46f9d0fd225342b8ae58ce9789f9d8c4b5282feb2964bc7b2a3bf588cbbc433b37479f7feb6a77bc6791ac3826c114c54db24072e206e388bf0584bbe7e77b090490541166970b48c6afd5f9ea2b4a1c11564b3f096eca69ef4491c56de6019bf44491e9f8d0f017;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74139d7a95f0cf19504994d261240c042e4ac837ed040f16175b40dce9360dd7fa4684ce1997b5c6251a074619d86a0ff7b6f62d2bf22c24f0b47b3b19eebc38065e3b0736a509b1f6d9e7d4767e6bc43567a9c853a07adf8129ff4e2d05ea6c9ee3b378cf3c6b1eb43454630bfead2ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3ff37d2ea0536b035a3c69286f91adbf98b51b5ec1465557d98159f8acfa9addc7f02bc29419ad14da9fad9bf109603453a0ae592dcf59fefc271574ab0734353cbd9f247db886a9b5cb026f64ccce1ab7e38052fac3853f7b2f40e47cd322b8a1cb4e119532a3f00ba8d6c5ccef9b87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f3929a711fb1f3432d10d64f1f36db4c69daf6c2dd52c80fa0930df25ef841ee6f886254cb1a6401b29e74716a162ea3f6f998c524cd9f48676cf4bd29864e237e67aaadda12ec5bc67313d4e6a8104fad1fedc0a078ea15be81d3924f04f41ff449f39a912f2ae05eb1a39bf067ddd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc76b580eda9259f89043f641ec94e3c73ac0f6e10383f7e92946e918283ddf26a63e66daefeeff02b0b342b764b8f99ce5c146627b2e347fc2207626e60bb18dfcfba9cb515512ac546854258de8c9e1f2fa451b843b2e69617becec7204f1678cb25c7b390f453bffda8b4ddbe72c1a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfbbc08dcc1f6aaa680de4cd2d11c3666a7fe724cee92a39e42ec27690ea2a9c1650f52e62165e5159cf3e7e9db055792b41d53fb844a712b19f0f7ed704b6ec314eed64d6ec1d814818e1d1703bdefb24be1ebb30cda34a0b6ef7a2ecd930550614f945594c6eaf619e4acb79e2f936a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cc2fb25913c17ee9465d8ab8c982ecb65cd55cd04f59c92947b87ff9e1130d6ac851d33e422b1f4cfb5b6e33da9fa4cc4d644553800df2119b16debf51f5721fa5997a87a92f9a4ec3b565c71a6d56814626d5849fc2c07f25ffd5b1438e7674d61857edc1fa1c5f87b156addf32c340;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb51e10bd970e352f950f518db9f410ce4525784ac75d8e8768198534e3fd710367c19ec0a880f84ee228c2e57ba9130a6aba56adfb96bd7fd68e447614b55c2a9319698c12f64184b1c65c69e807fadc02e21c492ef015a273ccc2853e0dbe6c4ca1d3f459eef31e6393dd6af7888dda6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h414df49235a8afd790d4337aa5e802f842e558cc740d0c9aaaee4fb6863f99e06f5510db3dea63e93c87f9227f0db69a91fabcdf35ae655a3763a805187af7845b34a2bfe1c834dc58bbd04d0ced8e8a90307786a47aeeb9ba1327dadb1b5ac76600d7076ba4fc72d854b1c7ebc14f41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9f6376dd179cddbccb694d049c3c2b6b3a6c4f73894f7ec3fe3a7de99ddec86eadf328df6078695cb4810cf5418083aa9ca68c158b9f68e39fe79b25f52add9c854abf407f3883d7223efab143d5ca0a2dbc4b9872648ce906277bbb9297db751bc80a76feeb14e78504effd3aa2fd0a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c7fe80e5ba3425674ed1436206720f0b81d7aa78d8d8602b688ca28a7a65c901ff439c739a114889b5957bc926b851b35aade64391f4b63b7656686df434ccca3ca2f350a23c8a444b4977f8ee717c900b35f29b627163dacb4a0a86ef2a4776a151208a8d344c9859355c4c627b8edd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h788a2a7de1e0573c1fd3ec23ec737492fc1e87d3af96bae17f034b0e72580c3bd5a4d3832b751d3e5100e096551b44e5b7b4835f80a89ababe0093e8010bf3c705c0f41828e7981865a57344e659fda055cce302a6e50ca3540727047eec72fc12f7a7119ef57cb2edee741dd59528008;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62b9d549e45a5d4a45187f52d3acf6a08a61deb313481cc13e13f06bd8e0e14dfbf4d5c82b82d077ae0ca34a8faac9c74d87d6633e86ea320f44ce60a1bed81567a18f1125982fe94e77278b6f53bbe027484ebfd4f05137df7b285f252244bdf1dac7bfdc4c9e076fd11446d95115df4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb27cc7a31c2e4e352db7810402e663d6d160e5460d889018c091a303d1f9f873d7701a706b3e003db6d66b3ae7e3e1722bd4d0d7346f58ad085c8f9044435e0c5e0525ae679c13d63e371f2e5009ea1d29905c65076a93b73412e2efec7b1229733e620d68af4ad72436301aba0b4c06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4369c2a4ac42f6c7fe334301f393235e90dd9185fe3f8d468ab84954e1419aef019ffd8a6fcca5cac5a364a52f5bbea23962900683658c321be46d7e4b8c2e7c88699f17e0fe93a42fd1a7b45e53e56e9436b8f8853566c6a312931addcece853ba0cd0168d5167fe84ce458bfdd6b7c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf244f777addc2814c12d1492897e2305d277a12c7a8f1602415e088b889018e644237b97511cbc087aee47d6d1005d06ed81a891a81131bf91af88e1dd6d13512a4398284fa4fc03ea662009727abf20104e42eda6489d7787dcb57d815ea310b830d5d6c9c95ce985ab37e79874ab7fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb4f9545c1ee5339ca797f495b32ce3ea62bc698701de1ab617a385905563c9d7523718c5714c253d03480fc8ec338940d7419577510b4293c17ddae5e1f62c23b3e35704d45db366e9f4b33d050ad49b7b4ff1526ab078b26b969bdb1bf8a25dad8f989e4757fcc83b532f0a79fa5e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2071502fc01ae6ca81dcc527abcdc6ae35ea9b2dc668f4ffc6fa561438a7cd3f2a16bbfa8f3ace092f618164b49c689910769c81c745f8c439d1b4ebbfd158e846350d788e7a7f8637fa9a3b37db04c5798789e9ba0152874f6ca082a349ed791d8ebbdfc1476efeecc33bbe3887167dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27f08b0880830c1c9d0b54d499ba3e9a8711b3e245b846ef287df1e8d38466d4b5317e953425cc73916fc60a4917b0917836538a4b7a2d7cfea9ca81b3925dcef989ab2a9c11e9b7bd9693907dc0d46367bb0a14fa49609c1bed4f6938bf05f034ee71bc530133e7e9a4290412a6f1bbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb78afb2597aa0464fee38198f77d66fdc263954899332f71caa4225c690643af5d37e22fb0e4f6daedd149792e35d60ebdeb7d98c1dee2b3c901a830f116d459c26bc5efe4af01a9bf698679fd6d3c431d7db41c19c4b343fd675b5f0c8c2f98e5a02d28e4ec07989f636c04d9207a7fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce8871f424207b80d5febc2dda34872894980bb6fbcd31903a81c9e0923fef0106c6e796d95f555a7079dfad6b8660fe6058b55cc1c82eef866684a5b6e7839f444194d11feed01a8aa655264c59714c514de5525b517865084b1b9c6fa06ef2039f17b5b0a33657b7adce5c88b55f943;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6c18aee7d0b94e7f9978e538f5db12fb89e6968ea5f27a55584548e8d6f0f91afc60833a4fee770144551eb2540f00a302d37722ba2d865780916ff90ca26fb74c4a1a98d25352361160b3719cd9db8254810de7859c556a0130fb5029b6fe3777b34d97a35d265ec05dadac54670280;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0007560bf8b9d3e888dca4274ccb0d625fc4fdd53054d7be4f8ef1105a7dfbf129204fa85f6dad1d012049726be7eb296c9c14ef358568d837d7f761188beebfb9220f5012ca899d403f249d6274247092e0cc1d0c894a3e8449361d07a51dfe4b8d73613116982849ec996603e017c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cf2afdd03d49b0edb3e8b35223a23d0934777b986d9885f3760b933158c7cf33bb82df9cd5a8b20b8d65e4b6dac8bde00016b1d3f7d663bd773f7a8fec3d3ea4835a8b626fbde17d43178c3247218c5c9d65a6006cb0946d7ae33b670747cbe023c1113871c51ae73b775de072202e4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70e5d6ca6de4480eb99eb51031fc98bcd1332cfbd9dc215f0618ab64353f0b36a7421bc4741e9dc0fde477cab7af169d5ebf07f29c14814a037d0f2793e98663541353504e5b24aa6193828827bdd88f13a0c410af367ead543ce97185d6e013a47d8763537a72ec1dd102d27c7b4a4bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58af9a58cf4bf898a29724b0ee4103e8f70c8d1654361c1bf23be7d00ba4823a28a2bed45e979fc67166ffa3d4640914a804b0f35a23def579bdc366b1c0f8d0723f801d7735dd08e572a0961ad8bba6eb67a7e059adcb212f4d0ae0dba2442ef795d075c26dd906d2564092ab9493ea7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h130dc3ee1637d3a2f9519dbd142efa18ebfab296b3d242a0e5069f56c1050bf65b87a8d55e6342218e54371b2688f2831d07a2d6cf9c6120b37712a2d4246f5044815ad850cea7654dd5c1b7a4f7f2aa229a69f90ab025dbfb01befc3706c342236c8f7174ada800bc18eb1bcc4d6973c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce386c07f82c4a7c03f8b8ac7ef1f238834970bd824dd8aa1f50d0a0c0f2cdbe26a4ed72c09050a95a85ec7813613c1c4e8a0e4b9e1147fcbf8571e22357d14583122f876ee2868d85487a708a86c691328f6c2a21848c0f2508e6db24dbd955f1732b9b9b0537df75993c6d63bfb46d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3dbe791404cd2150f208cd7d3185d9992573961967df2085a7188f5c58afb0add30c175772e40861cfe588fdbbd5b33003c050acf88b4ca0bf54f835ed2157f687ff02b4e5808ca0e8062b7398fa055340f021e120d943b8facdb5cc2e818a1cf99d36c7a496c07f86c364b3ae128a6f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5e3fe8f3a908acd39a62ef00dd4e0b517dd21d8828bff4c91376a5ef1db4099a9f8292f22af14966842ccad37632345ad5bc2e1bc9d56b61d58be10f395614e15dc00d313deb1dd92956dc1827504cfec6a558c45e99991db1956ebd937b925bd3e2347d1019afeb073c666062b8e3b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb4eab5d23851627d76862047f1dbb899f45dd7db61ec5148dcc1f88686f70a6e6cd1ce9fcfd0ca3318013e5061e60bf048a70d977fa1893e5c900d7466bc402094386f817e47fbfa7c1e67311862f1494461067e14089ecec43a2412973bf853f54f9f5d4f25893e7de498d97b87a6f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ffb85d3eab6a1bd870a4ac9a8a643d5869338af4218c513d1102e1998ea551a4607dadd04aa08df90a0d881c930f7a0fc7d16ff193fca23366b97431550c0d913811e135cac2aa50ad0b82d699803fc6e37f659108cf049590e75404a45020e55b676b16fcbc38b978eb8ffe405e8438;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd0b12bf91b5fa42afe80cf9fb2cfe982ab103092aede1d9ce70ed1c25a15ab6aa95682ded8d4535d440992ce37ed1cdf4b6df59c3790528c03e7d52ef28535068a23d6daba2e0b9e51a9dff364b55e39b0f1e2da973447c3164461de67b60937372c83d3be3de4dda0de11ddf597ad37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbec59a5b18208a62a5d2e6efeff881c5b5d2f7fb8113e9d59a015af4bd819fee793b737ac878eb199525ab997d5677fe910876baef60062974155fd6f6c43a53007c07a29eee12fcaaba2c440aaff3842bb43d49f11c6e87680ddfd6c2ae90a33ebb9b6994146b072d87b9a02cf731c0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb59be90c0d30db7cb0055981b5073019a5e6cb84f4861b987d8782a7684cc30af7ffa6f1caf169c880e6464dc23a309b96fbf64fbe4760a8881b49febf043271678ef9bea432bd803254a1fefafa4cd52605c78c9264427fb2aa7fd7c0cd1981b2e23b81fbc57fb213b074d01f9e0c5f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd50154b59117680bb31e751ae21292fea396616b6b065e7c58d2d7b0a8520c5612cff1b0171c5bdd1e3e2957582f7d7ffccd924ea5c6deb793d5567cd99a29d19cf02447643a52ca87215dafbd89db937b35cba818152f3269dbd036fd7fc4fb802d34f12793c9bf8f6ede08f97390c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e811f803257698ee1839b6e1515fe16b0919c5c0cd58af72ff37ea97212063ebb1e0eb7bbe1b44fd8a302a155646a0f3b4761a39139f5a2b47f002fafafbc57567ce2b98ed9458970d83665e439abc759d643c5bbdb55b2beeb3bd06faecf23b637ed967768e96eb49205007a39a3c93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd947098c1bea96afcc37b0792b0cefa65d648d088af629083c113b4ff74708034d996adba71bbc1ec76cf2175b65ac71c19eabe9bbf773ced3582b69d0305e5afb7578e7ef9117e6a715b1ccaaab35727444599537eca93e3a458e7e34be9a490caa3ed9ce14e9d35dadd3cc5a276023;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dfbdc03f963b8709beb4b5e3780ea7b5200f581b339ee96ec6a14e83d81786fd8628b094c52b3ed348cc074721900cdf85eed606012e46e344169bbf304683f478922e6db77de7d1aa75d3a5c06f53bd35b58fca3940523941a79a84fa8e3598e93ae39c88acaa2f70d9a9ccba7f0680;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cbb00f75907c93349dd921dbf9f0edeb25d6ba76c0cae68c19906e140ed3a8ff2cc3ae5cc90e0f56791714b02b59ecd1ecb74f47d007255715e6723fad342cf3b66ada3b7d2c29b81d6783f37abe6c41a4605337921ada36d9a99c7954df075ab1d457f9737516828d76b247fe0fe8b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdebe2d539d308a5ada0973c66122588a831f0fec5d9f9681be4a544e4dfc1c8b2d3f816881a24b1785a977abceabdc9dafbc87d73a42fb3c7fdbe6154def29da4c402e23b1142e73efaa02b20a243d307f5215ead5f4fe61c433662387c137983a2e4d9f5f6dd81366ac6996f23f26d91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a582ceaf1ac9cf5737b37166a9fc62383e4992271ff0a0e75ef8d87b6e22995b7b715de4b1fb640bf82f3d6d89d6704c8c1dc14feb60abb63b2f478ceba3a2c59982d438cbd929e1a5804bfd6f54bb75eedf72af4d9319494cde34fa628f5b943a85ff34c27c5007723f4365ede82602;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heac4faa119fab0cc28bd74154ffa7ccbf1eac2ceaeb8a7005663d0dea7249eb395aa852039bdbe1d97f8606932ed57f81736540114ebe760b421339e74f18a33ca9f1778e44b4384315ec9c9fc5fb5fc5ff77c01fdc0d0c4a4138b209cdee9b401c155df301424c64e5e770e79dd2a079;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb43879649a15e86e2af90460adc7716a9a9ced7bb6b3c11bb387ce723e38ec1f96d74756bfbd86e84079b86d73f660b427c7da75efab40ec1417a6f94da0b0e30972b2f94f1e9e7ee3933b80eb971c05039a75f5052256e57f0d5f2cfead75ac944010c6de443f2090ed4688fde6cc6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h737fbd60e776107c029abca14f321bcf916c673e74649ef462370d9598fe77c2d9ccce7afcd8c6c3fff3af27b0d275baff191b96af6083ea685c35201ae39d96b84a11710ba9a7b09b794c1e2a26d6a7d2edeb64d329de66e932e0eac466c93b5175964657a9dd39f36e26a5270254e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2da8ab21d88267acf6fc632b01235d8582d3ee108109197e7f199f25ef1d30b9b82c4e3ffe4ffa58ea409309c1c0718140ede201b28dcd3d6ed3edbab60a9b408f6d96a9d601b93b25c0bac00c81cbc9b775fe1455ffacfb3e1e97dc1adc7fc584e09212f4fbe78a532df8096fe0d9035;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf71c3d348fa4a000dc482dc65812fdb63adb2322f81b427dcbe2332e70324121a09c69571eb94a327414dccb55eefe26eb0c66245152a0234352edf9570924358617d6e0bd6742d7e934d4fe565110068f853b3052416f3823ff00641cb6a507d21e55bf26879f81898b5a55f13d91b33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1371ced722b2ee72c49981df951c2da677bb389f37edce20afbc680920868c469578e095fd7a3ab52624ef63ea0cf8ff7ed8e2d2a4e2f7ce8f757816f0d98c91935dc0b59f8c8c0db19ad14f183fe68555aebeeec04c1e7e747e5fad2a7e2864bfb7e8b0c8a7d7859eccac2cb6c16baae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1cd5256a3e9ded081b3626ac5ea2f9a1c2fb0ebb1d5ee627d4920d437cf275a438e16e11bc2f35c2571bbfdf82dc56980892eca25b547ad6cd39d3cff769b78e4789d019b6f460fc8b89994eee341beb79248a8f9d1da14026c3d1a085a81adb027a6a4d5644b8b1c34562206b3bbb05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7233eb735643e4abdcdbcb72d6c579cae097b1f80e6890680fbc03c1e60dadc930e476aee2aa04d7b90fc270734afe8090e50207d3994efed2ea74b7c5c04a34ad5392157f78bb10fec9e5e29ab7964f84b63f9c19baf02b250843b77d809add82fcf3e20e4f6372bfe484d3f967cabf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bc54b3da9cc8a57da2b1b2a326101c57e028aa62b1194c43c991d4e70b7eae7ab20650bb264853bd4fc60ac0fa7f31863c8b22eea8d72bf70a8509d72bd046b8d8b56e7b2e0358b1581d7d92545b897fcac70cde72c014c61f4f7807d8a412177e62e350c71cf2bd8cfb940eb997899e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38e243320ecf82db9a6b222e74cb8eabb1674c8994b7773edc176c193ce498bc7b8efb84d6346a45d49d0d5b9c28467f8ed0f705e14530c02c0703c7cdd69157876d6bcc4922b041a2b8f67cba3ea353be191de5fa734b498415529cfd7c223d3f5631b8edf86aafdcc84041044e42f89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h368bd61209ad0b0632aa53b0503893d0bb3f85f7cb96fa2ba26a985e9f44c922dab91457ecf325753b1a2c16035146a4f201356f6bde8b054cb31271a108a4ca38a5b885c99c4ba3652e9f9e23e31ec363f3279bef13bf6499c8d4b2bdbd4a489b711ab3705c129308e71b0805ccfb93e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb183e8a80af3e1dc282c0e565059105002ebdb46e10ae70d445e01c27db611c0f828045572a589c07340fd1ab1d5775d564b58789eda8c1ebf118fa7a5fa5fc48111f4fb58cf6d912355197bf86e620fd5f7bd47330cdb8a41b17fe1822927fd1d3b7eb34a9451db848f29d88f86d589;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41fca6cf60278ac6e4d893567e03a697283bd922a96c84b22a96eb7dc459a78bb3b474ef37b61571f252207132a72f34a27d4d970efb1b1500bd98bb29cf92e0c817714fae2956fea04d96c00fba4cc143cb338143628153fd0bc6c680a8aa4a5a77e6b3fb239edfba50c8843e91abd24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1ddc0822798091d7474df9acbb979459a28f67a1ce69f75a0ff931fdb26ce70afaeab7789389972971a624145abc7cf0d650c2b22672d96a6b806eab578b153cbcbc34912b65a2deb14d6ab047a3a3260d8124d9ff5c7c38d53a825ffcff7f0a927e05f01ccdec5ac404881f27caff84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fb4e57ccee801b84ad5757d06066e9806955a21ffa0a411962682654c8effd5e5b6c655d695f44d4e054ca8a90a9ade1e79d914d819f7bc6b6e5e37b14aa68740e971940c8d791bc628deb093906a9b84bbe43c19094c448f581e325aad9e39abbaafecd136cb59707e94eb03ad8bff9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae66026d067d0782e3ce4c4976f826a5c5d743d712f9969519f242593fae92f35f6e584cd46d827a2860b6ebbbc66ac0e019309c83d12cf43db39513c75b96e2fa5a92ac6c9e075bbfe2822b4e962c81a1a803c0c92f1a2a328c502877aa950c246a30088500f5d2dc1de8a205474a377;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haba6dc2e0625c5b70af8baa30228d4ae8155fb29d6d1cfb0afc462ebbb672389d2772f23f55ca30d5748b350f01961fd92f3eb8d5543c4a7196356838636408664120eba724206ff9fd35f6cbadc03e6e1316532d529b5778536d3b23dfcbcf1448bb72808ba95d3b19a4251a8969505c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4a9086e10a28564f931be6ddfe1bc38f63c9439a75dc682eb3d21cf817f9b9b0202fd217a4f0e93f3e0515695ab79b77acbce57914327308ff6835da53d697f05f7b098daf654e6b82557951bf0aba5dd9752a2a21317123312e35a2898d422cc4d9f89bd001fb8de40308031ca0f82d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5944e82f871df85817f8ded719cd6857513df8e67097d02682db808b2ee652317bb8c3840b4ba5c15e0cb377259c525d811f47f5bcbd23a5682c8797d1ef2f7b33d0f6bb3fe6aa7e8e02a9223f5555b8f11a3ec08e2d00c235061b1ded3661987c8fdac4cd6c8c37dcfbcec0cbad1907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22830d759ca9fb4cd4d7330f4e5ca98acd70c8c4dba661fd0b6706e6455bb8e3534e984b7b750e2d65c987bdd6c4a03ec6b5d330e9c5df92a63e118fa84e5b6460884f20ff2cc514aa90135950aff2facf42af9f4a3b685d7fe083f5c77bb37738e6b7c5e2916320793c895fb5025835c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ec00a820e7c39b31d6748b6d0aa1f7ba110a09f84711267bb9bb04de12f243d3d725e954d664ae020246d9e1929bc4affb2e533f0dbf96f80b41f4dbb135817501b4f941b4b66940aaf32f3489d1bd8228b8237ba60fc0e7c5ebcde11ac712cfd2f642daa45ccda8e6a2ef40597f2ffc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15ccf031cc19dc2f66d1235144e5351ad5d8900177a60a66674305bdadf05eebeb9807382598f66adc1fc790dc31fbd5a8195d74d5ca7155f5a75ba8c31c96b095928bf1c10f41feb7574ed1d9b27ea356bb489c76777d59906189f697fd07fe579f4d601d1adbcad791025d1651b6849;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f356fe9580cfa6fe81e3df666672c854bb34df0bae1f288aa78611069a60feac3a46d1f23ef31155fc211f054596d914b1bc69a58ed15512064c1c675ad726e9237efffde5687c4c1428f146d8240cc6f7b2dbcaf28575d1953c8c679cd584e4c7b8f1fcaafd3fd7f0b1d3d6307014c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h765f9ab86ae73af010052f13a68d5548dd4c7830c7b5158ae5c4a7e5bdf1a75cbb99230887d9d7bad177418d220c414ca3a3141d56864edf66763ab96b831f41f790f9c3577165933cb64f828f85e3d3296621133d7911b736afe32210882560a2b155a1a257d992358802cd491ba2226;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb03335d12ec9f7bf84edd6ef850876a004846b72693c7d3efd61640d822d86215feb4d75ce429933a0d062d8e241d6b042b5c5d388b40e57caa2f2cbde998e43b4fcd8f031db288bf8145f32c4c2ca0b73d5bbc09d6a904e5a751b6e654b838496224e0c2a4580026dbf73a0da8b3dd8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a697f30ee029b30d5d5b1b01f0f38ee255b30c6dde96b67c3295abfd4e9e6fb68a848c39f8de27cec5d9a85f3370e8a460ce7e233f88a4a0dd5c16961f9c09ba80de987e0b85b50bebacc9ae034b952a7e08f742a2fb85168dea23898a29e320f47b03b7a228d5cd9316b0098674b551;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b2d6539b72b6fc033c8d1acc7f85f5c441d4c7622b66858f51974f64fd1a6316966381a1e935012ac2bf1fa2c9910390aae0a4f31415a81b017e1c2baf2baba042cee3059349f4fea1faf1e7747e1f2f2bd6e56b8db812f0679328d69b89fb06288dd93beec2857a554d57c91044ef57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc24b4f64f45b2cbbe5179d4fabb6fbc73252675d5c47bacd28aa027a77d6e3a2087a42b93420d6a7a17f281875a7c808f542b9b27ef7c0ca80716f92022fe98c850ee4d23a4ff42585f08e8cd4c64a84b5022eefd366657edeef26ccf2fbaf6bafed8f319c5db323accc22f64e160eb5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6e8b384d83b89c80646434e0da63b25439db106f4bedf3cdfde44bf094d0beb47e051d32d797faaf901e138935554056ae5ffc96fe714191ec59781d4cd15241638656a704a55c29771c6a896c551dccb18cfcdd139b0db34414c8c93fb4ee3d13c41b36ed71a3d4de2c57bb5a72efaf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e1c938082f602649a94a4fe01450bee0752291729259e488fdbadff71798a425b97d75c879de54775ad51fec23b953d993649622266a700224ba9f9f771add38108da260937e8efea168296527b996cb783b9f65fe7c189eb555a138587ae06c495cbd27289760838492a33a9e63657f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98033f614769883ae1bb92ad43a9a3bb997f70ccc8ad7f711285be7a3bd80e640a1590b7539a343c70ce12f77c019e4916cd84a2ffbf78ea7e40c2cf561169ed8c1b8796cf1483b620a19ed68b72ba76e45ac8b191a0dde9fe624e4a38dcff5073bd015560cde56a1518fdb15b49130da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h903ca7221f82a0da512b530c353b449d13f661e4f00d074456911e902dc998d9a6ccdb90df1003c6629df4e016d1d9ba70fdb0c4aeacde8810283c7b4f16294ec19df140b3f8afb1c7744f015a03c630eca176c138264971f3ae8c747175cce198f96bc8fd864b9a84c2dc36312a0cc8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24df768632c7055fb85cc08f29de226d9bc895d9f1fc17619c55040921e2157c802c4173efdda6d7e2d613b87279e297aa9f9082ccfcf84f3ab4430af293de66a89926b14402346ad7db938e3906444f6b971845622b53f4391e55b57251a3e0f2588c1eb3e4534f461782de2d24b6b13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a752d3a333373cb0cdb33f835a97e551a88bf63102418f68ce7dbb045cc6369b3e2499496d84f754005755f007d57f1dc6bf653a4d13e16f38b264afb2e5b0f16b09b57ebf1362830555d21895ee44d4a423112b256de7f6743edcf789e449dd418d0cd9096c2f9a871406d598a439a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h389b5a2fda7c44a5a813a0df607b0dd53216533530a67f4038b8b5be5dc7507dbf5086e2378ea8dccb129667368595e774895d179edca5d39f0ebedbdc999fdcef5073cf19543ce546311f2b2549b7bc53eaa19eab6ed5c171a3f4d13203f3195bba0fbd931e820fb086f39a708e79ecb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7489716213ecb896d86bcc9af833808121edda91fea7b35165606910e9d8cca96848aa3a344785eafb7321cc0750c791e33592b02bfb64c7c10531289a0cc584af5d508ca889e9e3f2d9bfdb3cc91a84378501beef0fa533c378acac4ba1e62057f8bb2d30c3690d8da95c801c1870ff7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cc878ab5d2c4609b866417e515672ee116076b13b2d13e320f70277a32c41a2e23a6b09a28d7547d59b83bc6f8188be10c2fff0ef0d475a555333a0219d140bc6e9bb7a5c9dec312ea2e51d9aec33f850669ff9417d38144dbaf8f2feb34e31c00a584b5f7bd61230ed704e86270c51e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c06ebfe87ca2989e9178581bb1df1ce96b74406c42e5ffab1a0fac3196fc7a558ec2b446d607098af46b45afebecd1c1d7356adb99eacb7a5fa31cee4e241394bec7c4e8d491760c4831b02285c891015fb9f908c97e71676210927f01e94bbf38dd1505da9acb40846ca16214876e28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3d5ae57f42e10bdbef3cf3c36e1d8c081d75ee1ee1734585d5a7413b452480f6e30050cdd193975797f8661d37bbc649d99bc924c4ed570b1e5aef328f98b0e7bfbe924712f88758b187cbfc73d15e7751559e138d7fd4638c0a1fd4a992e798a61b3709d4d5aac49122fde31b79b06d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h748387fa10b97418c553381cdf9f97af4db34dda48691c9f2eeec39946212ccc37fc7c4712b18871dac76948da784e225f52bbfcda0b559d3472ad81566056179099234b11d187ecbec16ad2794bbac675602553f02944116711aa07f83523e0a32ecb2dc54b33573d0699b4306e3566a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14b29af72552b44bf6a91dbaaf410c4bb37fcbdd2aa93d6f0f728e32b6c0f173c76040f87dc7598a1e66fe961c34c1fed0ae2e4138312206da9121adb4c3a868083f702b2f9f84b69d8ead210c201802093288c031423bfd07f10ae80599472bbdafba2b12e0cd6ff6cb629cf2168f964;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda5eefb39bfa29026ec086d6446078104bf4becea4da7ce5e7bd12d458b8e6959f9cac178b8586daf44ab989dbe6a9d1db6d4fe814d497cb9af064cd01ded872ee81081291a26da28bdb874b9e5ed5f36c840347578365d7762caabc41eadac533f01b6207a149a91187f681ebddd9a1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h304d34ee09ef6da69f63d5a65eca4de2a3375b20a25c9e3e7ee7048970e0cb39dfec404e3a7527da0428217e7589265d3db88a1f91154e4201df3aba2bca9ff394e74706454248237e93ca2761a523396d0c79b7ebe86db430f61f395d77f6feb8e8a3d483c2031bfcd1190c52f0a23ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eb66ededa1b103add380ac75ccbadfc7d39fa040c4a9f0dbd054c3ad5e967d3297fda8c09f7a452c37294741087046934e9c9068c1a78429ab2b3359e75a7e49accfd64499eff07cf27bd0b9945358d526424495d95349e2cc10f2a9b182250c915951523f48178b8dfe77c28f35cf14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41a365579783bed3b1d1f555039c32db56575383622231ca32f78a2d5a6af17ce0cbc203476a72bc175448185a88ec091e2bc47d6ddcad69e264a7e49fa722990c745e53342b131c8b1db0ba846fd7394c34b57dad753ae0a6d08c33506b741eb6b19a4cc89f3eb1059622f42d5c5befa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58932e7e6bada257629df5de7dec7365fd50c73a4de01f0c086f66b680bc6122918a83f5bdc1d7f673bf8213b60fed0defb10176c863e1439c87a441b8d6729e49333c88bebb964136b0715d9233ce7c421a845d81ec7950ad88f54856490e1c1453b285cf8c0ad5beaa09ad3d69fab8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3925a0959cd13a6cc5378ba1ee6fa8933074af3e2bf6566cb404f8ee2c26213c996ad9d7af5addb028cdc5e22f487b8f86125fe948187e4748332cc5eadf293caad6735828cff8ad77259c5ab84fe9b2b80127f9c541e7369b765589b07abde84f1456e67c2dabf8fc01ae90cb8bd29f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb07d20811ad70593d313c19927198bb614c8c64212fa7064f18833a87aa04d9fc5f9f3c7037a2314cc7a335ed8a0221e5987cc0aae38a424de53a45f0cbabae74c7494609c5c4ea2b4f77c43a416430f0323413b0fbbad4ea4ff7dfe857abb4a64b53df1bc30987af92f5f18a4745de00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he59c5f0dee88b09f7149be2ec87bdf3558d4f24279fd17fdd74934581cd4ebc53b0756e34ff4ed9df1561885b0c67db1c9763b81b7599746c0c63e98ca2f0a4f8e8eb6ebfa3e4494a047babab086ef1d644802998f174a61aa745515c4d84c03c0ed6fe60ea17226a13be1b0f88b7b2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1b9ca9a7566b2cf19f304a73c89d5038c287e883fdfe8cb24b26f7fbeb341a8d9b6b46c728586a13e8893aca9ad2d67f0294164e243451f622fa7a8f2dfdf83e9bd595a6213c58f79c35bfd86ece91e9bc43c04c250ecfe7fe7f325ea15ea4898baae00fb2ac1f7a971e594252ac0a44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38fa5fe2f67e2ade4a5087f5620b8eb6e8851bafdd4dd2ff490ff2553dc58cc385edeb43723de1ce8cfacf638164443cead04f5d911861de72d660a3b6b5ee2aa6afd36398db5a18b6591e048b116fbdb91781f967c1b5348e678b258bd6cdc1e1d4cca5b20b1033164046c874526beef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37e863608332d3bda0691dab95b6d71c5eed37dd3bb49b8a8ce9865a0368de22d81df117f3e4323c4fa7a76839cb1d423870f478d78050e78506b7806dd2aef1ab35b634f7577cb5ee5bf7271a87e684d7d21ffe665b81107c0ac3b99c30ce869354cc4f501dfb9b884f5cd24328fb81a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b4bc7340770a3ebad5e8a36f7b4c4abf6eccc0172b6327fe6852190d5bf7067fb78a9e8f3acf7f6d536c03e6b5098f7a571e778e493324aeff7ad258b1039e74dcf2324d46ada6474ef4af10273d0aa8d394f9c711c4155bd4e4ce5ea476b94b9774c010d7b80e4fbbe7b242de49948f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h279c6ee0f0479b1a7660617c2f7f26418075b45fc7a75dc900ec005fa357195bc4f8ca34b8d4732da449ddf4c8b158bf1abd45c95e121dde84e0fdfa733f40e0fb25e8b636f244b0b585005a7baf7521daf892f54b5c63c0077bdf1e09fcf44d51441eb065a7beec9bdf78f8c0af25037;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f5e1e8964c9339e4912c1894d0a120539a196fb261532c456bc29801654e4a0ea5927b9495185412048cec8b709bf676b9b4c266b1481a71e1c55d02bc33028ba6219d9d7fb0ed633aa8f81fc7efd7716be0aa8b8727715cf0474c29e8a96a40e85168c6c3aa03badbb234d2d962048c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24bd5f0137770a00edf011ef6a641cee7721f50e211357bfd30d112e95f856a50cf41ffb32f8ba9fa9dfed7b79a9adb7a679e88643f0fbfc18cc2737c60aa80a1bc9875937d1204d6c25e0871183ccf58791b0ca599f83e7aff4ef6a44e0895fe62d36407427ac82e0fb0aa2e0db446ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bc0f17fd0a48796a39573bddd3df3259bedb4f4e832f2232c458c97f504f1f79f2c2bf5d387b7abd5df7b448a910981e57dcbfb7d2f1c960dc6bb90195865a07dc8b99ca23d6945ba86833e6e4efcd9907cb7684e1b06c19f36fe386dc4b3d32029030698837ee7cd7d93631c0834a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdd01b0afe36cdb43ffee0bec17f8b93cfa2050db9bd0b6293d946cd0b9ceff6a03813e6e823072488f8422654db27c10f369f9ff46f416e28a78a9207f6b8a38eabd8eeb08d37d26418481d61c6fc33d4d46c6376f3a928ede68db8ae0733602c6ef98ac5b8068d3101859bbb5cb4970;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfc52d87267dc0640fcbb30be7442b719106f56803d192bcf46b51abff9dc07c13fcd2ab3607a82f305a6efc29e0a40ca16f04700476c23b68dcd8a0a18c49fa8a648a2412eafa23740f58776eb49489a5a52ca6be7307f76e0411515b3d56c746c66621d842ce1f187ff34b1188252ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc680946cf4869d11a0887a05dbb58aaa52bae87af0bf03b7a4ff09984c937ce1aa3bf06f84e55723d6b6b992fed139e03098f5647c02cbd3e02f3f2d0c39af371d5d542be350eca878f1393ac6d1acfe2a8a67fa9b72823a4b40ab494c85ecc429bb7de17ecb90c93805103a09c7ee7d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd90c6882a9303ba40fef66c3d088c58b7f190637234987bdb43bd65c05d8e05374d477b3aa3f4d1044e3b7bbb44a1643eb06c945521727dbe2799bb45879d70be727bc1c474dafb3590a6176dcc8aae8a8147707bf2225b6dac2959d6cb400c8395db40a12a22f461ee2682d76effd40c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h324f5d07b9f9bf6db3a75c214863ced19a3664939fe7d5890ac22c40ec528392901d8d5ed5ce43dbfcba27a2f5cb0f9be8e0df59f8242c8021e7a779c92b996ed14c23c06d4075ac736e18767768b5f9678d66c2e3bbcff890beb8c7f995c109d412d9e93524049104aecf29899b480b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b3e06d3ca447c832d670fc5ea6dc3e6c6e965cb34e9864a20e092a07730247e4d95a908c1bd08c76457885d5d6ed62ad56099c0abf092016bd72b950812f7e162ba56cf4ad215e157ba9ac3cf527ebec25df50a842f75d82c39ab84303b432bbf19d5363a57e2a55340a076b4e24c8f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1447dbab1774fe1708b9cb1ba5e76a0a9b175810bd136bb45abe58d008aa12ddeb778c8f804a23cd963b4bc8208a1c5f8212bf8828bbb209368a79f5a93d2450b1c4083643062a4c969dfd7bc40b88dda171a4e96a84c27882d16101e88d3db86ffc46bec71d812ed7af10b44379e5def;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h564f6de3d74a5494d1f85e2fc89dd9ab65a3005523481acb3c6201dddc6fca4752787d38ec5c7f47eae3a102518a1e49930bdff6f16316145a947ecf84d82e822f352eca2510a72ea7ce9096ce315b6b5afa8c4fbb181794b6cf8a1d3b654dee07013ec066a03547ee14e6bd76d913f7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36c547a97c22601aba3dbab9411b4a8504a07ef850ed177d8e4c997b2b9d772c96289f8dd58df165a253e0f126bb38851127560d01a83cc77bb5e204769daeac2b9848d89b356bddc3d7405874be913a1de035bf767c439be7fcc02f1f35130b33ced4239e52cdd6e7f3f23a2e7d06012;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2560c4b001de2b6ca3013584def69e6f3a8129e0f798cfcbad636b3ab437dd0d62040ed0f3d2acf77645d7b4a900f9004b86a8cb181bfd61dfc4ff8caf7907bf7478b04969a061c8c5facb57b4fa8affc4f6e4fbd27b23527d562f31e01dd1064f6433f490851dcd6b82e2205d3279022;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d37711a1ae2b3deadd2edecebe94b3cf5d76fb60a7aaa23c1891b879ee4886f7be5c21937b98297e4cfed5dde174490a5e8ed23f1c9d579f7d68fd98029688fc2a7bec01838b21f908ef59b75eaf56a64910cbf3abceef29470b5226c842d28acb98922e775654a6b74cdba7d9297c2d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6238b185e0bd84c5ce86ed7b5e21bc89f1812711c6b14eb2d58a323b70d0141fc0d655e68860e7816b8709e7788f247fa5a6c49a77f0dcee3681a92b8d9afef8f5c35712119ef7d196573a7e7f2fc7cd04055b6b8718ba9f7c9ef40ee1861096906b1f5808393f2eeab4e29ca6902e0a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b55fe966944b3132ff8d05c0290ccf136527fa62c0bbe8a8b33ab9a75aae9b76c84678b83c8bea0710832e0cc8f2eba26316b438f31e2f8ab9b3904e727522c58513f3584109df417b82a73502f1862629a8e3f2efb7c3038a298697f66c4e97f5166d9adb76c906c49d834bf083aca9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he34e78c178582c46b9ee48a6718594ec4b2bd2960762cce93b5b273850b81a267733d9f0e33458798bba018939724208c3728111e7c2864f7ca923d945cd7e8ae627c9cdeb82eb86d019e1ddac941f1dd1b16fd1e815104e4ad683371f84fe030a6f6b24d73d57fffe79b92a375b6994a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d16cd3d58215a38c3c53c2edf679b2a283ffda7c5a1716987a380b991e99b64b5c932128310b21efc79a4271449c4b2ecca9be8a22381f8bd862e1b81e9ea222cc09077cc8fb4b463c9f071ac5e3249088b58c6cab8756f857d7d9804515e8985f5bf51459cda5aec4cddacbcd42b8a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h661cc69c899416c13355285d2067cd447c5764db678cad5d3a077d87eda08148d97e255ac095731a5b515a434cc9a7eff79f2829261f214ee6bd4680acda26d054aae8a3122a95dd1dbe7095c56e124914377e11171a27cba03857d444dae5a0c06fb52ecb3a043ed88a0b8d2118cd65a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4c64ae0ee8cdf940b53bce397a6b487000cb5f408fe826eb541ab421a029d7e358577b163d573fc13b3982bc311f90979cc677cbe0c7ef4694d19419c2858423e29cedbbad758f6ef191f53cc1892babd6e3ce18d0cb584e70d4f3a98da1653f9dc3dfcaf89ffd17dd155317f5c39bfe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h638253e342544867b12263d8b9973b2f6dc184a4e6c3251c08dd0f67dfd6188cb8e1753e41afb7c22470822ac608c4f754705f002269ec8560546f149e2129ba6b17f3258a88f30b2f070ba37c1e5d088a1378eb4c5a06022f40ed8808235dc9568d771eaad42fd8866892c5f36c28e45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6f1592a8e8ae45de9846ffc4c2015b3a74fad2e9070e58bfc77ae7040599465155bb61414d7791c0640d78b82c1cc29441303c98194aad7d9a707785459ee5e427921f7ef242dc1e2208f73c1a8ccb4a9c0c8050420ee56370fb862ab314f9246229c769685ce9ca86f6c9f24a33fd54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6f9bdf37867ad4d9e3d73457de5aa56e3aed86493c874d6015cdebd1c012fa8ff92192fd804619eac325f4665cf5e4d38c4cf7e09cbd7f7f2d0dfa4fd4c4eda27151c9dc11175983e267be6f6b420e2452f73052c816aa54502cf0abf69665ed60c499901a146885031e5b579a93ffc5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17de98e6b577549f5dae4612370097ed5bd473d7990c46d4b92036c08d288f63271c7049a5caf22e333ccefe3813a0f729c257f96e84bd72bd114d9b0d6654f2212542b77d7be2792a02b335d3a231683a681092b069bf7d0e65ba7c07fb10243438b886c058b7a9e9087b5455dba5152;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hadd9cb566a99a1b3481c6a9d4b5ebf1ff56e8bc1f6c23691c047c79ff0510aeacc8b22363f531782471f6fd642a4133d96532b97bc8f260ad10c28b96e3ec1ec0a15327be13816a8d97b109e420669cdec8f1bc9d8573f50f19d9138b3db3ab76426576571c3750bec15070db645f86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habdd4e9eb879ac4a6f4c762a05a8cbcf2bdfde8cf92a1a23ec42d78528fb4865e92114c84e926bec30fd390e10de08b390627d3d039567dc05bb47af0c3a44ba5f58967c1ffa3f3f7b5f505ae87f3fef2af9cef0f6fede70fc8c22005ab2dd377e2eb5fd6e3bbc44cd7f18d77c5a679fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7649298bb029e2cc323342f4234b59f393a2f22831d74786709a87f87b3e84643281ff36eabc9ba1886d53e12d128041d0153037a1e9be951b3b513a1e2ff7e7f7c2e326a3cd58d038c4021699a2bc77464b88afdafcdaa72184bf87dce50f36e889546e990bca9249f27d76297af9a3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7dd3192b5636d57cba89cda68a44361e8c7e51bb0a41b1b805f9c642184a7cea9008bd0ddf2b043659a6167a4ebb10afba1eff6561d7b6b6a9435ca996823c158d4c0d85cae9486e98a523bb9ba990385b694840142536e6f5db7e8213de0a199cc9e96e09ef30e76b3e6d05629f326f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bd43c69e0f5d9ed0b94f7c46cd244c14a43fff20267d25ddb337885a0ac354f62d4fbedca900d09d18eeb6601a3cd97093b257c9fc65a78cd1b1e44eca5b9ee9f1adae673d3c4449be00877d5b6acac3778ff4e866ea1018788be7ca965475c14f590609ab68e894d245f9cc4b967547;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81595905f6aee81c6e9a6a20f0120bca957a063886fb42da754a8798cf465b32809e28af2e7e9a3390197ae9364f606a695b2f122346cf50e4de85116781ab4e0ae6c0d4e0d3c24ac43824da883c1869f339bea2b13856c24a8151bd2f8f48497e552a2a986ac8b69e4705315464ebae3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2555cfd266c6966889fce0c59d190f397244d536085bdb4cbb810bb9c0c4c4a815969cfaa6af74e4b23c094c564977ee61d970ae33e928fbf04ea65270d0a2c72e557b6ae0b68b8963a9e8f180fc39c6270072b0e9fdd7efe0175fbdf9bbc4743d340b4b160c2ea81ba9208e52fe486e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6619b559842c8dd204a02c18ec425f7b4f8dd45e1dd8dc8e1f523937c38218ce93a0b0d81b6921cf6578b143fb3f3c4075be863fc96a7949fcac59883ae23ba64d6a26d5eb6927e2bf035cb49ec08e36e6fa38dca4392e9e52a50f777e0e1d6a02dcdb6cd1931fe69ca86bfe41535b5ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h354a4c4ca1973cd72687c31485e8eeedeb445ee9cb6aa128416290a47a309b3e39b9b00682acd57524dd540720adc9ae79a2b9bcc997b76a2a47ab8d293795dda96f3816b4b4b9101bd2e7c69ab8d9f9cdd7cfd5ab79a0e3bd9fe940d2dfdc7f41d4f1593bd5bf9186f872413c7195332;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2938b9962283049aed00198a0f49ebe957b26d7486e81b9e0ffe3fa7b451bf1485aa9255289eebd76c249db01ff2fb124974ce22a3909123851f3c770c69909575f59df717551f8a437e0b4225b5be60d2aaeec37e30ba5d4e666b4021cd7590496821261c2fedf9fb943fa9c28f8d0d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fcf64bead7d62e75b4121ad0ce852aaab23714ece6bc9b8ce586077d98a3a617bba214c58c8c88135abbb643018e92e7135d0e005bcf08542e524131fc2d949910000aa9667297156198282849bf64a5b82824daf2965f056f7b71a2c4a523fcd533dd744197f00842ae270246a4d2d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h255f6073c56485368b4c09297981b8a87947fc3def13782fdf1550836d3d2f27afab39aafcfbfe02162127c9dadf99b9fd0849c6452dc0afe7c13b4661b4babc7dd5b79b902f63af62ede1e2abe71d1f3cb17db149b09fa70a54deadd013c63be4c70f4dd65e66f9a531762135ba297cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6532a977159af5971d6358337013f8d671404637807939acd4ff96f1ed90c4717ec82ef3edefa6581a2ffc72b64ca027471d49dfd6ff9a9568f7feee7f16ea741946ffe2e08ae7f8ea89069c1e03dfbb34eee64494ffe92aec8cbf7262d680eeca88bcfb6b19df9e94613474fa5858b52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h474c8dcb48a5d5261bc88b50b445216993fb96ffa30f0fd9d3125c03d96c7ca85fb7d04e62b16c96835fb8a158a32e63ccd14aff167fa87daa032967837deec36ee1d48fae6b062f49102722030ba30a81f3f62980348a823ce0f62292c3cfbe1055c4737851128c03d7e25d45764fd4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64677a8b3392a5e587f669c7364f55f7a94a1209b645b19ec9b189e8794548e2ad1a7f176356c3b9177dd206f1401dabc9959bc0a8e446981309dd2e74ea54de14c7a0bdf0fedc21bd354185674a001317503ca1a04b493c8b7d09c4c6736cf7ba97bbacbbadcdfc8fb80cd990e09c504;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h330d970c00260fa4d7c642bc1aca6323ddd60cf00ca90c94b62e0585abf0b89c36e4455401245e6073b9a6bec0d3c88b0f30cc4b39fa7fd6d275c8a2e7f2626b6d62fc90dacb27d7be1dd9208c49d9ad9113703286195437f908c73c03ff8ce750e424bbf4604f86521eb511a49e3990e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h568f53acab11c1e69bb2004661324eb0ac42fd75c46a60d175982cd3f3a2d0129dbf03f20aca4a53331c59d3eeba3e3e6a59e1e94d8366c0bee46aefc110666d59fc71ed4e516c4266eccdb9f0c546b82f891efbb64f498001b076a06c4f5725dbb9edc6c4a7d4504abc54d175e2088e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9526df14cacaa7522a069e2e91ce29e891a50567a654abde327406c2bb15e570e0b04f6518ebc262171f870fcdca0de86dafaf2177cb6cd914e2cef907302b7c920586ca119c9af8f9167628ab2ff722cd39736d6cf0afcc8576344d63206d397badffab59cc0450a290cf8b23cd2962a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50c0d0ed5bf8906b1206563283444da3b6f0e495152a4a297747e784f705f8beae4010d051a60340031b55d2a685ade758202802811392d8e436b2c497318c3068a254ce9048a052d979cd16c1a5fb88e1f96845a19379cb2e0fee1c090c36c9a342fdf43dcf6651a95162250261a8b31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91f7568753e1c0714796c2c4cfeb82bbfeeff6aa3c190e0e401f0a326014b8783cdb3145cc248d07ea6c04f04841daed0b80c2aea3084d76ff686814ec0e92d534ff5115c004aacdac252360cec75c90f9ecf2dc54a481914d909cbd65c363bc407d5b6cf0a8e94adbc18865b2bb227b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he773daf746c9f1cd5070ef98f4ee4fc6be855e786341cc84e2b215133780354f9e07088caef540cd2aa139b8aa4ad7be17bbc1d7dbcfe5350ff2693997c3fbb9aa2fab91ff44f774d10f923e666a09b25c445f99e65c156c25211327d6e9769c1251aeb215ef1a25784962670d880d645;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5167a91e8748b9fe767b41e30a817d22deb966e2e0446e6f0ab7c3b43f94f0a1b5f40c48d7816cd9283c37409f343d742f8e2d4c65ca591e6240f1f9037d1dd66d52ad746a2601f45a367788fd3907d6cd67b2f831639a752f3d3e6ab7200a36da47835dffcc99cf1a90ed3bd553b22d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cb9ff26858b5106baa89091c29e29f8f18a2eade2770720c6cc636cf5cb63effdeb06c3f9787b8496de266289fc56522a7984745778071ac9ed76c767f0d4b021c7022350e0393e37970ee6696eeb6a9cbe48fce8d2769dd8676eed31301b7ed0b4530e52beb4ef042e32177b032a824;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd4264ddd13af5fc1011952c036692df6510743ceb70cab69bc26f0dfb91372fd131e51fb81e5b0bf3daa4329d672004c3efdc46c480bbb763e078798fcec44d43f6b7f2b4d15402e5c6203b30f207332c3b57dc00a73fc9219dc94c7f69e2eb5624bcb67adb84e5575edfbd746dbfbb3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eb9da9a770212b66f349dd55ca21e7c72dd230658087595a33ddfbce43abfa154642feb78a9cc4322f60911c70ff0e6a6b345464d1002f4164be4bee2bec56a18fc4d1d649d39048ca9340b927faef5814637f0c406c2d42db115f613420960cf4ef87fdc8f1f6005291d278b804d73a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd7b30ca91a01f833816b3c526974d0c1e3a8a547f810a504e787df97eb08e6cd8e49069d1ea20f9f42b65560486732b791528f62ac181feac957377b6d6a53d3cddeacd1154d8189fe464e24bcae37c65b39261a2db5b4b76505015f0363be810a4fa4c0ac354b4ef7dbf3f8a4b1fc0c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde067bf54db8502f331f81481e4381e29f4845dbf198655dc90951979b3f9ebf7e715c07b1452e6477ddf2fbb30f99fbf8aff270167657bbda05cd369f19549e7f0af5230f2b154a417b76265a46cf515dfc9ee2054bea78a232601bb784b4b1a99ae422f43419e07739e37f79c12c8ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h555b77ad5587ca13cc40d1c1c682751176abf61d271e4d3e12812955f9087f7f90dd09ee11d5f47530c3a9d621bb1a51c664154702f59c0a31fd509f53f303c3f6aa367f88b5bca1db6a6aafc6e9c2bf3d08adf7a617222a20a11f4fa1e8ffa3486bd30e39ebf23e41ec24df59ad6f2a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcfa4ffe977a1f72cf92448b2f044af53d7829b21583284c08c81a503ea8bd4e61b8bf03074cb7fddde10934c1a2c0829fa928793a0c70431c210717e31afb576540a2365318e43611d11d4d6b3fcfe3a6d96af35bda1bb9a2dac3e302052a138e74bb2e0cfa18335ed483450a6c3aa77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2fd6483876a6f10450be59c9238db2f3f29ccf0bb9d9cf09ce6af67e4edb8c48680533fcc28faa99815f6e8cc4c434207b1a112f6c0a1c19d69a2254827ba68b8e3cb1eef00d41ec59a75839a9c44a08b950ebb24449f6499f8c22691f2954dea6b2c02dc04f52596c5d80178c83d032;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h468ee91feca392925b7551de9e5d51bec2ef25946cc699a522483312ddc332a05a9903c7c94901c26df299d53ff270246a4705d9622ddbd92e4e975fec438031c8e73a0c3e6cae92dea33439e2b4e1e6a18ca119932eef786ceea7e09e320b3fbe725ffe9d9fb4f2bb527bc2384a556e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f808c3524c612a1bada1bad1fb12ee0d7367fbb826c16c9174d1c58486dcbfbd4e769e66f06a1e488503e2e8ee769676346804c8f3bde6192c932af836436097e1237bd1a0e269492f9c36ced129e2cadc07526d8b9fec56e56e92677028f554aa9027bc8d86c4135db77762ea1f61e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20bfbe5fd556a0123f0b3ace28bcabcc15937936f9d2cee7dc231d0342267f0ce824150e6033da55cb488f9c73e1daeded417e9fec178fee3e701c9d4780464d3918cfebcf76c7f88bdbe10cfa24b681c432dca1691ecb102402fbb42b121d39a2f245a7596262557a1c75ddc9938dc32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he90d25a27b91724b85c6862cc57adb3941e48148a1d1489b2892ebfd1d99093ce99cd1f19d79042aa9a550d70c5ba6a92cf772686c6ea208383c90095b67ad697d7a11883b07e7dcfd8bdf9753d175933ac3817c6e9625b5182cfbf1d5cdec80fe0074a652dad679592ae95d97dd1c558;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3f19237fc9aa8ba5537543571245625225446840406c2b44d4cfcc4061651e2fb2d6b8f5b83da68b4c2c8bd33a6a993707dd145229943e52be90c6e1ef29e0eb188000e6ba8b657a3af91d3e87bc06f0df400d36735269f07afd6e6df842fac2fd6d636a34cdac9c6ab955ceb922d1c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbff98198a10f6195f40b9f03560f86bccfb40cf7555b58714a07f0b641f7cb4be6e7fc4d7ee1f85228afea233996d68ab28244fa13a5c26614b7a7300862e79474b1e88bb60625579b14c9fc3637cddc6e89afd3735ba4fd282b35dabea2808c1a0d5818da7f9228d63d9e4999e767073;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf55772165972ef8141334341125c44b45277a59ae67dac8e0899781c4daeab92359f11c3e2d5e8066085292f6fb593c8c80e93e14cafc34fa9758bdabf19d9f947fb5123e9a0a0f82d67fdcc56e9bbd65317180d238a7971d066aa650d3212a44e0edd5611ddd063db96bbb8f6dcae7e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h946fbe2dd581115299ef3c128e834dd1398a889c1504d1f84d7b9a7406f32ec15f341c0e3c7d8db2bdab80718bd1f693058542171998d322fe89430c41de55d71b7274215cd0a5eda935bb00e3d73820181ce8d09d4e1e17df97f42d89dc1d1431d7aa7d43a3bc2c9e87548c66d594a37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c9dd170945afd3ed41e84584d4701e9c2ee9af6db4980a5a945c494d57372e6e8290e25132a7b7ae4dff3da07bf4abed5b79080e2021daeef5c0662dafe74c6d89987ea3e7a2152c58c0de283f7785c75fe7bbf560337bda8682131699321f36c1f1e3e42e77fef00c46264db28b362c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47d5b9d248d7038d8efa12cd809c0f0d00d5a0d24b1baceb85249e9fed2782057418408a2673ad477d4419e398e903ccd9f03dfb64c237cd11300c2d419c4e5496a10fc3a7b16355e83f5cba6dcd7fb64fc1118f59bf6b15a7f2878213e2aae83310bac4e77b36bd18983bd0153b912fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6083c7e011df0a9db0b20de65a6f7b77f809ded4cdb22304fe7d2a293230b927108ec0f056657ea8ac0d0d3d8a5398e81b47060dcc6f0d14f3c50d774ed2085f726eec2e7a73ff8aaa6485211c2bb211a54eb580d771b1d305e07f4dd164ba903dab0dcf085c984e989f8ee60f1b1a536;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fb3510750e0d4dc95981d5eec901810be5e3def94b5a3345abce67d9dfac95d78030a070fe4b30c16b33f835afd7b52a5910d119ba50f51fa14b5c60c4ae1b155aec1f9fd74e31c9cd4ea87ef02815c981579fea8b5a3af7c057f809663c9b502f7929a8a116bbc5f5b91483197799d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd41ff549a50a961bfbf8eb990e37c184883acfdc8cf5adf9f25b9aa335a774365e618b444af57bc78dd3593a37a83a078824f6841b95f165b258c02b5c5c6290bf6ac50aec8b76ee092bc8dcf7890998065fcbeaa9ad2ac7c7c335da00dc637a1be35e9751e971d7c6e9a14dbec61327e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8f5d06ee3c68d868fb69f78916c149153ce6fb2577071bfeebd6a91d2163e0d65b0cc80908ec4fcd9a27c6ba3b1460cb8aea6aae5c77bc8f6cbdd9a1ca0618fb401ce345b11f77b43937e41242c1458cbcd26aa2c6e397b87b66c76d633a84c656612b8e105ab57e6f197a5c7d351b2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h647f838c640d3dfc79bc84e29c73b8596ddcb1dcf37a585fc36c0811e3ffb79b09a65b63d4463a859f4d39351a68988d692d1581683afa77414248321c60239c466c0f164580cb76a90b0002c08bb445b3425270faa8db937139294b3ee7de2185b3160332b5edbc3b4af4783c85907da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30bf4b911a68de1938dfedb59bbe081caaa9151d0bedd5da144404c068b201300551a5d31131373d37d99eb9577572b95e60d722bd97537c7ef8ff2961d361f2db043f71b21e5d7b2b1f68fcc13d4508890db6a2114b7dd0be777212db26bdd6109d4b3da7c968ff9c29288d2ad9e7dd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h791801f9226f31a8c5794b77e5a9b0a29a6060e34196154cb5ec982f3ee47eae927e584b8513c019ec32ff789670ed0fffdcabb3fe6d5bb54b1824905c40fe2c0164f4e9d48a37743583fbbbd7f2f371db4ebacbaddda5fc63171f53e49f215f19dc456b1ecd3e9e0e71096e0f7ef9d1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5975db506192d51f6dfee2fefe9d1a3047aa80b899ee1273f907242cd205720bdfb4a64c990fa4e956e53770401b625b80743be5ab5f6b7494db9528832203b274da29bcc1f5063a893d3aa682ef78a7a87b8c5c6a0274c19a7fc69902f5ed245004211bd35a1d98fdb77cdb0e3715d84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb982a328b444707e33bb758dbc323d361c4836d9020ad0453322669eda872b2afb17877734a717b4834e8ce2ea92da0d00c530bd3e66ad376862ec5ab0feb631f5d3afb4d8a801169d49b890f16931b496a589d205589d7fb71035235ef14dbf0902a08581b2ce07fa0ffeb55ccfd5d05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd54872ff1edfe706a6b543f019cce22ae2205f3d5ee00f5236c934382659576b51fa37a5c87c1f82bef20abb4cf8027679f1054d5dc7b4485e7b29b3953c253cba45c2323975a8e5320b5cbfa9e4e4ac06af9d656aae775b1c94dc2e90545e6aeeaa4609de1f8816bdb56db62f2e6c1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c8d5723ac30ed33fb4dace7f8493c33cc8bf1172a20466212e3f9adf58a6a7192ec17fd77461349a12c231fa825b8cce1cff901a7ceefbb88d87bde7b0164ae707abde8b7eccad0d55a56e449f3571770a79fceb9e2b372ed99c0e6abeb226c2d3073d5509ea6ec7cf29edcda524216a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10d33baf5a53b569edb245b03fdcccd5b61038ecd112fe31965c75528859525862c9f9ee2d46cebee2c5b4b6294615707ba96ab9e98bd5d0a4184b1000823f70b46269dfcf4112391e29d94f9e43a26571a48088b3d75184e2fd38f7209bb0c01b758b0885849c8795849e294c9fa5e37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16c3287061df705502c171a03c11b727c153b3b8cddddcd0850abd01cfbf78d447db8e273f6ce8f720c95dc7a29531ce3e0767b82ae530a1272e1c43bc6ba779d1280f003e83e6808ecba8fc0b30393d94c4e00dbd4554b859ea66d6ed46e9f394cdc5bcf5b5d3745e2071b83d6c55b28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h166f3654c15a29bc61cb306440945c8ae71c97e704d0784b19309bcc70d4bcc1cb735df88b49add8889c5f3f04ab1376a09249d11d292e9b73d0351f5866f577d9a3f16d01ad2ee41486328a5201f5b034f616ac9c2da9abff2be588b9a86d40799571bd120a86ead1a66a9487fe131b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h271e9763e9eed86d0965cb602a0d0f3d3ad02846924a9dfefb5b35fc24e1588c17a501bc3c97b0144e18679796b45dfd25231528efec292edbecd16ba1d20c88149435d8b06e5a8d77af9972fe75f998fe84c38e3cec03e29c7a9838205321a6e362a5f10d1cea04b4b7bfd09011958e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15de9fa4fe164f68fd91495019c8d2105b10653fb7677e6ba2eb4ee8d35fab85c56301b8385f59e35f4bd94e6c348c03090c4979e2eced2aef43d96d2e64f884ffd57d751571801945bc370bd40960cabc8f32b3751d8e087841b0a84fe5596b770f9cdf284e08cd6af8dfb8d37bb46df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4524f8a1cf497ff9564e1416ec680b9d246ee08ed138c8b062fac0f054a1521270ae59b75e35f7991561feb255975457047ac44b95c6b79c4751accbdbf9e7e87cd9635a44281a3060ad3886f4c987182831cf8edbb9c804cd4ce070228db7a5c34ac3fcea34ebddb402fff7e9b9433ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e63aeb49647bc5baed49639160d6e09af193a468ab6cf4f168e7c89f72afcd8f60ead67b5f6c0febad332d0ccfdbb56c4409eff89643ddebd0dbfeead64c24aca0c75f3f6a4e2799cc32fd34a05a432b0e8aef068fd06c92d7985c95af0c19b619058dc98648c52062d9728490f167de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88c356a81b0aa0c9b5b6fbe75ef4807e1474d48f3bc0ea710cd654e935a10d9a71706b70f5d81294b7a17715fad86940765965f500bd15a9b5814dc1f996552e1487e6d2518920ac952828a6e1420c1c3de044d4436127270b33c6259df0d50a0a2b7b20801a32147fc2e85733062ae7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd5a465d431ff322e86cc50c1aa4b448acf63b125fc180ae9e3ccb044eb46e42f684653985df05147bf312f154d35dbb9b6cb294b579044e1cd668af51bd6a1fa2ca77f504a99eb65c6db5adf92803c53fe616213f25cf15bbc5420a1df93ea6d3e3423c05a9b0c0c3a88b777476038ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39fa4e510dc41d6fb6847863e0d5bab4fba1b7fb12e8737fc9856d9cfad97a7f738c0db6d32ab6b64c32cf81d4989958fec2abf15f8bdf7caecd30698438e494d229f8f7c5b7cebf810c89df23184855371f8da163d8cfa2e0741febc728b9e02b1c1fe78db5c50b846d48fb0b1a32ed0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75272c159860e47829a06794611c0bf0373d5e7c6beb18687c7de1b5606afb62173e60795799d389c0eafc6ae7436cd1742ca1a55f80a236e7f62e409e5c9452572cc44c1ff007f34495007a79322ee84d05cdc9f1002f9c4f26f11793ba94b453c6425fa02026256c15aa43b72d7dd23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6390ea0e41d9277de2a6f702cfa06bbefe7b32a09d511c1ff85a84c414fe26990a78a9c0535536388b1db461faab000427672bcca1b4d2fda9f85daecdae2631240d2c6671bdadcc909830bfc3c2712efc0a89d79672c9b72fa04538f9ec08f404b0b47107d7eed2226a821668d31b15c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc516dcb35175b781cd7bf180a894e17ac8097839383ba2304c447c2020a039089c692759c76b102e45439284a1a5ae287d2609ad2c899254449500c26304ecf56457a7d072bf31310d5a9321e4d06233de15ea83e28a370acca295dfe904a25c1ae36f963b315dbfc2d031820849c6f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2a786b8c1fb3d7790f40b1ad2117bc647a4c6d5379aa0a8d151476131e7b8bff7cb3e94fb18e75c062a70a988374ded7f339498e5a12427991a3f4ecb8838c3bffb2e11589bb789ddf0509b835bd574119013c00b0c05b360a6a175ec076cb3f38084c72c97a68d053d61f2d30a787e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he09e27d7c97b0ead4f74a5cbd131fdbf8c9d41f40330cf901e9518933dc68dbe316a3760ae1e134fe281ca7d65c5fc44bab856a365e263f4234b6f9fad63ac7eb6962108621257e47a4abc79b44584075ba0cad20e27206aea35a17e05c38a24510b9a237bad95e2fd206f712f9a10dc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53d71e689dc42b46297434f457cb955509b53b039eae849365180b348037fed033848f731b2fdff569814f7a267a2b8a6ee9b0fa8bb93ffa58cb0f7285ca60e7b86577901460fc84d277d48ab75b25f435a65df042374934a2b19a5f8bdcb6c3af0c4d737e13effb06fc6e9d3dc8fd457;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80bc09f901ecda171f577f375a0587f9647b14dd0a071fb36d7b661aeb4a3ef9fe0d85c24307672117f82fa81140643a5c399dedfb15607819a953545f6dd212b5175ad23ab935d798aea5bbcc24b4e61831a532e90be62d911699cc6b80cef385ce080d6e8a7f94fc2ade970949758ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had3dbe2a504e1dbe63d6372257a843449499cfa0eb6555e9fed9887b32ee7ae4261e262626a86b861feed92c78ac98e4ae75f07eb628ea448cc59a7f39d47456b0f8283473f74d8a27ce95388744d7a891ef9ab1bbf2d2f866760491e01a35a7e950ca902e45e554fe33315cdb36b6ea0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde27b6bcc639069d9ed880fc72c114d60765ac4deccd912189a1e1d78f4751949056ead778f3ca0416bc3c7a1b5ee16c01d10662ec23c0316c05acfb480c0d79a212540b29b29c4693fea793e6f7352a40b1df60c4f887fafbaa70005961c2774aca71962afe09da41ce0fb17bab69e7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9712f438937a85c49662798b6f4fa1435fbbff243706ad644f1ca01a33e9ab353e63dfa51d222b71d1a05dd87659de9ef715108c63521823def30313b58f960c137a3ab8279dccbd41e185c117b34c275d6e54a09535ffcc78fa5f20ab1a93574b22ff9dab48b8edaf3dcd19c62b2bd47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba95f5d26ddb5c64c38ed84d5aa1e2e67d44a220f51c8385791004937aff183c6bc3bdae3ec97d60534e959d06a3f187293a315d7a4be80051208157d7b250aa8e15b8500f06020886ffe2d2e490422d5865f580ced1878fe586dc08404b8fdf4d728c030c4803bd06bc3521d36c8799f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a6852ecae2e6dcbca31f201290fe704d8bd0c00cdfb734e55961dda250f19c403cbf1c4d0fb541b0536ee2a7e514120bf655665932a38cd04e2ea5cd76df5a4e4f801bb9f3c78866ced83e38e36391abbb0714726d4f9503f60fff30b731f5e2dff7a5107a6e62d3a2391043f37dc24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebe800faf2f49c31054bfa7fe407ea5bdb964969472743f7770c3f90f336d6ca95d628f7b5190498e801c2760e73e7573d9d2a5d9ee36258984aa1d6779dcefc627112b15367c80db6ad1106811d40e211aafc0e2346b6741ff303f20faaca559274c50feb26711de54222ed010918933;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6edc5fc30754993172e88b69e3065b7342a62b84f0beabed17acae455e5f4b837135595729265f0874fe99987d5e81f64df27da53e359d2b891ba0ca79c41f76daf3a7fa84a21d2f5da0ca999dd72b476349c750e4710393f458494520e74e8ebfe3c0ecd9ad9edec742ad333d210025c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23f67e73ae770f34876a88e586abb5050b944cc9b1232e1ac1bd3404e126fd1cd4575c95a3f320ac1617b41a8bcd9fc95675a0cf2d711cb77ae4121958e57974229b3109263250b3b053ea6ce98bd7b6ceb375b37e649362d9d2b84b59a54d350ee3642bb1a592b07d64f07b23a656a2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7eb6b847df22a66c7b1526214d0ff6a5a510fe57bf70486f71b61848404fe08162349b517fffb20d7b5a5e958827865540014ad05a132ed6fd505b2f469e3b0ed96916dbd4d900732d824a8f07968543c102759eb3f09dad25c98474711afd66172098c6e132639d52bbacfbb90009594;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9834e3472001ab261d16d42dde01e9bb00475bc68fd2d00e525071cc7ddb8c0b3076252c512dd9bbf9286b7e128626e8e8e64000fad839b932425adf27bf9be5d1bcb0bb6fdb3bf77e733b2e129db6b1133b70ae43f097fd0f79a26b8d5b2764bd4e82f313e22fc3d71817549db683e48;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdd15c70b2d5752647217a039c818e99e70fb8f85b44c6b08b7fc9d1740955903961fc5b4c565ddd8dd18f0dc272310f3fc7ab4a9d1593033bf8764b4352ec46366b661f5b54bd73c808e2a1bd25f8bf77c1b238ddbec1f8ec24c4fcb6a0e308d479718c38fd9afab50a9608cb4bd641e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb66b2077e46525689cec1af12c55f924689dcc0484ea38ef62d36d2d68e8fa78fc3dc6898981167647b8ebdc4122a6875aec23d4b1c327e480d4589e20abdfe1ebc36ba6e7a834b2fbfa785a6c6ab3cd820f0b3e9d31ebd86fd850eafa0a3d83139bf94e62423837101a071cb6d90701c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb162630e481473235f025d0083a7511ad1d9c54296cc63bc7605439b3f64969a17a779b0af94ac6f72c1d0e51e24293a95ea69f073f074c2f6bf58097093effa21c0a7fc78c1bd5d310972546238b606829d5efe9186d1332e540b25d14d2c4c8be16e849a7e683abb326e014caaf1ada;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42630a4d704c0ab854cac2f9817c8ba10f78c28d050996ab6a06f1c887dba7b100ee47466abc0e7b346ea596bf2dd72bee4921a090c207a928b79def17a08694c5e1b72b837b7e353e264ba3bfb9cd73aa4bbe0f8ca4fa088ddcece98e6ef030eed710c4ee477902e4f396882046dcf9a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1d8e1d8bb036b29a86eb85f5c1621926d73eccf0f51ddd28baf981f6a2b96a63ca97d044ad9a567f190267f7327867962defc60f17b554075c49d33dd783e3400f679b9ed80857751e9e7fdb48486e65cc4d6f2e0036de247de12a2b9bbf3c8b3758d612245dccd363416438c38063a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha83e7351cfdf15862a1b66b70c7c1eca48d13075630183ae2aa087cf4281205d9720c4e58e7f85834896647678caefe9a0ed5dd84a4c9474c6a34ffb4640b837d44fe8f27ea2e11908ea6807681bd1a868ab968183561574c9b44daadb432c9e497152611c173107fe9c50cdd21374579;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9477045dbe6a0b8befe7ae598708b5724c059bfb8ab915c6b441bf025f4a8f608987f0ec594e604f09af58f003fca81a85fb7075f19397dd32abb2a105ab4c6b133bbcf9145153a91114dc394540d0b4d82b9e3e6f9e6878e1ad51d72902f74c68cd8c312c396d7e0b6495a34467d1bb3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c02508f020288e50e828f77072959bd564322a6692aee418e9b264451b82505dbc07002f8d703f8879f027704d3c185cbe381af23d053cfe58d8ab12a44c19d4c9227d9cab3efae347ac093062260bd82b2d55e61280f570ca86a2426ddbe563f5730ae8a7a4bf0b61a581a77dd0bcf7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28df5f695f2b0204ba0fd227ed0d77ab28ad436093dfb51f603164c8211c9a7cd9134c9f2fabf75c8c1379ab3ee4b5edaa5d8c4a406e8f47628397e2a6e0711403d0e2036fd9e180051d18c38c2df72edaa57af27c83b3f31caf97d663fb2e5fcfd16725e0d29fef6a7f4e4000c8591f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78e8dfedcede6300852e00fe39507e4ba2c99d34d7304e6e5807bd25901b201efc0ec16bec81d5c2362804144a031abce34ac3e772a0f6cd3887f60c72037ea61298b8cad1321aa26975aca8da032c248aeeb249acb7be0b6ebac68c02665efc315ee41e820cf85b9b35520fc5609445e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f3c9ff82f574c291d272ff668330da4f892e566f1edbea64098ae05bf0f4da26beca27d6869d37527c4f952ae1229530a1c928d47f861d334dbeee40b12e9f511acc7da223d6cf129591276dec860a5093106811aefb568b0d4df96899b0502267408cfa2bedac5befd3a43add8e7e28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64a9b7e7c3a219205709dbcd644ad4726fe8b9a5bde5ea3f5fdc6cf6f27ec778cd313f8784ced5b8583839bcb82846ba37dae448288c78fd159416d2757f440d1c85b5063de9cd0cf9bcfbe873241a9ec1119f68cf43b895681ebb0fec6928e58c257058a6c85f48baa7eac398ffe9245;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7fb5d6c7b552b336360516bffc464cdfcfb6f4feb001dd8a07f4f1aa69f86b8d5d081d5482b58edd12173cba5c367dbe5d489d3bee52e13a374232704bcf53d8b5c67567e04788e6ad981144e6e5403a6bd3b097ef5f0d03bf4a5fdfc5a550a0d52e87aa4ffcbf796c6ac331c267ff53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7215f038499d8bcf8d6aee45c3e02aa23adb2bff7f9d42be148d74349d404d6f9f9eb18868600631bcc27bea93b2a423872d9846ca7ef794cc9da4e2fe302b6eefd564d80fdb1e031eadf174955e64327c8f7ab0c923eeb0dae116bd9b4cd71aba2242b9cc7eff45abcdabd58890d32b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h365a445da9832a7fd66a7615f87368381a21269cfb881fc2f189905fd55d53acee323c51d1ffbd69004c6e3581edc0c8c29127bd678a58459a516ecaa3bf9f72af4b5fa697b826ceefba0c39fdae85951e8356b1d8370af2c4565376c25afc604fce610eaf2b81e0891e68b7bf70b630e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h891471ed8970400403e33670434bdfb805c5b121b0dc009c59f29268b269a7a776a1cdb4557d077534bf527565b2bc3e655db59a6740fc38e00e46b7092e8956ae586d2d779642d67a09d9f3d8335813d0407fc7d53169290243805ff41a3d2df9e9eee66fdb99ea11b8e85206f57231a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha863f034f087d81d6e4b0a8f8915cff0aa56da59b99fb1bb3cec83cbb05def784257b5ea534665a10c46acad033ae91acc0e878268d2cce5d1c5ba919c30abe42ff831028bd707375c166296f85d566f23c5963c62e9d2ae2db2f00e509f96a1ec5db3de75090696c185fdc5643c20d2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11e12e17f71a0125096015834de4ff9036f89a7bcf7f3c8a560c3f1658d84b551b3b8732aa6555285db1a10e9435430fbb7b2eac98be254f6ef0faba1ae31d4e98355d4d98e3ff3c41b17d2e262e8d55de6b3d30194956ed689898644e73196010636f4c8d96b1f2dc90b76f596ea9624;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ee9969eeaebf237d65cc5223649075b8b91b154c26049065ae6f7d7965e4d838a78e35e8b0fd84af4b4b0b252545ad4d6abb7f78252d2c658632f2c08656414b825ba2172526aaed2061492d97350fb19c6bfa53c5dddd95371818e6efc287b47625525a82f4804755def26b9e296cc5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hada9fc27669da96f1eac0e5aeed3a2b9b05c5965e455a316c0d237743fe6e846448a19874c48d44f94958588c029a43638d527d31693809d9a3672693951a12757855ea205957e50518dbbe23f04075b8e0c1262c69bf17c90e327ab686f4ba938e62fd878f8fe430503c82f61cb2620c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cba66306d0e54d6df457ea17b051e993e46883b32d973fbe7e690ebe33a08adcc7863f82e0a7f2b058b0408063fac593d483a9353d8bc8065921ab4f9b29a5cea3dcc12e15dd0f523eff542e36c0cb01b2257f03dae614078cd6184abf4d199a17a20e8a998456eb96101b3da689f950;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e33a1122988b05d3f0a13150ac08b8cf7b348f08e93f135de4311fcd18993872a33721b6f478a6a09a69aae85fe5ac192b6960d235b2b15ebd288e8012ee1b80d0c3a488f4fcd735710c839d7f2d6f2e2a137bd7e605e980bdce95469e4ae44a7c10ed8898a3ee33e4ffe9f720c67ad4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf802fd533074671b53ce1475e74df794396ee150e5b5b6fc999de678250a427a2a872ff82200e464a6da8b30412c965ebfd263da90e21cdb2f85107e76c25829220af3059ef879c1927dd1332055ed5534d97c9db49e165c62b2dca74d6ef5a11b9d845641f0908d4e9f5cf785e3fb22d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9b0ac4d02f183fbc94fced0946474d754cd951bd69a545fd08e948a14ee82562a96a1ed5486d137abf712d6e0a14f6805fa90cd68504bb2a27b6477d39b9e3a45154216d91851a013f5f18b86026bfe3e1ab1678ee938ae295462076ae5ce5751d41bdad8156c10caafb5a8542fb27d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1af6811a4c27dbd35ac84c50b9a0e863edcecdd084880ae2c86f33328afb098749a23015a7a5f8037ae052197b9cb5872d962cabbd89b5dbfc097a6bbf25d7249f07ac79f1cda0c27fbbfe0297401be70ea0d92c6e2a344b17821998e9df9ee6bf88b65ffb1b5fad57a358a8b19140bb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbe0fdc369670f2498e2c412ad79b8fd146e8ef821d8bb4bd642ff0e18333bdebfc834a64da1216d451e1dd7a1d54134dcfaed50f625664df9a4dcd827d747ff66606ea2cec614b9829e76730ec9a3a6a0b892f30c4c4fe5b9b313418313598ba6cd62f385eb77b3b99af2659fb1983db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bb894370b35ff44dd4715c80116a5461515eab501335bc33f66edccde28bc8610677fb9ac72cf1bc97471df3f8f9619ea826eb89580dc4cede76b48ca0f9afbb55da71951201adaedc42ea651e3cf405c6f6dd7313bdcdc1e544ebc1c5b7c482f2bcdf93e6acc4f10c9d3b60c17b2685;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h166d8359892d40b3607f9ba07a4ef6a6f11beb547b7ab1c52728c7f6694e1674d5f4b31d1c073dc39cc0d80c171b0f29fe707466b8f6f5e985c1d83efe139fb3ce3b7157c19eae9eff3b875c3a1b56d73f682726c52b82b97d905598083937d980fd93611a5f2a53fd8c95382e485e104;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e513b88e153ab8b4e990f8fda0eb27daf5fb95f59921bc4506409d7cead09c634f78c9f039daa0b407c63bc74664bdf660bd3ca5db547d2db359a61dd1cf903c8d71958fd962645368f3fe510b99124076487fcafa56b18cc3b14db2a7da16f543ee61cad43abc632eb065514fd8e864;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff01a2abd77095cbbf28e743501c9133e6c22b15761c76e7c4d509548862e35e02a41deb829baa385488aafdc0c3d008c2669580f45dbe5b76b5e42666ea38bb955584e111ee8d5d9ae28e14f5147a67013e209fb671f8180ff9b97291f4c5b303242dea765cfd71c098d926ebe4fcd54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7e07a360f18207c733559cf78970c423286ca9df22ade46a45851b6eb5a4bf755093fcf23f98d7c4ee72a648eaf68342557738be792074872a25bdf68fcf62eb285aabc4e95b58e428efcdbec426050e078cc231e4b6e1a46e29865302943bde2f11941d2459d2037de63e88c1c623b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3b89af623609021d5fbc575deab8cc90ef279c46aaff39a2d18132bc9b5ab15fa84ab2d528b2e8eb3d86e07297717a2b7299f148bbeb34b6d9d635da9dc39fa97555cc939882242677ba0929cb03170270fc19734dce99415eb0c4b051506eb70b0f6353a4e281a76972fca8ad3a1cad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62244f3b4cb9f01a1fc644cf70b94cfa21d459fed31879161bd26b35627bbf2aeb85842c1d45f49dd8ab52b4f5cd36b221ad2854ba76d03781612d6828d1376cf402d6231809ad7769e6a7a63bc6dbb364f9239476028fa7a5c8c02309c049d8eb0adc505ac83a6e67f2a5c0d505eb6d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36ec209d3544cf6c68d3959f8cf44f55928e5e158b96be56e2e6fdedc8f6b5a93482377a6e2092da2f8ce4ae1f9ba031c397f6037696443764beea138f32c6a407c091bf630eeb29318fd894ec7c8a44c421db26707beb69e910b5c055a81a16bf3dc6caebdd0b88b1979da31c60c4518;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h397cad0394c5c666b5118c4e31b384c0fd88aad1ff774900fa9453d8bf352e7dd5017cf33af7dec7a6d2949320a7bf09c2e9b37cf1191ccfe55539b6d8d416d229f0e9e304baf4f8e21edfaeafca45520f01b265af471d108a57e4cc2e9fc6739e665eb20face05e03ed26012abe4ea3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39e7a45461e7c2965054b6473db6d53413194770ec2537249720661e6e6f520bc3402802cdd971e19ae0a077da7822703e91d3c8607370b681ebf233cd2d91ffe96536810c05ca0473a451e2d566062b4b63a6090a19f2146bb61156f891bea8ccfa3108b0fac58c708d61e50319d7d87;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h504dc383121572027d7e9e908c11ebf266b72e85ea655d516695042ce3b2fe67a1c78592997540a20c63bbb8f7b81d9b9ecff31828c08b4950676d88a894e2b0ee6283e802975237e30ef7b868c957cb31defd8bfc3e1ee88d4c12ae5db18591fbd4f8967a04857738ac2ae8961ef6bd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee9abe3df8a260d50ecac474c73c77d95255c3a6b8e0b1a45c07bd7cc93228c33789e19ae5e882fa8b017bd4953f2fc42714f6ab985d9b0a4677a2cbf256b00c1a17c7af7bc88516f6631f11821e035ea8a850e889e2e723ad046b09b3eca3c936dccc8a6abe1e171b7f1e5c8c1493fc6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ffa3a60e4ff24c11a0b200427a2ad1ab821473f5aa1695ca0bc2c528ba541efedbd709d8ba47d575229f1bf9f87cfc02e43ea76ed9abd4957681001c9bc46f22ddc91becdac9557f84670105aa80dab65c7ad010a7f7c646c9ee31c95b8a62c9b3c8e9766f1e4642ab41994fefd067cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd069595e871a66c01874a1fab1df0c94ddfda71f2e3ad04ef9aae2be08907bb120c13aa5c18a2a938fdc09c9dc386e9d0d368956a0952bfbaef797036991621071e98fa477b02b1a4f48465845318d8c74927d88b961ddccb8e22a27ed817b7b1da1192ef7f615afc6a7db743188231bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a03c6f8195abb554fd8313d4c29c08b6038323a298a73ea1405a4f16a7626ee15fc091e7042157477746877805a4285135a3ca2f2dbbe76449f406b9cae74ce5608f809ec52b2133f67576f730b0652967a565570182f687ffc8df7be05493b75d3307250904e392ad9f5f10adefc667;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8229ae1ef929a3b8f0c679bf8fdc736b3aa2d8895c36c621159b6cb34888cfd9dd201ae565f2e4baac3161818f174df7d3977c27e573bc2bbf4db9c385cf7bc652400d1dbbe5078081e11a8cac53b7d33f5edebbd1a51054a188b0ff6c71274b067b4b2780c26715ee20e5914a6ed6606;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13bfcdfc103ea2a8e6fca2cfcbccf9f4025acc8593bdcd2ad8b0d22dea6e5598f21c1e01fd65827a1023d6e1dea8b5d4ebb916b88ae7ce9ac096af093cb5f4ad757d7edea081306407c8537b5ada68b29ec79175ae22bef30c3fbc3b9d5e61777ae2648983f9df8bdbade2b4377e18ec2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff153d2f606e68d26127d5bf979b4aa4253f7d64ce9e673ddc552bec1bb872280778473155709456367054bc1fc617b84d81394628140e0dfeec60172a5b1f980b085db8b5d16c7fa368a2fa167b8e72f61977ce797fc0fe73b60952503894b08319af2329966dc5d60ec4b4c51fa34ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44c3879f2ec44bf9028f493d19255547a85cec50bc7a621e7d01c3fb65adf1b963b6f01b7d67e4a3e56d43f2e0b3dd5c1ad432ae6e6da735aabf82d63532181c97cf601a43aa35eacb4b487de2c775ab37d43f5ce601f8e4de0598bc4262c1ac33310a654756ce7a18a4b2c17902c19d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc5e5690a1b715ba8258118c3227ffa90691deace97c2078ad8483a15940d50855dc151e17eec3dce71835e916152c0568050879c612e02fc2f235924583326e092fce62114792783133788a8c9dedd8ee444a463253a434cb5f2e9519e07aa39a6897ec09e922caf6d200df14a0f93c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a8215a493aa3e6e9f8a6c6836adcc9ddb9bdfc77dc5a6a6f00abbde491c6174b5088971fa0b28a065768f72e4ea365fd999461927fa5c1d77d14a8d48ed5da29e5bb9b1d18eff80d0124fa322c6b38f210b6d06956688205fa2e751381106e1b4a60fd7692584dc6736046b79f5c93ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f889c169e4f25897e27ef876dc1d96b9f0a861d16e993cf6d6f59a82b969fb7011931904df11e1ac807a48d670867ec9104c5d5d3e7ef25b5af109cf60ed8d249bb49e32ca5cf2a601c15af7ba10941a4a0f56ac2ae93b2d2a9ddbe6d34ede37d8a4b5ea2e3e01c6bf152070ef003331;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6835fbbf8b7417806f1e226ccd06b78d0191fd1495c933ae8f19253d9643c184403915c3c98725dd173e4811493a6220ffa346635ba53e27d266afd171f14332f4dcbc626cdec3dad940e80d921a9575b20411b777a9819697460851f777dfd8b23cc3fc89db148f3d4ac90d2c02d61d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha08e51429cffd3127e2b53eb76365cf898c2fcac90ccf1736431b9c2c6535146b494323f9cf01bcfc7993994fb9a92c011cde888817507b09afdaf59def112026a52608d6400944cb3ccafdb9ad87bf627696b289983d284516048d454c4860e388af8e1aa499a85b1aabe8e2d6e40e22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77d3afdf35ca49d5ea88e8e1bbd00b560ec6d6fcbc7b646a830dcfe363625876eff416454ecfcc454fbfd4f61a6c2d8b050faf288b80be968d5386e2db336cff2c591f80b185dccc20dfeab057eee7f00d9f3e6c3097d09aaa2e0c8c2703cd86abcc549365f268f163bb85c3e236412b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b17b87fe4b85fa1dd3a9c3617151e6f732aa5e0679ffdd7238c689a603dce53b53851704320983b12080ef997101c9e508ff02b2fd88936de3c66a5ad5e4b1c876d8b51fae58c775b366f1ae9f731ce2354120b515ed558d942c51f2221704c0140a3162a070e8137ad31ee8e4de69ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h700a9bc850d32ab345f0e31616cff631967f23b1ca1570a24d31c67986675ee37a39a6901f4df12eb448b0f894aacafd350f24a4447b1cd2901e254dd99613d242a8f3dd973cce033fb01cdabce0ecc2fdab359bdaa05f101403fed3285df908123f3306da45f4b2c5e31852d84147313;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4094f5c5e5d686412887272ae6707b09a0c139bc81c454961531e3728c442f1f67afe5fb1ecfe1be2587b477ae18d1138f2446549c90ed6791d57f306195a6a87ce23ed63a68dd6190548c4c1aa5ef50510efbf184ed406dd13b776d2eade9341c044c319f70abe03ec6355e82072f80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf57cf191b9b25752159a75fd2d62b747afd8ab6a3a5e0ad4c82d82fa8243fa804ca267dc19855a481ec3ce7c33c984f07e5e02da1bb228348da553c0407a74acc3874beca62130c1a411ed2231c83cc11299a459e9618f0132fa774bd879a6b33e591aee15a45fc9ceb6c6ad98614a65d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h909220aea51329a4199fa72d434b0311f1ff928b4096c6c4123485e7aff7a2d296516e71940b6f9e2707e4fcd018eaf9286303d40cdbe1cbb1662655b3ce18ef030b8f514e44950ea33902f77b09a5b5ca1a6b1fb3a9db7cffae594be65e2a9bc459f5507d48b7654a30e3c8940390bc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc927eac55b7def5b4dafd0bcdcc134ab54e629e0d0cba5d540da471cc10b210b616d992f8f05695538cb6c981a73eb4e771c7af7319b5115b679c9aa2cbfa159bef2849721b80d1ab4f79d975d47a30bbb1799db83b886049a329780b3d588a5bc98feed27de35cb81f6744dff3c548cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6eade55f920e1b4c947146b981ff2e07665271cd0bff9417704882ee0c51b7558968cc18840f1d0e6ae6ff1ed029f9180a2d19ea6ced81a20bdfb69b45771415d8234a801b0c60530b681f5402451a9ee5559968f8a00257b9fe2b8dc5f29a297aca65cb0531d4e17fd38e453a7a40a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54c317a35f8b1f612b65858fbaed3f949d3e8962588f024faca86dd518dfe14d11f486f4a8e5cdc0290bab93cd11c1b1abf4e8c02c3da445b541a52a6ee736e68e461467a4e684bd2ce1a5e6a73b99496ca6a960b60e6375dd78d2cd58273d1e3a993826a96ffae69e6f27062a6a3fe14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97d1687ea0aa4461b6a0a5c9b81682b8d3b49432200b62779576154092277b1ee0f7b0978471f32da88f45538a94b4009858b8775c089efca101eb9830807d6b3352dda23e21ecce158e6cf472491b8c0a6b56b0fd8cb1a3401712f5b612a0498c9068ee08d967d1027ff766d59fb8471;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he86117a6c14790aefadb0079680b1c97bf79af5a726f23222a1f9778351cd9163f35df458eec7d9eef67ab09046f0f4ee439785557be622bc5ed54bd84ce4c20d880ef27e714fae9ea69e909d168d4c0c33da51bc7db6812954a6a70f09dcdf4c3413236385ccb0064e59085dc3383497;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee8adf058238153bee222f43e6b080d28fb6017ca9bc535181e1c0cdf3d39e42888916e0e34eb1b03f5a982331c7b85c7f81315bbad6d5aa3f70e89f6d0bf6f0877f254e30e5f7079f9832b7208aebe8ee3884ef1e1d2511c117bc6c68d0b0b46a4e07632c21068e07047f2db17fb9c01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89cd8cee6d27fa3fcbf5ccd3289ca405703dacba130c3e1a66ec1bee23e288c3e67478eff0fb70c1a716daa2f73e42aad790720cec33f3f0a4f8d87b628b355c22b94cd03b9dc23f6c0593983e000efc756492c630f1b3ed5c5f508b93ebc99c143751c1cc7ef297520ea6b864822d952;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ef97e15ed4ad3f0fbd376892c5465bb987fc2d01c8687aaa372f86cbfd99ec844f423e3b22d1f226083327688230209a3e04f6955177e73f7efc3e06b9f425660b6e107bdb68ced121b447dcb9040dada6c262a9646b973219d8fbeaeefafb4b4b12711ce126a7a45b8dd72cb3c95d2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4167df5fb465d6e631d7fba10de2570f23caafe5e5f1451e4c071a85064e2943cc1831b7b5bd29a485c752c7591a5c510a30fa41b6117c605c61023df71a5d1eb75c32eb7e36b2ed3ad5ac6cbcdeaac5885afe9da3974b70fa985a74b8e4525826c66088f1282b6b17d5dd50c3c349c26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0becdcf97740896653a762c18d98c01ff4752bcbd0c7bf1ab080f3e098a21c7e7dbf47084c06acc26a4d3588189b0404b6e056b7c83394861d45d602a0ef3f1c829d3d49b2c9ae3cdf7c740369bf710b987f04e73756b3f91ad523bf90a9d9e95cbdf538eb199f1e1e0d4a1f58c41bb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ee4cada3924e0b9a813804d509546e3ca37bda30f149b2bf327ab3b4bfa79cf1565c563873b2bed90f9c54417a5147fde76fa0caff6854128480d240552456887900afbbebde6b9af420d3e5831a358292e85c4c9121ddd3e4eb4a756cbc04aa965d301f5eb3c51f0a26ffb918a7b383;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88a7863364e38247aabf80492520575fd969c8564c6c6ee933173d3e222dc54cabe8a1dc430f811cdc714dfdec34e85811be2225c0013a4fa3201b8fdf883d2debfaa84271718aeccf78a2df543990ec51dde0414e9de2649e029ed3b128e8219727e90ce1f620a7c8395f007ff34c2ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99c5caa181f16622eae3f06e5d71a9ac9815f8c9885782ce178e82d0e0c8738386431bb9178d890d38f0fcf5ab40877673d6cd95d463ce9a3ea76e930e77b13c1c0f3e61cadf29b5faa6fecb6930cba9a8873b8670073694e7ed1e0a25ccda8ce0688e64d5aa399a909a16465f25d6603;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c9b210285e0277c1786e4bf408732e9f1450eba6a7caa2f45e086cda5ed0b790b6353928486d5b7e59afbedad0c471079c316bc61bdc9f02fbf4152cc25e0db2b638ebc733a98c830cbdd0f3fc152312890bf30441847c6cb611bf54ff2fdccc1e048cfd611e706e4156419291610770;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha77057aec25cd3396b1af2bae32ce66fd6a84355a5722bf7159e5de57a409c8a90aecc2c89b1e0af856591de42cc4c68bcb2c069d04bbb18e08b7049b58f57ece0db32a8cb0786e5f91347463b348992e60b2c5d9c1d4dc42e1bce8368173697e63c2df8000a0bc8ea99d8d8e8f1742c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32cc748c99c1248046984cfb92d0f91968d407353f88c526f962e4c8950228e9cd14ce9dd603a3a07aefec59ee91be4fd42b5c165032c6839d52809681430d2a412d929d1f54399413842c49e0c41fa4a3d6b8799eb6c654b2a9232584c390ef83fdb8e12e97a84dc062dd0995480634b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e78ace5fd729e1b5270538059af4b0c8227e698690601e9b8986cadf52de7a859474b6af0ddb311bb29095177be7e692d0a7eea198a003b2dbf23142bf208b8ad72692bc4eae630ef564fd544cbf9e5962afb123b530b6f0ed3a6cd42912c8abc564d46bb6e0493c7e222d2660e1e048;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21c74cb6451513c6d8040573597ce683e5ee93e374471307b66056d273126c48c9bf6c17e76b1ab8fa89323ac71b3fc6e0023fdf13969287ab019acaf91c52ff49f89ce76ec308b594b4b1b3b72df17429fd661cca412e6aa9a8b85a1255545c07bcd2d2e7229d9301abddcb08287d229;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc75aef038bc1245d5e98952b175d33af89e04a23b93e33c9fd00894fb90358bab362519a1856f9d5e8a5a3fb0029b03707500e1ba924dd45263c2b09337977cad03cc68a3acef2c2aefbf04267d0a649a99031f98eaaf780726d9f0a56438b10eb7fc96b415e97fd038aa624248608d9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39296f92b96b50a1fea2a446e67c9a51e1fa899306721c35aaabd84cfd330fc1dbeb28b657dfb98f6ef9001f86a621149e796696960251594e4234a4d93a4f93afa0b40497b0497ec08dfaac51a22c51c05cc2f82b220560823e6b32b68e11d4832ebb634b7b6e36bd7bc02bbfc4ba485;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50413803b7b7c628f376e6f421327c55fd2fc6651576bcb6541309edd902eef712a2c8ac7846e7f19f798dababf8528cc2afda4a160ed8c2ef36b9073c32750040a4c1ce0bbcfa1ab05c5e20c69074b0f07a7fd262912017f5531c0bfd32705afbaa4f2e9f133b2ac0518e6a30dd56c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb558f1d3cd25c686ab25c3965ff1344b141fde5cfa6afdc299bd2a3b1c24811a118734c9d0d7851bb0dd52390d80a31019b0f2dc8d7b795ec4076ce626ea15a02b10fbe49d30046a210609ef63837e673d5d53a56d7a5432954fac389e1d7ca55e82212224e2b26f4e27cdbf936d7b20d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69337147a1776590cfa37dd9e12d00887488d6cf5026b661b1e56c31cb099286fa5d3ac9312b03b38bd571544127227773161e9e7dbc2870e552b47b97f1b3e417b544fd3a145629c4c2c2d521c49e5f6a71336c8ab7769ed08fa2dcc2b311f03ee014092bfcafcce92184d27b287b822;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h304939a1af01c8321d8780577232dc2aaa644d8275ca2a1d91a96b8c637d008632267e77266ee07cabcf5dd9ef9857b01d1077c36fc314c3841076a01f3995aaab1ba601027b4691e4eea6914233ca6d9b576064b64dd037b89016711fcaf2819a424861fa1b0b5647fe7d4b3f1f8e446;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68ec4812e7128bc7d76b2d60b46acbe3373aa818256f942c193efeb8a54992f26b725e3dbb24e5703f763ae049cf89c177a4c812bc334a1ca518c1e2e2b6de87ac64efa524358f4010f1933393730cfa7fba363f5104d82e26d4a259029d078f037821acd889e32264e4df040b61b378b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1853021cc87ce5a7667739c8de4b3bccf806606abed3e14eef70d87cd644682712b7ef88fe29e2106856d3e2882d1d2226686b326a76192df956bd9a769853aa61d1cd56de75e94a2de6c011b69874a8e8ea7660092820a4f5cd6e90cda532f684a9df262dd1335362405c593928064f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdc130db0e04fd451242b725669897cc7e11d520bf7d3e00326ca857ef818dd8dee4e8ced7064309ae3b8ae0a4f201b5ac2fcf9dcc51cbe0ac782b4c6fb5d2a6fe12b215378cd89079b2ec5945ec19c1f785bdfd68087b5a5f71ea901e76ce5933bf408143cb435dcfbddb0da1774d057;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50fba42670cb4b3a72051eb10bae19f5d1cf015d4edcc61e411d5c0323382174785a2f7e7cbd2cd703dce3d41d13c88be100ca314e03047a9e6877074d5a3ef6075a266df29e90f26ed6f1bfdd82e026940a5528254badc40d0f7e8e25c283b18652089c5ffa0e70d573c059a5d3c67d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43b867793d36e667bbafc36df5afd3da028ea3edce92737c8695879833b1f4188844221adec3d0e7a4ff99d09b7f7da7df3639a7d0573fd78bd2c5945d658d58c81d49b7740869a2d53ca523973d4ed7dd8238fb1b72419c5cff171cc7ed5323b50e28ad3174cc1e0a65f7af8066ff6ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5373fc6862f457c5567555f69661cce267a0231f8590c6c66fa4791fac278f56e9b8eed73373f33adb3ad6273732888af0ea8f1654671d383a661a8d5ed339e0ed0968dbaa4608a0b117be3236c37458c2837f52dcf42a1cee4e9e674667f0c3926446b8ce332a08192cbb3ffc293c322;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3179ae6bfcae10a7fd85421e4fe6ed42fb88953ca90f61b103e8949d8fd617317b473697b383c2c4698eb35e0c83574a6cbd709a55bf51676c3df1d2751a265603a00e67c389bd492721581c66b93598efce9244084c3cc9c3fa02acf5e73ee01c4bd6fc5ce3317dad58efff0302474a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e016fc9588624acdb1a4caa1b09821a9714d1135d03be50d0306707cb141b4412f017203b68501e2860f27ace81dc6caa89dffed369c77fccecc1f36cb5c2fcda1f12e8badabf40d343144cd10aa03c3033040b1261c9791d5172663c17e84cb0d1c79a3b8412caad1a53ba4e41085c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5755e89167a5d8b6b44fdcff0b99e075880a367a31fccc444655e0675b4246e8f2b3d1647c1d7cf9487bf55912e30b41aaa20e7197ede56dc0a919b3f342f58b9d4ebf820d28203aa53baa04e5d743ed67ad2c089fd9e07adfc288e844f128129ee10de5fe2b94736c418d8d10fa5e74f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h459a13eb569cb53bed30da7732b69cd0fbf3dbf7f17fe2e094349fd00a98723ab5708967e34f06bd6d37fc615f5ab31205b78c1c22f3b7251c5676b18f2c1513364276b7a46129055a3cbe0d0a0cb63ada03ba2294168fd10f03e714152bcbb567d6b7872f59aabf75d22c809ac6c240;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67e6f42498aa036df7489643dd35f2659cdb7340018966794df7de6ea6a7788929e1d885d4c52db7217d3e7e46df11c5d091e77fab684666800c7a27f700fe9bb22461f95883d16c4609e6280277953b8b216af48c925b1e24f536c97a0c1aa5084628412a8f648ee7747c5865a8f51b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0178cc9a616c13569210b49e436b78fe0aadb3d82329f7a872765654ff59c7d676521942ec866f91d637da7b76bd85cc301a9f0386c564479e9bbe1bb552930019d81f4e0a72b43537c3a56228f7cd085145b9692cb98356417d2e9c6fa4e73e66bbe92be32ce5f2b8aa12f4461121ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d3a371c7621ede252c7f312eae7a154fa081cff4e9cc5298457fc281acd4f3dd56a6caa02fbdb6e4a61b3f1baf27fbec2574d301b5377d972f86c0c484ce13c2511e6ea1060bfb6d6cbbfe292e2258f94fc9d84f8ffb5683f096c180d52a4b0566d2afb594226e381488f2de03e86d5c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15dafcd413e822c677268198d74e77fd5b66867e7b2968699695c3631457415b4baf7f885d2c3110e5f742f128d1a335a2eaa9167aa754dc4e2a2cab07412c8de9d63b571d891430cf3a4a8d1b7edbb301808e640e386a559e0e5bd02027d74c252fb3be1e6d3c4addca676e6d93ab253;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64ddcd49cfb3a652bf7383512721b2168ca4808595a40f4db8a07abce4ee7df32cbf97bdd1c70a98f188edd61209d6d17dabe8fad320af492e5157715474071f19d06de8f4207273bb153b15430ee63f38d521dbc66c87b6397f8cbe8c8ed1596a1b520b318f50426a91395c22c0e68ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf597dd17b346da8a6a5ad5ccb5bd3e6e065852d7d707eb8f8cc9af66c76f42e3dd8498a865a11a867f1a2ca2cbaa978347af93871f1ab73ef433cc42877ee6a0f817afdbdaa99d145a69241fd23d7344ec68ad048520079b8930d0ef04ddf681804bb09b0eae63a38801705950d5614b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34e19fb67f56b4e96a22040b16713bc972c1beb1ef337e31c822f95325dccb1ade965c9a77c6b30a6ad83dc0d68d6a8b0fb3731b2b7f9555087cf769f52c12be314ae10eb4d830294f9eab61f64f54674fe25224259c8b0f78216d482a7331aadcc6e0003f2cc6ce68ed300591010f36f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd47dc76a94414ebc41eaea493fd94c40809cef853973f3a424ba8872782267548aa6db1d36b2257613dabe2bd97aaedc90ad0dd0fcde51d211ca2e95f9fc91f8567d04005bfe4d1e6dd5d81b856d9c1a12e62b0f40e2cfdbaddc4590e380423be9f33a326b2107bf63fdc49c3779d0a52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c2183eec0282681f27589778f2893b4a94389e94232c0ee6abf9322e4ebac738d3b2f85c8c347cf8ef4b23f4003ab8ae1b024c43c583c210a65dd6b23bafc1cfa66b17a5851f2c39539050d9f63749354c05b6379fa6e25f79ca0f864f34284aaafdedffa32fabac8c6e578707f37d2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcae247e13dd99266da390356faa8f124a03f0419a1a7f88b0bbdb9a26d9551fa70d3d8dad48680851e6c2b5a13626fa237cb8efa588f3fa9e8ae277b6fe1e35182d2f3e4ba2707b62c6c50d9ef62e4d96b7629b1d7f82afd27e6f54f5a98a0f3f1df8beb28b05b72df704d124c6d4bc5d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafc5b3575f69878c6c18b0f342b734c414ad6a910d290a269456eb4cd0c0f406a919c68d36eea2396b0fbb0a70a4c5b615803f1edcbfa2600701a0db63b91afc6b5aeffa5a59b6ec3011a8109c0bc9d7ac164a92ad96b888503eba24ab1f71f39249fc15fde58aec18c877bbb1f691e0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3c52ac9dc1ce0c0d540a96fc720f1e2191099a5cfbce753553837abf291d4c9fd9d41e14f122d1e96b03fdb7467a89ecc8f8d03bb1a002af250d0c45c0d7b9c95e7fb7df2d92ea55ac406edf3ebd1f7187023e09d5dffb7a2a93565479288ae6b70837cb3d8f86f8a33e4cc3fa5939d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb48de83d8f1213525fb0222060428a61cd5b804ead5958e29373faf1c5d44ebf6bb09876203b6cb59f4f577a0af22f7d3afbba1dde72e9589be3ae4ffb040610c146330244293d3ac5afcc388bd0a03cc818379c54822d2239c925d376fdb3bb930bb1691b0f3a260fc832ce0f6e8d4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cbf02c162d636c8f5d8827da314e9f0195efae4c60472b93e1011c1057a7a2bbf4b7703a04ebcfcbac8d5ff1ecb223e5774b96ea2d0699e11625c8e657d6a41df6f347d17a3eabc3c80e854a3fa1b3c3e16df98d71e6eff209239385f9ba7da6dc1af84e68b236085eb368bb9f117601;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f2222842d15e1962255c50f54c2a121658f80810f2911cd8519914dc591228485972cb2c19e740eec07f1ecccbdf718d83b426a93226da5ec81a3b0ffb56c0f069bd76fc77b811e66417ebb153d99d3cc2427b5174b69395bd394d351a21db7419f1135ca3cf62ce5d52aef493ea074e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fbe6d65eb655da54d0c1e458de3e4b8a3a18fab07ee40f6d866896fc571dab2403266ebeda2326072c81e8ba3068617af03ba544ea2af60b1d47004be79446373d7047e7ce075314dd3961ecd3b3d828ce0bbcd01af25d869a62421a2b1c90301c3c9b1c5602ddd42d0a98bd3d327782;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e198aafc112043037f37f8cba715d4d0aa8dad961c74fc2379ecf4c0677c430e2c1d84a7b93a22366f4dbe6cd5d48b76e8eda2ae78926c7ca5ccd9adcf57748e55a54b4b792fe0cf6a06b1a744f5893917791dba5ab258a122ce7c6e0f7f73bcf4c4e44e4c9310f1582306c0888a0ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hada6eb2e6bd039f3d2b096e58f04aa42d9114521be7dacd03ccf2ff74dbc7da251e9bd8bd3f9570f1cfb2281f2c9a574d4668e79d9b80d2650b4586428cacb985c00b893014e0bf6e66f86c69f763fd12ff96cfe81a03c98ac89761ecb62783d8bedfc015ef47126f9abc2bbcb6097507;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb47a9b2bf70fce3f726ec6a85a7588c80b8dfbdf2508f5b28c85635ebbf3347480cc7299a5f4f49a6a46969fcf25fe873706aab053b615eebb7184a4ea5b5d37822df55374db418758907c64787bf415b9257a5e05f81c566c999aac7c90f1c32016d503c3a489faad9f2b10684dec373;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2487c010218b2535a4b513388a640bb5f1e6c0fc71aba15b014c99916ed65804723572dc64008062e8f34b9e940b1bb8ee56e1fca2e453a61d853f84496d256ff2fce2d283ffde69a631b9f04c2a5a0a87ee5df310b618ca150f0a2d76c19658b1a95d379a16512585dd45d4f030ff9bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55c17bae8c21e071294d3076afe2628b3627ecc8b1973600bc0dc8b5d0a686a96863fee8b45e5411adcb5240f512f8deeefe14f61a8d539085651b3f5ad73066e70bb50ab5301adfd26af66f98e65f25942b28dd15f228c11f0976e9736ffe538b09e520d1e4de082471a4e17a4c679cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf253c718d4ecd5f9f5fe8a7f9d8a2955bfe4fb404abf3c106804978aca9832768e26522b9e966aa7f4d521972c280f811dddb9f5f81c6083593bcefdf9196a52e883a30afcaaf12cc5fc5b8a765122f121e70bcfc4f887f7b1f6e5dd0265d381931ddf637654be1bc95ce6053a5f11b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b178f81e25162370c0184e53713883a20549c0b0080c2b5e0c0a25e6a4c3311555f5fa63121b5c80132ab1f8df744fa8e343612b79c39334c1b310b1187be784768398a2a3f6b710a5e12adb131e101a13d24d9be6d5d1b9c950b3a0a5d44bd019aec4ef947da5a855b324f9b4315c7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h772f7d693a7cb7b779fc210909342a0b3e950b0b38a10ba2be07c41d4b3ca82de4a9547f7c56f0319dac4fb86c8545e13227510274f5ed65fe117331b51d2bcdffdd06cf21ffaa48a141acad2d78ac8129f642b274eeae3d8981f8f6786014157a6d0508fb64b3a272dcac993ee19c1cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47209066cd5d2517e0125385867879a502c05e875bf22ae0f5c7b0337829e2ac622f50d6100b0a828ff6d064d0049beb4a7e5b3ac927d69177eb1dc2cc41e2e3affd637b794913249a387db5a064dfa9a0aa31d92c0bee366e198c42128689af8b9cf9234d5e0adf8febb437686e21796;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h955e5fc9925f0e19bc79acd29d6e19f917d44b21a304d669cf26a4d6fbf7c6c9c2ff70e06912875ac951b29d88efd3cb66520657bda4df470741a367280c3dcbe7d80285631b2e9edaf457d622866aaefd53e9543f19409740b94709761a84580abfc88fd666b074eee86880c3c444f81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62b3c03c43702100da86b80b77cefaaf6c18d06c8ffdc06bb33865760ba9927d61c2adc922f6c79619766706d32e0fd246fd840a0a3a4ece5b04678ae13f565ccbe8555c3c212ab7b8f886224984a893a8f5e4aa9e34976827bf1c202d0a0542688a194caa27c6b2d3dded70e9b96a629;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcc9fe588363cb2357c3db6a8871c1ae733741e5cd30930673aeba880c7743dc4bfc349b8dce415b35136770868c110c2c9cb481eb155bb00e3d1c2bff81c37e17970611304b928a46e58ae3359816644e5f3eab6299ce6f02cc3ea0241cddf2dc7833fd7aec437330ccefb869c878651;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6d354c7af9a939136fdd24dd3683a74e4058fa8be63f77137fe911c11d4cb1092fcfc4aa2acb7fde198a123d7c2b792a68025870b1962b1cbe1ef75d48b01a44d604ebfc25d3adfec25d5c540d0938fa1960106ac245478592a3315c43ba1392a234f0c1475ce2f7ae31db623f313596;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h340f562fd3d35175de2db87d3a8427e9cdcd921a2cd6aa110065be7e996670ebcb485ae367a4137e5ee90c0e025c02cd2d9a7be224a43d332f9763ee60fb23dfe8ebd80e3834434f87f6d606652d367e483c6f5c7a94850a4bf4956733d041bb252b24cd12a38bc41861631fb300e5658;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85ab5d9b3e89b34a75c27622bcf1fc62857b75ceb233c4bc49bb39f2d8bebfd316306ea2394966fdae58e9bb70f7ee70a2e8487d77154430be250525c5b4a1588dbdb64b10bbbbca9911371fb79bcd38e11bb86cf3df1e8dd4e4c5bca739949a63e00bdc4c6b462e23991b8fc0b1c3094;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h654874c0fd967f8a40754b2044ce991b6ed2f9aa330514d6f4c3be745fb301fc4fca4b23c87404f81aee72d211528d3728322a00da5e79876b79378f1cd8f92d87b6a65f23e94d608d79cb3587163a6a0c5ce898addb19115cc6b1235f45e31617969fdfbccd427124dc3395d2b1a1822;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7e57a9ed744a7d7b067b5bb654eb5c0eb07c3021abafb34930ac163000bc93425b3b39d68ac886cfd1a66c15960c08b439103a34e6fb325931210a068b952f585562c9d75d87917d73d3755cd8bcc496be534d20b3f88182b2dee2eb949ec2975bfda3d4f0caa88aeedb0824011bb822;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h798f1b4e56cfa581a0dcec0befcc89e909e7fe3d7e6e8fa34ccf3056571ec6ca6013fe690180cf7dd6b9dd8700f97268c624ec3027ac2bfb19f9c934b9541bd778397a1115877219deb47c6786b50c139e8c88d3031dcfd462542a4f9a45b40d22e3376e2c8ca9aa4a75760326926680d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e242f65e73479dbcb8a18dad94812ab7bbdc9e050281ef426125d7444286020a2ff7043e395b9db474570cec2d5a236347a0cf252248ba2fd2af0889cf53ee609178489c9b7f0cc113070f4a00fac8c03e1bb9027bfea93630df18a3c8ec2713172882b62ed4a5b006ec1de0c62a655f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf13aedede5cb1793b959af60a45e5c13501ed27a68a0a617cf27df8e5c41ff1e9caf63e97537a725337fe85c0f1e76cc085c1c26822c740fff90d8a447138a6a5b444337b41da6c5cb1e0a746552ccf4c32388a216d64cd02d7b444f457350a08feb6fcd159d6e16a3479ccd294a84f40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha36fdbe3d0fbefaf0d618c234df8fd6ed458d92733be50624a3b4306f34a0210da649ac3160a1145476436f906d694e8e86eff641ff520c616b0daefddad8a9c03d345e5937329ee9db299b4973a43722121ca294ca6dcbe4f18f56614f1809568d641290e9784e7f1f28ac888370403f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29e83441e7e30709c731064eb1ffcc431e5e765d63fa3e626a25c21040375baa1db0c535e17d686798b50938057bc629035b4ba89eec5a81863e96e3807059958c9594722bfe1828ea1c0918bbef6bdd58e9172fc91b086519448269714a77fa0f25ac8db84ff6e50c36efd43d5fed50e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e137837e8773858374bec0f8b71e599599ef111ad477ddc14545220ec81d7b3fa7e7d2c7789a34f15a6346d66fdd397d6cc0d01a2d6e045c1e5913453e740f187319f79d812d7667963faf8240e1ca4b51c1df5d5447f773a78caced20ee05913bff4530d31f90d8e0c04188efd83dc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76389f62c18fcd54d90419c1c153815e0628ecb4555507fc9f93d1eb676e8bb72cc7cbcc9f74bbde8ff72a8f9fd5ba2c7c64da396d7782dd55e12b3307582a8f328ea6aeeac0ed556c31b35361a34f88c1c99fa2048677dae3c87cf5dca21dcd4ca934e1cf6087ca046e476d6a57b35ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79b6af82fb7de358377a5457d80de3f9aaf1ad32c05a2510b740fd36d5e698e9194a0e8439856ec3226dcff163339124a1a15ea67422a7dbf517cf5f2e5f8a9da698a4e72d8d64660fa870051b790da17661597c403b7ad62b71f72ef9ada45a44c755785b56e0c10e10c6a5495040f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2bb442f5db5a9b55f12a0fe7df1752df1aa60ecd3fb86c442eab7ae9e11541ce85db26125c67ec872138d541df4a3b04768e505d3e8356ee7d13e8ea0d73416790700ee2696f74656484ffbc132013841979a28a6c11d992d1d587e6adbba7a6d2b881a39812095eb516b47c7d089c74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aa76ceabb6463c25d23614f5cc6aca015aa3b46baf1ecaa35aa5e054c17f3e54971e834931f815c070c059ecc8f3b5dfbce11a651c60a0adbe4b1813c5969dfa0b6041fca38cdcbdfc465ed970abe58da8afb9c1a2db6de8e7e122973b14505d1bec0826f8b93d85831e3663d034264c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4741d98cee188a4244009c6d0ed7e4c7d6c12b3e7edb8e24f6877c048b252be80409b183ec512b9ef2aaf9d64e37a6260b45022ad54c8bb7ce7ad72ab41e918b6f0901476039b990f0cb7842710ae4c80874303c61f347099896d1aadaac0c0c43b9ea875fd9aabf9f76d9f1727b8c47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2e6419f6dac6df515e81ffd7d574d980de8788368bc3c58c702e345ee3baad268a1519847faa8b984e5cface944cc827d4ca6733ef6b6cc117507c31d3c211d5133a8278638df3aa1b46093e9da7ee7061a443f7155cfe3ec04996620cbf6b14e7089603366df717c86dc0ca7ebb9d02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he59d08df34853adb232768211533fa16c12e7dd3fd4d3a09f1530f513a674604f2eff420a1513f0d695388203b6c834f5fe88a1edd5d262b336da2dd2239638184a5fd21ee2602e607ec964d8bce320c8fbfae16a0d5e065b8d297653d06eb76698f4243db98b2efa4ed04af3d47c8994;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a207f1c36cba0abe2c91700ad583d2baf0b532661993de1065bf166c0fe46462c7953437ae1c0aabe5b5c72a941f4614b37c853cec8cc1bf35bd5ce5f840a345ea5da48a03f27db42cdf7e16e35fdc9e5904dd4c19ad0761f9365ccdd63ddd879bbbd6ed6fee03b97cc1acf30296d3f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcaf858361d9ca4798fbce141fcfafd9b43d68aca0348545b69f2b46069dbd81da1fdb405b0c5f837dfb75dcdca47a49ef1951c5d1476d87129485a64c6eecd2670cb829e013ef702895e34e5bda99d63974b1863ccc05cd5b2cfe7bf75b523fdb6639a486781e643ea42a0245c5a9b04;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32fad87cd3e81b09e506408b4726a822dddd91ae3070cf14071dc890f67c5898cd4723cc7d92b04fe9513420e24179dba7feb6de0fa88ab852b9b75cf6732d6166a5397b732cb80fa3d03f583da08d987e799a0c961eb18212843a0308c995cef10fcd6884f29d087bd7b70c28f51df1a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21cd7e31496e10b7f418f63df683c3ab5a0f78e57d6c0f95c9a44ceca174cb446ff70dba95dd3b2e6d8d753802962697b7ff493491e3f6cd81fa09590b0285288a97c86dd84af061b362238a60c909551bacd102ad74f08ca5acc279af21d7a179e610335b4dfe17c20d8b2bcd6a7aaf7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87d70cab7407e6864959d7cf0850d8ae888a701057ce6f336af0b0d465782db71c4c77a166d47f4dfa542cf25715ef25821485486034e5d1fc01a3c5b7cad6cbb3d4b35b2c33689c3a5f521ab55d0eb1ed5371eb2a7c0f860a42d84ac04a27ea5cacbd7e0db683fb496d4e442382136ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1557982efff20eaafa561f8d241625c5d3c25daa01acd6d722d7bea24711a7193da7e6ded043a760c0df19eb39e3fef989306b778bd31e5933932dcc9909403fe9fa01c254e40ba7c45de7049bbafb80494943c22db2d7bc8c3148c5c2ce2ed27735bf502040ff436ee0a7178165d5d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf57697a1e07f5a2cb0d5a8871f584219f3935ce2df9b171d058366ae5f410007174485efe546483a8f3c1c2e45dca5a5196b7f9bf8ad963d1343b7ce8380aed666dead7e85c66e6526eb0dff95b361d55f783f83f8fac18c1edd99b555c78ea938c3683fc65e67872e20edf828731f024;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he859ed91b8df22df89ac8dc118adafe72ccbc26d08937ab63195c4f7cb07c723b67978849050de3b58f180abd4a424fb9518aace50ce1417a764b775bddc1e052ee9a2cfca9677ab196647fdff92a84053bf3b3fd0a49e8ba02d1a9a8c123fa671326225bb92d029bf2c05518437d613e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h249a6d5463738814fcb3735f04781618abf9992f84ffebc0905c4df3f1616bc44ab031abd34053175d517cb97c09b0282ea4ffbffd22a23347be16e3b755f35bd5875afd8096b07a9e219e8c27ad84568fa4588da850d6d150579c2f14d102f7f553c8608c48a9c306af7b720283bdf13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ad05368556e7b22af819707cda65b4c9822e92ce45fa4ca0d515593687a906f279648f5b8b769289daaf197187e0395e57caf425681ae95801a3d611390ed743dc064bcf5569cda78c10fbd77705a6e4803c78a18ee611b903820937f4738d3b956dd584a0063be64c9728004ce9e9a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a75ad8c9b647d0ed895201fab55f7c66a84dab66790231259d9fa6aeb8eb882b9f92cc89b33967612cce63319136e8f2ac4f4bcd400e49c5619ef08294d401b74e88a7a55cbad7d506dfff9dc3e55ec67aa3bc7d2ca62748935fe9e7198c995d3ae5e32e910cb8db3b7c1bd840036dbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cbbfe1b75f4240b2d7620c37a43f8a922ef7722c5d495d260665833aae715fcfeebe3d2ae7373dcc7b80ac01ccca69f8aae4fb9f04ea0415966fd67c38de12c9ff76860033c974983542f411a907292dbce93a182b47d613e71acb70e06092f668719be585970ee7f152e7e3d5b6a3ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dd3bb704a5e8a7e511ad3de57f0c164da2afe44e31fa96e44dc369db3475c460d51b2d9438bcbde69e8f3505fba9c4bff5c635ada39f11a7131847a86bf57d9fb9c73c247394e1f8fc2a3adf0d371306a60769b6ca7ba806d302d02c715e31261dc134231853d45c1e5cc45b9238f94b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he39ffcdce0beb199c6b1f51db380e3cd6fb989965ca6a4204d88030d52fea6eb4f477cb94a81ab830ac2f7041f6dc239cf7e508b7cf9552bc832f3203bb0a9f382b4bd02d5be5381762fe99eb82ebe87e81d40942daec95a211b0ab1aeeadb8d4971fdb036b84150940600f8ea29524e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h821b57b13e9ec413302e28dca9a130ac0a50dacc54dd6a6b9b44fead65fb926505b52c2b0644363a6920c634ea1ca0c6027c5071d93b4db0e8f635802e7d0f152d88efb3141e4cdecad4990506f7115337001478e2ba5112c43a97e567627dc4006faf9951238125ac3358143b29eeb53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h305dc02bfe5bc3c7c2852823419f5382341c3e38c71d00f4c72faefcb95db6dae580f812bca51cb9a669d3ef0e6cbd18f32479ab51de14946d7e1482d5ef1d79b5bedc62d38722b037224336b9ec774047e0b8ae9d5cc8fa795f4acac4c031a4aa434a2f56bb1cbbbf0e498cd70a92150;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82673ee72ff4ea9bb65d9a8e09c560ea48b4fd34665599f356bff888df9374ada45e8b6553c2c051abac80e9e670bb6693c15d3e9979a05f36bc7ff11415b8ce6a97167bc4aae6d789cfc4fcd3e605c22a13c524e75bb84ff8fd68ad8ee3f4d5820e04f8032f952d3b6e31306195f7383;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26b217b8cfaa83abe43db1cd3922684b7071b73b0753389177302fef6928d813e45d9331320f531693a37ad7613b48429f025bbc0801f5978288d52959bb87a15525f1b496b747154e4a3d38623ac85861c3bdb675e62f21e8ac00ebf960fe2828c49f82fdbecdf3ed784765c5a3830c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb448c5d2e6493b26dcd61b7d1e2baec524125bf6d27f2b79dda207768cbce0831b22ee448e2be17c52a07f63c81b8a2295d504a180fffeb6c3bd1d4775fba1173f646c335171c8ddbd72240133ca919ce4f39c32062d85a792330977a90d952da1433fb4f141eb60dff68232b273e1aa5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60f1c6dd03536d107b619673610c708d279290d7ed932a646ebc0f292bc03ef289b1e0c5b3558ad0d9ec65037e539d750ee36ef2be22bcfeabd750c4672c1bde607b46bb17780de197e31cf0a6625eea8ee358eb1d1a5eabbd43a1bd14a384815211b36b0df8df1557ac4ab6618f179f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f2968118975c4994400d6146537c8d4c22e14571e7018046c5af5daa6e1c1ca10f7e9f4df9fb1ed37b0c5390192efcaa4e43934359cf94b71585d812952e2250d05aac738210a0fee1aeb28a196230a5b3895676fec11724f0a6b10e6daae9e3c3aa17398150fa1de42549844aaf3a78;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8a388cc9b4e3224b49b0587f8586a399d00ec371ebbd9ad63c77e7142610f61f4d3d5a3f98c46df305fab1bfc401785ed8f173a51c87a6c438ae03211e8d4cb6c13c0fdea9a2b9c2f6e98a07dca8d248d52aa3f1e085d3f18d1f79bc121be6fb1fad0d267dfb14ea61a708cef9ae4772;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb60ee9e4fbc23a27aba1e8e1ce3d330506130c2eaae38f3bc49913360c7cecdb4ff8a1644fd9a0a2b1c4c69317c31b21aa5ccb48b888f9e3d81a8c6cd8bcb8a14d6c6690b6262aa962a6d92540bb1c26eb2683a5abfb91f5f902ce62ae7302dc970009ba15ca6de8b11bc2d6b900cd7eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb5a1e6aa9b360b929ad689577591692628497d9524e5451f22b90ff51c23b64d359206eae691ffb66cf66b3ed0d00a20701699c52b3775ed97b2beb9cf7a1fc6d703f508a8f58a36030a8d16dc8ac7da3f0eb5da0c5d48261e96c30e6251d5a650ff0b7f2918af32082b88afecf340ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33165279acbe0cb1abb6d1fff26d64b3d6b91fa60dd22771edd3896cdea07bbc18ef7d12d301925911a9b963a0302ff658e947ba905e40863fa8070a8881809afc46567cb746c4596f188a33eec53522499f439a7101e4498d9cb882309d71530b68a1e4b9fb174d3cfb1989dce67a31a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4455ef4c3afd410de045154e2fb54d4f0f3d4785817a45eab9d8038d8cd9701d1dc96ea8d6b9cc826b3d04dc3aeee0ded8eca7ebcf1feafd87952c33db5299e1f517f24ebc4b5c567e647848987d97d06133b7a6f776aef23760e4464201d4a41eb0ee4cfa8d72cf5e03058120469e039;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59dc6a74ca657151070a20736c498f65fb0ccf3351ac2fe50dfc846f173c9307651b365601603e6e20255f6cfac4704efc10d50f3f07c6f67602cce0fb5434990e1c3522b9561cc42e60822191d2f30e3f9bf678112fa5358ab8a0761c73f717779154c93a9bf6ef31d4d9facd5590eb7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd87f218d9a65145de325738c0a8279f8cfeabb9310d57b154810de81cef0ad99e050b9cd1bf2984ee0a25eff3ea5e3ced6270cffe2460140a86c07f59610a22f4df99f8c50448f9c0fa0ac7ff78037bc9f4598df213b83b8f1cc42b10a964a7b3c6a0f5822bd05010d15d95dbde16ba08;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25fa63a2f0e9cd282bcc52044d8ac7af32fd80102db314fd79e906044ef7642b95c1cacb53cb75629505a5d734f31ea5dc7b6e10d9509ea9c2be3e8f77959d9d93d2ed5a4d7d46ee184b86b7039f85efb899f95338d58448c368d5f44ebdcfee95961b0adb9720df21d5844a3b2782413;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fa2998cbf3313dd93b3d9d662a7080c2d92df4d859119df4b5613bb242df49a0890f384dfe7b7a77d92c7302bf6e750e8c278d60a491a3052243a5dff055907efb7191d30cb734070ecc025b24efbe9825f227b253447a65b87b6a00601babbb9f425005dc006fad01453c2cd30d034c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99b8c830c6b56cd99cc6cc962f0455554951f6b5f1aee224a30f4d4eaa45966fc3465f392fc53285723b6631c8dae929814fe811adc96ab0ea3faeef070f996ac002fbba15383e634c31927555e8f2737372871014f0fe4a66e44981861502265ef3532576f504881270f1e528a95ab14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb6797bde59ed5cdf8fca23562840f12ae2307b0e282e7f1f9ca109a28e87f1938cd9f76f38bb3e76eca3199ff2423c390fc45db32f51cbc10e2d9b5f162246892f821277249818ae52587b0e99278db8f769f238d5f9a04a65cc7861340045567a870087dae1e134f9758ab7bff9af84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18a85469488101f6ce9594047d848ad8a969285af619db17204a2bf86ba4bfd0b0c927273c897e3849cd455b0fdc5efbc10cf2d2c22f4e0a8460821baea5cceff98c1fed9dc5995625f2e8b72daff784b9b5b73540c71ac68014f1e8660bb7e81b80b31c56411415846f349df5746e936;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8e23afd74a3d7707707c08ce379dd1201b259ec6aa0f5c1b79bd516906a49fd32ee54daf2e5a3c8acfdf502f84e971c0587ae0f2fb4395bb7d755c224fcd3771815d98552b87c1b39f63e268f6e8d73b57d0ab18cd7dfdd6606c3bb10b5b7a4d17531d2f52d0502e51a7cfd6f4ae2346;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30d716429220e33f2c23efd1caae648611f34f9fb6b6a4101ed177a0db396db3ff1e158ad1f112e1a01876b7807bf8315e25e2037c86ab692be452b57cd575b631f5513fff5fe629ca8cca88115df266b4d1e33ab2c3ff2f5af14ce5652c1235e6ee422c693d4bb53c0d85e2bfbd6fe72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff194ce7692a7a7a665f4de207e34c209c8e735448285fae0973b79221ed0dbcbcbd5c4aab422ec0c2df58ac306b266e20dd4cb95812f4e1df1ecee5441e9e6e9aa82b48ad85b92ff3099b89b038e3ddb10f363d919875d9b26f5e19d89d8ddbb5a868e990f76379f4289f0f7fbb1a284;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6bcef779e6a8e92bfda5f8e3f84beff32e00b46716e757afa073015be3d37e439bdc80969fb33efb7c39c10c50bec83ce08a3e50d2eabb9cc0c62e1e36e26bf5c2d597866e89c2103bfce51264566de9753efcff1f55798408a6b92f3d7c26f1fef971e3bc3e427835e64025f75a79c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h565bc251ce9f16cb74eb23dfe99c1b170912295d376b4a9e6ba3a5e2f2ae602f75d4bb810c16fa3b84706706387978d56f7fa97b61e322bd4b13591aa34959ad0649e5c5732853dafc1da5835669376bac6c532f95bd1250bbcef44a935eaa829fe8a09c779ec2c329ed709ee0e0d91da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6990e71c7ca9462f6131e1b6bc5ad0af42e7f91221a38de143d13b99131c94f695f62051bb29753c920b96d9bbd65b5803f089c39407deb1d0c26ab4f98ad649b1acc0fb0f1c8421ddb5e8e4e90cc1e56b74d548511d008157bed05fc427832a5c444c10593770509e5d61ec0d075733;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff5a42206eee688e3e40f45b1a3763fc2fca6843eea9f56dd63742ccd0caf1ceb6bc6d044b86a5e9717c8d0b131fa17617f2671cddd961e398ca0a658bd53cde11fb9135b9ed5b695dc1fff9a655380aa494546bb7103ba80afdea47a7e4b31773d5d672c44fe5ab6e3d77aa6cd0cbe97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2135817fb7d7cd0ac23c218a08a9e1f41955d8cab8df6ab0529c5e04bd0952adbe014bee95db4464b60e40d0d3dd522d5a687ccc6643a2a5493270e0720c977c3ee3f7e1c3bd22f07ebd28141af8c1a645babd10ac2f021d72f8d181e9b8a98f7a24fa8fe197a13e5327bafd29a465df4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ab0ef15b2a82f8b246aa0425c901c8a5e36e57ac1b576aa8204bcf26dbd99f122405a38eb5cc9f439e2c34d9ccb6eda90f1fb3d8ea5bd3b547f6cf0221f266bf451b9a95349d2622ea8087cdeb8b15b7bfe8dae9ba314d4fb56df0846cefb43befea1df42ddf91ac3535718fcb9e0c85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80f7a1df7215ed1fe444fa92c00aab1db6f22aa88a49b0f4f17b3ea543934a9e3cf069449d160c05c37bfc5e516951000943dd3b96328cad31d734a61757d06e604637bff447088589a490aa2a3d20a56b618b61ed1a2d079d9457d550c4db9ed1cac7fbab208a9a4d29fbad366d46721;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0311cde51a850f39d8f3a15f2f9776da5415b4bd6bfd0e5f3131b959a7a92ff10a5fa5d70397d8a37ffc7e39a3e1af783c929f230cbf0a2708b01cbf86aa234a99190208f3c8b2b5b837d2fa42423f23744699d097fe1e45905a4c11b6ce217c2903c8ce15c4ab8f5a3d2e9abcc116a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7804c5f28f8b6fcd43777a08d0e7cb31a412626d054fd45cbef505f9b15d48d4af688b06da3b9b9a0f961b7b0db31b5a4e8fc87fdf342952ac94365d650fcbd2894afaf1e00719e007cefb34cab749d6d252574ca2a11af0c90811d2c2ec1e9f4203a5352322c48c7977e9db62e448239;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf8e1836c39face01c3942cc05328b4d7f723de7eca0d06cbf368f3ce560b5d0e59c07017a049f14afd65ac93bbab806483ae6fb0192c3f88303647ed08ce17ea648f925dda93841b2fc980cb11feaac854905bcb5a0ab701ebc70e034c49eed706ec3961bf9cbc2b9dc9ef6575875131;
        #1
        $finish();
    end
endmodule
