module testbench();
    reg [10:0] src0;
    reg [10:0] src1;
    reg [10:0] src2;
    reg [10:0] src3;
    reg [10:0] src4;
    reg [10:0] src5;
    reg [10:0] src6;
    reg [10:0] src7;
    reg [10:0] src8;
    reg [10:0] src9;
    reg [10:0] src10;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [14:0] srcsum;
    wire [14:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190faba9874e24ce7c285a8db6f5f76;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ed86cf667ec7f69f143f8c4704d6b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h506cd4977a2edc97902d8694dcf0ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d1ef46bec0b6fb5deff135294097a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134947104f6b15f781122256e16956c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee7e08c51ee36fa22c5b3f1703d82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd872f81ca22c0b47f2a8f73ae7e07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb9886b686982e354501853c85bb59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h146ab8762d6c57cee009071bd3653c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha67243ea9a38f737cb3d57616fa770;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb69fbc60e852334c4a8cd399852ab7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1e1af15fb556c66592a17dee26f9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28259e41a4b1af1764d478972e3fca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102e75e5a900e92227d79350217e281;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2b45495b07f200147fad348898e2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6dab6a42894b5abfe1af7d5605654;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff85def006ae3fc5f511f9fa7f1e92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb729a094860d71dc2b1d847cec4116;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e352a0ed3da6cc4e4485bcb179bc7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f3ab6bd90792c1abcd37b7fd700c32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h742cb92935287e43a79bc0a83ad65;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cccc4130d6d087b7aa73917c1e6ad7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8335847667af4300455378857376a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c17c59f600b66fce8050a6f8b35202;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1633c88977a6a1be22ef2b64382393f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3bd4b3e489ddf1eaa6fcda6ccc4d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8da4edbae38eb61db3b4f57b212504;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb14e8e7bf1651e5e465f11d13f575;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e3de47f3ff89a69a04ddad341137f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66ed5c6acbc970eaf8c816c86512b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h685ae53939d4b5a0cbbc3732d7db82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha35b3382ce692ab2bd50f46c1ecf57;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2a76d19be8ac5b25db01da9587e87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd33f64278f8ce97514887125434226;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f16624fda7d9c12356525a67d1c48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193c6c22c5d40d408a0bb4657a8dada;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ed16a56173bbdbcb9fd8f0d631205;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1babd68c89833d63c4399c8d0be5170;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3938e61d74ef33af1c98588a5d790;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13704ce880c9548667381c3dfd6255e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd13a7ea7342c073bdb671068cbf7f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63ec641a872d0a394c73fba34ddf5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5a4484f5c5d60429f606532936256;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4bbd90dbe14c5b6e6a5de94b251f43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f73371529c57443ec43892a1e680df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19375939ecb5556a988a53668dbbf66;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1abc07237094137ebe0d8099f6061f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc2835c98e53028f5797c032f9fba0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65b8577d1f75eb2f92f281f9545fe2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162a3e3aa48a97b0cc27d0a9b8fa0f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f725f8431053799c584c9643e3e5f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df8b3f6f7b0ac08917e11a151051f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4c80ee202e568cd8c04dff6999425;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1355500826922dd033303be0074b761;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc806722350e3667d4426d9ddcf5dd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d7a0657feecfbc7df921181ad95f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h676b371eea73739799c9f27a35501;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1194628bcf70e348afb85e8dccde048;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2cf71ae756078077d89e7fc4eabeec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h595341c4f51a0a5456f690b5b8646a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h74b7f2dc96ba46fe5892c3916eb595;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc23a800af8533fe1dfa159ba455c75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6fb022f5fc87df8310efd415748c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h673797070a0adaca9974f3d71b6a03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6682e8e4668545f521f880f0ddf42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f3962fc55c9ad9dd89b206564df55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144937aa3111b584fce9070e9b613c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3549a49b5b659b8c06f8c294a157af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be4ae771015a8ae250220313f10d51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd38011f7482aa6f1148d7771d08ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ee9fad0a191635fe582e74a57ee18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc89f981df3b7fb0e5f6c0c900850ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1876d346ee987a7a3c605766fab6424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1146668e94858e48c24227a99c179c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef478e07e64603259286c8b0c3305e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e41d3e4536928e36438b2b45bf938;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179a50fcd02ab017656ccecfbdc37b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b741df45f476179b6f716eccf65a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e6ecea0706865215cb7c20e1fa9906;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a0826fa856821c725407518c46352;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ef6e433add9a8475d8856d01effc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121f4903913dc91b0c99c1066458b56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ec85c817556a65bce4fdba00fd035;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34c4f94cd30039f6a9587038c2e79f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf91440ae3a05c8e54b62cf4225f8f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b6c8dde73aad810b1d01f01893136;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8761c3b2a34fe16bb0bc0d9ffe89f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had10a863f5c28b50dabaa230d3387;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17dfd23304f623ef96a686f7fa47eed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174c5fc4f8a8d53afa25eef6ac02295;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h481bf95a0ce5c046b88ad4023d915c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a007ff412530a649bce28980dd830;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e5c0ce21f15a62a42d9ccdea1372a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f8bba8bd91abfcdbe82cfca04eff4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea9cfb8c56e4e7e7b62a4af79612b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d7eef48fc4fb7b25ffed3da072ed1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2122c0c5d1b52e947330be63733826;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h97e3c906643f40aa4e0b8b5f44441d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6865167bc3d9bb09368a78a7428329;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h38426ddba7acab91b194a0dda8e9e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26319f8fca41009df7507ea40d1bc2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h119ce46864dd05ac71896904f6c254a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac817e2db7162c94f8874082f4ac0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6954866ecb77533ed56465534a7ceb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b688af6e34d12352e70d119807f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83fa286be322a165e32a897db3ff82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76f346df7b48ea2fd235e390e4d984;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h402208b35c066fc8d65113f5dd1c3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92498c9d8b94e9afcba8073c78be3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ca2d10e5ad6c60d4308c45f77d400;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45c64f93bee7706f371bae5b288fae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8887a86974a7b7c026c81f8b1d11b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbff1bf4128f57a15081ae2dd3b0b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha704ad4404424d54f9d71f33d2c8bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h862e088ea1462b0fdb010917921541;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1507f433ffde75e289c6c3d693440ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1738932595c9a66c13b252f8faf4cfd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haaedfd1a088eaf12959c1593b3e849;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h689241774f533121726f1ee9d47d59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h914f2805727abca4134b406619e414;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11423f90f7f1c795f9048a1ad0f9b27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a8057ef95657c7733795ca19cce94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d8e6b8e5fa07bbc4141331c53f385;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf45d5cd11d175a4627117c83f1f2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1851345357e0ab29581222ce7a39717;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9aeb59b31a1e33c3c852360eaadaf6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h949744c3543100b3f9a013c183cd91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b0235afe29a73b6319721137dd774;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e204d936e7be22a525cfe163d9d25d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf1c924fa268c6d46806983b0a29bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6dec0b50a1e7ad4f76ebf10798406;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c254c51bbd849ff41082a2853dbfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11e996652e77f398e3ddb0a930da266;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fe5ca0ea25b135f11436f34450714;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153e317143471a48d3b3cae4223cc5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36d607c44474dc3c96cb821a12a3dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4754e29e5b2e9f4abb108d1d46b2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75fb15a9d6feda97b945fecdfa7d70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b756bbf912442aa27e2713e0069586;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc962cf4372b8b54882fcd5deff30be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e6983ed9d8c4d346803c6a0ec1080;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f280a7c6e1f88811681c83fa84619;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a7cbd876712f6f8efb2926f535b2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c49cbe4321d392758ca194099f5eec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6b4f62d7b19771f84b41dfe26bf6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6fa4f25b965be9b4606dc3fbca4f61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c0b8a1f493ff7a682025bdf613b3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1000582323204c86d83948459bf029d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf63885900f3d6e4710035a39e532f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd1a30ebae0cd3b7c418aaec515b86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1626413045900e76fa016880366e296;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91a1d9cf59343cb619a1b097b8a1ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hccb01e292d27911b113ee99e38d127;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c55fe28fe25dfd61f2827fdf52a2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69d0ddf343698b49ecae43174a5d4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111e0bdbc023a79b0539babfada40e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf9353190fd4402ed63d32148bc7b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14fed97105081d7eb0549e0b98cc61a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58fa0de896093a267525a4c58ec45b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fb772e21b3939eab7a6644e84d23a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha55c4323550b0bf4b605062173fb60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f6af474a9e41f701eabafbf901315;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b431996450764386b42dc8b27b78a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8be8be3b915265f6b679a88f5d397e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he92e6b91bd0589cb4b29aa559b35c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb233c2727a375a87e96cd93c2158f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h476ac53eb6831813674e09c75326c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c3adf7db0e08f3a83f2174cf15fbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed1cd201abfb50b89c94f4115bd1cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b0b306d90d5dab91a9051fbde3808;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8bc01fc4edec4062c197466cc38c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16981921ef9a56f23af202cbfd8d3d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6a64c0fb429a519025901b999482d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2399529274955b28b43ae354eae5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc636a13b70d28680c7c9a1aeaff63d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb48f33bc9fcdf391ce4a69db2b3ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he51064ba41d9007010e6da9d22472e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8cdb63c68cca502311cdfd7c28d409;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb4e662dd3747fdbfb801bd1e86029;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db7c6ac7cf53588b64b350a2f1f9d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb672fdfc82f0194b3599c6705844e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h690a3e1b8a39649d08d4e43238411;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec27bd0780ead23701ba6ce61c6d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81043e9eef9f277ea206436fb67324;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h165757c9137d7bedc4e729dcc787b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd428a0e02e0ac537b743e22a77cc15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d42cc180cab44f70aace48789d050c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1756a374c2d37eeb93f7dd3a94a7eed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180672099a64a4bbc7d8f8e3aa47d21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d578fb8d23d8ab5fb272e77df565;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63131f85d14bef8fc27c482b2cacd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34f49a1a3ad83aa1d0f6d87aa5a08c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf120e17feef08e4c18d96564a364d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167192d9c3a9edf2ac6db20fb1a9145;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc98af3d07791c1824498ffa3c2fbeb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c9b63f16736318642d08b42186a05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd33c40511ac4a9e62df1b9be29f56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff29b3407fedac7a96a820be13435f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d519743d2dc4ec9a8333ae26a0c544;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a4b47985d32a4812f41d80255ac55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3824f1794c6d2cc68ff8378cc876e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ebe1142ef05a052ced960df3704ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8041c6eddacc749a05bda8eb984d60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8ed49a87c9f5a0335a57a7ecb9255;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181cbeccb6edc2ad28284ec317d2260;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e537a652aead3cbd94038ece30eef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f76a571b56525e46270c81fd5433;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a105feda11bb8f168c7dace1a4ec59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e78c62743c13f1bdde0d7d1129ebd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c852071a34eb92f528ff6b551fe837;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc576b70859efaf2fd1890ee07cfa15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87faceb923453ccb1c1bd13e41ed02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h322e6a17a4fd3e115fb9bdddb9a17f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h165fde768ade9b848b5a23e9a4eef32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16857226b6733582f6069e62ce4ccb9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15445528ecbe9a43a707a8809fdbfc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60bd514720d353e7c72a9198337406;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbbc0a2a8369444ff0ce127a936053;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8dd40f765b1239b3de6574afcaf370;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b87ed0d090e5663a068fcb88910de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50c7ef2f312f41fc5792ec693a8bf1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4e1c4f51e03c9640f9070166a24e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57db32d1f9c01ff0ca59ddf6d0e9e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d240391ea7ed5284d3fe826039ae5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12fff4f580d4cbd5f7618a9dddaf85c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b2b4a776f0e79696006a68c94a5a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf44f6b0a01f27dd7ad0d9c04581ce6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcab4bee656a584e5021b789cfd3a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f54d06ac2424debb5c6cd7de1b0dd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ecc4e3a852952153a8ac4d39911e9b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4abb4bd6b20f53eb39f7db43527423;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54c1ef2f72dc243bbc08daf808d469;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b1612c63bf87aaa600c4ce0a0edcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8448e8533ff17c57738f82a363e1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9222ae107c8abc50bfb842e254ce9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14dcbbf83edaa23dc945da56e8770b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc4471dd1113a1d82b183f0053fc1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9589bb5cbc82e264f0874dc6f780a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9eb2dc7361aa2637dcae9b0f4fce7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eeb753583860a4b2940e27ad742f2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h738e887a43ac43bd53a04fdc44926;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108d7eeecb6ba3254ad6c44a6673b31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0e1bf6cad13236cb9c0d545760491;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2baeb8212b4c598a073d8907da3a4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfba58c4f4a1e62deb2ac806998a3a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b292ce92c45b7e33499692c16f445;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba09a60e59ee448cc8abe898f04024;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d40dc18205a0ad6a07fc498d5f4ffe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147bcfad82b90ae0c648a6f43df94a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4c184c501bb507fc5f2acded823cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118e7491fbf89378b0009ba6c0c44ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce982438334153962c648bff107b32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10990571cdb1255bdbba587391fd8b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2a4fb58a8db7f6c28bb2e53a1b195;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164624287e78db00060b3cf1f7eddc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9449c197f255382a2724ff4c5a4889;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13006221217962bd5d6a683cc131443;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87a5f1fa660a5c7f3ff6d836f5ca44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h122e5622c16efdd337b8c744ed4fed8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he9f9cf7914f0c03248ee37b72e2dfd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24b7ec1ca88eec76cea4ea71f281da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb7d39cabdbe39a49ef9b206187426;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1242bbcfbab77802dbf08ba7a10efe0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4c38c2c988687447da04860e90d2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa67a5e5001d3112a2921407bbcec4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha59a7b3abbc9e7f6dcc81166a14494;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1731b27d540ea4c72a7ab50025b6360;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf86241ef051efb8f31d512ca26591;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7499dbce60091cc1d09d73fa8ca239;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140f0e856f1dff112d40a2f07b3db26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d19d55914c1594429892abb3b1ae4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae49232306a8ce6cf3fb9616591c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6cd29395829fddd369f056284b168;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69b757d9478d7574bf407a11a200b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h537262b3cf0fe0c5fc37b945da8682;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd138834848bf5218b355155568c7e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c523ab16e7f907a546d732ba4c41be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd1fcaf65d8031e7497d9bf8f44224;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187f0083d9abb38a41a6e12818f0caa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130f39429c1adb0806883bfacacfd4f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5f20c31972c60283e84cfc1f75a28;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44ad323d17ec2710dfafbec0e15447;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd237be784dcae6aca33cb84feee272;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bf34cdc718ee2bcd53604a85c819e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadad0ef6e59bd3f6fd669996f094d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184e5dd7519cb409cbbbd84537c9861;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf62cff236b65f231d87879f4f25f72;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42e102b498d5353cfee27e174f85a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121318c146a52e1f314ae45693aee9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e21884ab651b7a56c303489328cbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1420a9f6e4a5c2c8f61de12a26b5626;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h741c56d807feb977cd8159c1d3a02b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9b07fb703dfe910dae050b5e8ee8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb770bb5c22bf6130446b2b581ff9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc375b99974bd2745c40569c68bc35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c363510c78dfef17423b8ccb5f885;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd02afd876c92541e922797c968d2ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f01e9757c2729cd1a984a98002099;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160a901e3bd42828fbc7507de5ec43c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea0abb5db06eb94f2a09a15b7a6673;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad186528aaf6823e1b2ed309387b80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b09ad67b558057978cc038aa353cbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144d86abd2d1abe660434a57c98a7e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6377205185a27376ff4f0db56705e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha1c6886b951ab70027d8f36f5f0c4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1417c91d56bf5db2db7c94ad8793203;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha160e5a72e688f3ed58f1ca7cb4b1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b74f0ab747ed8d687f3732c42df51b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118aaa32554df3512360bde8858441b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf13f1c975fe3a50eeb86a32bb5251;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c2b3e1a793454215c858c509ce4090;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124969b16c25d3003437e83c372283a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2d60f1524743a0b60c59f36bfb366;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc496b611984c4211a136c6deed668a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109c96b648e7b635c39c28772813443;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h104868ba9ac10b9625a988a66b80c52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68c2b22ce737aa05aa08949589021c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e783e0c85c3f83935b0bfb4f5eb02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h104e315ebdbe9c07b7e497c3c9e7ba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c6ae13c10139ad11b467096e743ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b1df225cc79efe9771185b84d3471;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h798c30082d7f3d2b39a6b5140454c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1040838d581c3929eb4830c7b4855be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d36b27e191fb9fc977aec9a0cf113b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0436a755567ebb88c26be8f8ca4da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1897b7a3999b7e5e65efe9d2ae2a64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ab309dedbe581297e22edc13448be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192e58bf630a7948bcb79ff6696ca02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1633bf23a3669a741833c350845b9cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4822fafe2ff214376e91825da62549;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb60d125a26f33df625cb0818f53717;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1419afccd1d4e708998e5e25ec432e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173ccb05452d1de8a85bd8090a932a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c7449ea48c269c01e3935eb302583;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d6b46650bede1aa989bc8cd2b2e7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b833ad93353d614211f37a57082eea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9283b04e4e3658c6f0b7dcb436395;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aba938e76ccf14d0c1cd61004a114c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1feba7d0ec3f083917e04002f52e4ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c800a110636117ab691352726d4a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h540926b6c4f32dd8cccdf8f8e9ed32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1255b138d4823ebe0237c18bd2e15a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6762421a1792946081e4ec871566d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h873dee9eac385b298d265381dfbc0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he88515d15a2a075a4dc2e4df81dd4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa849b5bfa3679ae8cde36761f8dbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2b13068642d0848fc87af0314c4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe344bdf3c22f92c2db58c9ed8683;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35fba468b97f970d254d7f3409f7b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f82ae12288e9894a3e7a3713504a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b40d9ffe04469d7feaf7d5a69f60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19cfc58dd718279ffee955e216eefd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58737e542c8e21c897ad5e21d0c4b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f46efd705ce201cfdcfa999c7002c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124afd22e04cff7e261bb14c8d00d0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h55184ffdf96c0d09333ac09b4db950;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a8079cca10814b1d39b357e3594cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc57a2b140b00b42cc609eddaac1c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb34fefbd70f086fdfa509a41e25d54;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he26e1d8a87fac7faafe87b32ea8755;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2925bca3c9b10d418ab49733a31e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72c0e774d15df8bff6b5cd8763da78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39d29c13e31aff42106d8b50f741b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16eab28418b2be848dc4d720ca8a78d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f925bd0954b7b428147fd2dcc24d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1bc25c34590660c5d0d426087e0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba54f52b8d3a0dcd4e4b2ce8b708f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cee06ed9d148898b543af84bf541f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3cae891bbe9f4eaa0d5f704555376b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d041277e4d0716351c2ee626e7e25;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efa5ec5e2d948132663f74082a7c9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbe78ac135cec212113715200a2c46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1d011a6145c768f71eb230e23e309;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163c5f6aa6cf0f523ff297374336754;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd322566ba269a91696abc6373a8f2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75899ba508c8fbc7ad278ca7bdab2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db44a8d0345a8e53e7ce081762adbd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffeb1b99dfe711f934e081d7dd29b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d79724bbda8c9d4185f470d15a9d45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1e395911a02d6da99592cbaeafe99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76f5833da80e3b2dbf52a6cb65bd74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha191cdd4ca9a4948b81cdca48e6c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155bf863924b0675225a56b29c30922;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5611cfb28fa175da60fd9ae8d21444;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ce468ae1b030b4e2e521f902e116f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171d212e48b2d6d1431ac3bd3f7ac67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he77f3214e8b0743cb786b221c18571;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f32392c5d9c1bca57f4fc78607838;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfdb4f5244dfc9636bf067b81e145cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fef6b2e922aebc6010a15d80f35310;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f36c81b8bba5779d1038e3c123ec7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6fa49924c8902de484612af34ddbcc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36b987bd4332b66ba7efad2ca30f41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1f1a64d8703a59d3e0b1e5a212a42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb62b4f5144c613215e3af6f1276d6e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92740a2e9d783d5d5d6d77ddfcc128;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53897ec2345e182ddb66374b0f706c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2904459ba78a34dad987afa5f1174;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8bd1afeed7e0e6e706b2939eaea43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd90978cd6f34617e48b29d58311dcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b4f8f147c75eaa11c4e72c5e3aecfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb22a917ac45228f5847e3eaf2030f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf208e7e4c7b410549cc70cf85f8443;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5f1736029f8a04c9435c38592d7c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1fb8ea43f6010184b27b673ee1548;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13abe71c4bcf16209586ca459e68e3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13559c13326dde175b40bf717ca28;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e3402e22878ad1f3ee5d6c60f1919;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h610c5a3723c645d382d3b7761f4a3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1b0401b421246310f09fbe00c7d5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1743dc2ccb087e8634dd547f2bfbe5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10033cc60f441fd9ea557ca7cd837c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1dd68b9a4c677d979891120e2caf6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f65ee6ad2eef0e9644d6740cf9fc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86edb9cf1dcbff302ae4f9f142735f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f41cd27a5ec4f7b8bafc589802a63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86a011393dee9611898665880f8c5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4583d82f1a251c01ccdd6f3896c18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1348567198e730a31d7bb687478efbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2088201dd078bde01cd15669bf16b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8bd081e637383076c82210316afb85;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c351da85cbf50f3a25f25f7bb846d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c47805aa239786ea5c9d3212f1a2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1367bba6f6aff7694bdd83ed840fceb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5eb3b59da0833bedd4b75d87a0b69;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h825a30aa8e5b118077ed212441a3ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56339537c6ece95a60599623fb3f4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fe0ae10d445f31cd95805e150c304;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14fa60a09dc48f891d1f8796a948bb4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e647ebbd8b8df24e057e61491c8c61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123a3d68a0366e8ee9a12bfb2690f2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d2f73a69d560674126cbda826b205;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1964527b3a0f57b2586647a7e3ecc9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea853ad6bfc3c8d17e88a1c9b4e976;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee1ac5c9eeea31bd397acacdf044e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e560ac6c2b10aa78e1e56607f3d298;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb63a55242f30835b5e39d7dbec21f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b065cc556cd2415acbc24533c0b306;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dda869ebc199d4e84a7d46fb753237;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157dbaea0678177ac1a0cc3a68c730;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11630d361c596697f63a33d0240f0a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffcc3ef27dd2bb35b818000e04668a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c440793a7a151758ea09bbe99127f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf173ba707d8775ac80dfeb80a9fbd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110f55adfb940ce4a2401097b489540;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb19c1efcebecf6cb418f13c288266;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cff58c86344a171944c7bf07576a04;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae4944a727f0cd34e0ba376802bde2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd33197f2c7d840698744b1d4a01483;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1151432e4ec63107447333cb76318f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9269e9c65d3088c8e772411383097;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ccf489b623743d9a8348a3f55c9fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19627b7686e93219fa71ac860d0402c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce68f9973d9eb501e4c62bffa9af92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fac9348390e5eeaa0d7942ac8ca195;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16bc54b4e9d6544f00cf1d22d8b0e5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h122f61213bbf336e73d7cc2d547e1ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3ce9e364e4f167b3b52302559a623;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc334a7db063d8f7144eefcd4934f16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59bbc7fd75cf2c31d7117325d330d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'habf98e0b7d3b30b888e21ca962fee3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4d578d0c725a416931e034119e22b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7475543e9426c4274eb09c9596be6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b3f6d9b1990ac66f04189c5595cd7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ebb8e5bec085e0a7a1a9173a35b6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a1d57aa23c7f243178869329640b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ec7ef19bfcdca9d7d5d26e9074729;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1708dd311d8b41a464f853f6b379bc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdad3ef4482d2b2e20cb99dae20c77e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179f8cd1e31974f96f55f6984e9be6e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha75da4d7b8c4baef6b8423a48c4f07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10bac761e103e0d65cf655a6770febe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163a40d387148cf4dd009f4125aa056;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0677b59661fbff2826c58931115d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184f8c9ad4e4c8ea104bc30159eb668;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1810ada6d5a7dedcc76bd57f49a8949;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16720b69786f2a838ea1d355f3984c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b221455724ac6ab332b4984fbc559;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb4d68be9d4244e858879aef94c6e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h20e42adfccd54285787bf63b9bee40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfec9ef43eda77e8e8ec07587b0d96e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df85bd3ad324a727e0598e30aa01f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf4b160a26f6345df3020cd4aa3258;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h811218d43904dc2231729936666e87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d124e0a7d78d90bcb2fff8bd3cd47d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28716fa0f23b0312d23c8753acfd01;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105fb8c4adde1326d974784c4b23df7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140d603d46b6e7e5539186ae52c145b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda46a89b3e0f59e777cc31fd0bc509;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1985f27dffb1f966e95927d1cfe85b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a64b6cbffff92833642d14c1649f5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39cac20ac8f85d421ffe3964a74c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h185238fa1bf196cf90b91e2b75ede5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17073ce28662e380ebd7ef292d0e4b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f715f781bf4fcd53295c2314442dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7b38f84f8437c5eec7368679ad4f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de33b3971fd70233886c2632c64d9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h750e2e30e81dbc650bd936bd0427a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h137080544d534b2b3dbc681b58e79aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he18ebaa9ad032855ff804667133098;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1547b511c1a7af9a60c2691438deea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a01f3d9b646eed34945a2f35f9aeb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d788a1067d98d9d929f8685c18df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6e9db38741b49471ed91bba5c089d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e6bca4456e3435cce1704e5b7e189;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145a4cfc42d300443745a2f7cf587ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73b946f197643390a9129f1828214e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd673fd383833294252c938d76fb14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1690de62e55318685d117e16b025288;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c3faf9c21c2bfff533d587edd66e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d5cbec6dc424f0ba0d44115c4cdc6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19539c6631379416728c997201d3183;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a59ec72ca6aaa0af2e3ec4aea6f52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h150b1dcccee9d810d35f6593a5f0def;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3d7371a864d3858dd1d7832c28dc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf0f41cd3964d7148726eb13a5af4f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a214570ba8f1baa6bd3b1426ccf99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c29d5d327ae8f5f51c36abaef2e6db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e88aa981b90fad4206b4277c7bebd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143e105e6496240aaa43459864df9a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf866aaf06cb6bfc3d9b0222bc85b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d373fa77004fd1dd70b69f1a271a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b78314bcad455e9a044e875e0a8361;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f0b85895fae3efc100e625d58c284;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d12728d1b02202e147b2ea7a513cd4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h630245c98168df495fdb805b100cac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4ba412bcdfdab9e2d5136b864a8dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153a9ac3873c11befa04f1c2f4a93a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdede3db6e643d2add71a706a5aee43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10206d21541d412e2cf6915b83cc20e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h972f53b87557ceeae25728a2789c91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c905edce5c6bcae0fa37fd7aa3ba2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14aa0f14a70f3d9b7f7b2ea02c3c0e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a0dc3ebafa6965e3cf96de9bacd93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d8a3f0e91b7d972d5e77125dd61d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a0447b6a6239294c62ded99a81767;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ba98535c382ac4ce0e4f4e8ce75ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15deabe70ac255687ca7b3f3487a59c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h560ae774027408c3da07b083a9bb16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59ca89ebf4a3e0e5513ba7eba91ad0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135bf4d4169f0e8a18a6afbe75fabb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc754471ca12c108fbabf9f95479534;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15924570792e091a6f64d64a1778f8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5bea3bcd6d43b1336881b97661839;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11182f38bd2a604f945a5fb2a777fe1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0a0d18a1c30fa44c333e6fb5215f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f41a4d2d9dacad19fc86fd62159ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b152ebfddcde0146a8d36d235ebd1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45f3eb2cd507f56bcaf6b35e730be1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc57e2e4a50c82fa0a9b59a403b4fd7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd87926e85edbfab927378b181b023;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d5c40a5a9f9ee920f81b7b1c54d4f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbdc3135d44e40a38d1afbe09b4d509;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h504a5b0f4eddb0bd410dd3b59e907b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff2bd2d99b092b985badc4bbc7350e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d259cf4715f8df2c7ef4b1c237efdb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9dbe65b47d4d1e1550af27b9779f5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bb14d49a11683b133c10a27b6be0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6207f249e918f486a27870152acf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92afe43de29be7b7d24a2f969152b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dcdb6da3650d8de96b4ed47e026d32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19315cb41da842d24da14f4a7971b0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a184d3b659a2f33a72e97aa614c72a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa5b82ad400362afb50e3e9079074f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1776ce7b2c8308d1ebd18408f6b1a3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7f428c115a6cd7e2520ad7551329f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h682c5e3b53d204dbae87659d2b2e45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5635abae1ea365946dcac08a7605a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0b21d3c4c7313441d581359f65977;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e976c4e76a4350a6a64f687ec77cef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18530bf5dba0b7a038d097a8b41bca0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h177f50389f23307d91463d98e7145e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb9a0fbd2283b845319acadbaf7d5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14220ed04b471afd723d7dfcc06a7b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf52d4ee7645d8b750ad08d32ca4ca4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f76459124cc1380ad29c932286652;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b61538efe6801d31a64cfed54baba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cc653e5dff7410b631ad25c8dddfab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd4c89b475fea85c78a13c2acc1dab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h529296ccda3ff8d18b18ebee1b9a0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c63a55daf0cbd93644e52f6afd6f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h154e04e81c27e2fc1b73f81c8ac9574;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f7dc016148e6f8fbd357525422428;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ba8ea8d0b2f25825098da0f26ea56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2af95e4f2e51ad8046128845d358ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe17a2731230ad8c335f6bd8d95832;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7974d12f0bc78502a830201c5161f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hca70e16c5a286ed856815f5fa35879;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33053016edd837afced45ecd39f67e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9026aa77f2467afb193ab33c19556;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113f1da44797de638aa6f38757657d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1105e92f0b56c9be897faedaee1b64d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1799b8e159b018d534c9135ec4f49d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a686996b213a3da7228248ada6e1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb890552999c57fad9f6806d663791;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f32d447422d93fbd8481610204074;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168dbdcfc35dd05fbcd9c753d6efccf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b118ea570a0288488a99d3bee6ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ac8e194225ade0749a95ac3aa80cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9e372b48aefa42062a0740d3f5fa8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f02d364362a65d1fce01d37971b705;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h294291c79c1c905cefbd2fb771b499;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c34b4edce4060d080ea66612f77326;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d71115c451b71e1afe4feabb7fb93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e2b156d49790254d511a39f5895f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he83f8daeda9c1f061a4748bf0a99aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af9a0a7396d0665df4e68b2303a3c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1beb46b32b832f23fdd79d7a14baabb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc800e4c829d0d0b0026632fffc962f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156a223a990332bfa73a8d61ddc4bf3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9eb726a141248193180b3af000ff4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cea4b060daea49de4d3403207bfe4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120b051dcefe959d01a0172719f59bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db886278bf7821c4d87f506bedb0ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159902177f270a0068cd2119a4a0d88;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5602cd6bae3402ebf5b7e712be74e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3586343166f0c58cb7f681d2a462f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h939122742bd9f48270e1770a463b76;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111ae73b4cc9ce73103ce2703b876b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heea6d64f42ba3d1a4f48c37cdc93c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb8659c2cd3574ec583f2e2f844cf2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2deba8b362f2dd1ba28265960544a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1129549363aaf79ffe65b20b0d7b5ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c8c8177af7299c03973cb547e28f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dc423a8b86ee3e1f270cee028c2e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ac5f9d54b50c3d9a653a8ebf0083;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8838f237fe6e98e7c2fc9950a5172;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea4756cd6b9db3c206b77df96439a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2ed47ba6438338a67d75d67b7409c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda713c8a38adb0701febafee1f741;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a1be80bf03113ad7c266c5b42c15e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdcc119355698bc44a318e5b979a217;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d40184b1de0c7821aa8e89f3f0814;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1f4013c85a50d4159b6394a31f93a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191d906bda4ff47ef4f9b6369820e30;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45fea1428906735751ba7e51247696;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a0cc5ae522128fab2c4ff478a6ad3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h302e7fee44ac52cbfb4ef5ed106e10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18417d7e9580c193b229645f8700453;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1373265e5a832e592f2b3bb340b2a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ff68c7416714d694738319e2f8edb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89dea7d25258185a516c510d8be42f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc86ac17d4ee3ce1d14fb8d925ad894;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f25f7bce36e34236c9a2dbaa3ad819;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a007d63d5bf3c39a91b54d2ed0116;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65a76329c27ce2fdf13226e544cbf5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1afda274195ec1919a44f399135dcb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef1861922194788a7c9c6a1e9229cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ddf3e92c0a6cffb8728d1536922a29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ff6ed51cfa10922808b68c6394b13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1546ba5f24c8eb26e5a4c366bac902b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4f2605e9498d59a951ffb5621558f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c74df63236fbbfed2f9d5ca49d3c5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbd0f8a79ea7d4a16c6461fd95dabf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cef08d8bf4b61dedd45c0c84a45235;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f1d4bd5342416ee62dda8d5bca349;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h351fed909a1fc6887f94974ecf1f70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8920b235638bc0217665dfd0630850;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8eab72574ce1ae92ed946fa7e8c8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1460698778f626f4aa377a2516b5d2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7388230b2551c8c2daa993cd940694;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b8266e8a4b68f3db29291612ee4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a20dd6151cbd68e51cf0e37d0d64a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a87d3439956f8d4e4cf73337b974cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h259007764c50d7cf49d948f942d6e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4744636a86eea784f0d9837991f9b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2cb0418a96fd4ab955b4f2c6f94a46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f914631c63a0b1eb82846c24e471c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141fa60bf8b9d3c92b812ad322d40d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee5159e34e5104b99c91f9c24acb98;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158ca7f5b2224636ef07ded934030d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173530e6921adff7429224b23d15188;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f3455c17211796931462d526d02d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f04d773f6fbaf017be8a5e5734f7c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e55ca48dc5b2341215b0b4e991996;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ca664d2d38b2807ccb54d13c21925;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11185511c3b15a239dff4ecbd55b0ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180e3923e5cfe08472fdf878c3510d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1790e16ee7a103fc61283c09c93fd82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcfda08c6167390b15c52a4e0967aaf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e3813c546c0a1258ed44d3bcce43f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8e78b2274a4b27cfd51ae2b8928e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197eed18604d3648ff0d80339386d20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196285b82e3a81a754de07d6396ae20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3bf9d4a956c607ea508574cc86fdf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98bd952373feb14a07b5fa7b534cb1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152133383fcfc8623bc6f8504f6a9cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108ee68f60b0b89d030136a7a0c4bbe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h219ff1b153bf913837be2196c4193b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c06a722125e0f39f86843c1fdfea4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1794815a0efc8a9e970527625b95998;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h373ef9f51e533359b794096d08bf2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e510ad22f16bdf4a65aae402f579ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182fe34e2fe991dbc8304afe6019aa2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107bf199ae2d79ef7ca74a58bdb5c47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8aab2ed36a698b1e2ed8ddccfd61a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h569519af6bd68edb2776514e8887ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e4a97b060d1031db1b6b12f9eeff3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha38713d183564a5c98cf1453932db7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84e5ba900a0c562ec7847f85279367;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce8805fdfc8f0f33fc5aedf6f9bb8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf62adf96c6027ec44b370635e6d845;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfd127dc81bb340f8adbff48f80a40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102f00495d9643f5528334d9602d0fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h577d48bbd3404d8a72b1498c8b9554;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f8e59ab0cdd9b8c219e0d416742e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9538027def42e7f7e55d14f7747520;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191d12ed99e3bcde534da2f3bf7b8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11932478a2439ef7339d061bf20263e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98c1a5ffef2f92c5edf93f5343961b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h268e113a98eff72153b97891d67d7e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3c27d696c330ec7b5865a8f74376b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84f26f3a83b10560d15202be296196;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d174d14d332dedbf3caf1f921306e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75aa58ba547927ac57b33d6f9325bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14df95f7aa0a675c7bb30fb7fc3ef1b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c93915bf3bb39b973dc05c35632707;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de9404020cd3fa80c0f2869ae586e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e585ce71107a86e568cdbc247aff6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c37b2b7dbccbff27d399f13b3ffee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h715cb408e5ef79133349c959b87f6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffdb8c4efe2f705876a31203bca2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h646a7d454af7f6bef5c748d78bc5d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa71e47816266abe62a658885adb94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118010125b0b1392b9c9d3270d89258;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141d8315fbdebbbff71ffcb72f317d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dee7a8a485d6454a5ad4d06007917;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dbeabb919b1e5f0faacd4be32d1d93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6f3c0f61ed1a25e1efe4de261320a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ecb5eb6a2c7a93c38dd94e0fae9cfe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181c72e6f39b44e36ed12f62f3aa782;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15adde9192b834863e40174680562f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91df835e6e562e648d021398f0ccda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128c79f2514ed020f845f91e8713ec0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1834d2a015f58bc9b84d9f236871a03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92c68610ea3b94c5bec5d7b6f7e701;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bd690a502fcbe843423077544109a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a49565885ada36cfc24a8b9d26d5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h706b54a722198e4b8dcc5a60ab2006;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4afdc63f0ca67af5849f661e9b64c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4275e084672c902f692bcaad2ab7e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45e1f0c491db0af83859b893336abc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc44431ad4eeed900b14051829102f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba6907db3a57be0ad98e305b9f459e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc6b72de94bba96ee52de54bfbf2e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73fd7a94bcfe93ee434f296269bbcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c817783424960c48d74afb772dd22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7b3d10d41ec584e3236d13374b515;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d1bcbcee57ec91b1defafb892e6e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9984ee26f1dd040f0ca109097f246;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h427b47b543e026f210c0f004a6c997;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7418e00455d249ed9f064e02fd801;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1316e511e03c090f886b76a3840378a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h20bab939ffc82ab83b8a30ffd637bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1430369dcbe033f1f773920d9e90253;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h397d06b78a189d2482b3bfb0915ac2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115e20f6e323ff833d583b8f42ac971;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6cf65b01f4911e81e1ac9d5ddae66;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6cbc534075a7ad4618ed8d9cbc9b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h713c2f1b33d7634c068f356e9eb5a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7017f39a0ac041f75898c1185cb8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a152cb5e991d25e49b2aab411e932;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188c1b945f7b2ecc5c50a27de1d3161;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188b2bd1506aff794e772ff15c417f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130e8d2cfed73c836c5c921b1f8f350;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h734608a395b4c696b13970e4cc4d23;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49d4e01c5ac9d1556da2282a03bf0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e6d2d1a90003e3f4f66ca90ff2912;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b56254f8149c2c3d3639ef14e50f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2dc4ea9130bb8b23d3504e3e547a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be311becfe458f607732f073779091;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a809426a8ff02c858349364658a3e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129cfa11c1de43f7dca3e99d0c9f99c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c479c815ff60b3d0c376ceb69fdf1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h660b25cdd97b2cec3610ea849f6018;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26f468252c1b91df983f2841d24012;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1956a11b5a5467942911ff251b75fe2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb688c119b7e278b7f8899b6667b1f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he79752a329929eacf637830c07ce08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c0832cb75d33e181310b526614a2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbffaea0000d734d338f2163c24e025;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b5d83751d7d19a8e42991b7fcd6e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0a53a40b891fd8c7d2b49de17645c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cae34d4bb60fa0d57975d05769063;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h641379776325364d540c8a50b56de8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1151873d1989855399321b0306cd0fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1807f961b327db45b25670d1b61de48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fe0478aad28233deffe4028c80b9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13aec8208039072dbafcd1addc0565c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e17e83aeac36fd1361b7b89fb96e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b06eb9df4fcbc1c173dcef8cc239f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1e0197455aecfa382f589e9d97806;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87c774c8383d7cdbd02a3322180393;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120626d1b3c17f9011e2d5c0a56275d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f36640f2102866d2f564017a07e3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b8078d6aa693e0b464e570229c2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3dad4b65e20ff7c942039df12c64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb428ff7c29929c3aa910a2cc11f60d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fb190461b3923d11203c0d585b830;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4dab18ade84bf06001596260b03809;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d2c1185938157983fd68ca0568f55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a7bad1cafa19dd61719950eb144e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecb6549a990c03355798fe4ec484b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26e2ca83cfac5460d364625e7c54a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dbe3a7bbcfa1f445118fa3b1ad1745;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b87bfe64b5f41466f3114363e403f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1958365cd5f7d7d92e1b518f6b6af9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d04f3c4f6fe3c1db103914a67247c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a8c96b9f9bccdfe0dda723370794ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1708fb031b64b5906734b0bf804f1e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad0edde3a69b573c7401fcd95a31a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a3a8bcd5affe3b9ec86333240b798;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1060a098194d0fd217b8df151455185;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bf50a8e96e69f424f548e03a47233;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ffc0210654a58f9bfab340f7c96d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143e8124effb4e77134bc4afe5ceda3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ef4210c57a62d99a0b417d57e255d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1771844642ceabdeaae727258b577df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141eb8d5cac9a56958e4f49d53637b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h989ef6276153ea638fe03d361be18a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfc4b86813ab925e3a815e99e27db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107061f3969347db2a4f3d48e0405a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d469e30cbdcc560a339bdbe62a996;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e7e5e61406fcd99a4bacebbe6156d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7853235d8e5b1ee5b38fa6d334cb61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13928d39a4b011362a0065296de627a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108841f090c70f100010a6eb5e22b74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10750ae0d7675db7856463affed4244;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4d8c9ea59a14eccb4aa79ff89afa9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ddd35432d1c14d4c732d22dd41324;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1da7c746f7417b946232dbe007f0add;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66482098a7b47c5cc2191f5bb35b7c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cee5fd3be884deb09cc29b0af646f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4c3ae055e5de1ed46e7501491ec28;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f9f6bd6d71d8db05baf8b7e9d005e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efaa387eb5a983c16f2a69ba9ad2f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1539ec6172cc5a7953fd76168a56d50;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e2dd882c4ea7f4ea6ea1ac799444;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10c3ef921848ca06888827853a3b5ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4c89473a72bcd694afc763bcd50a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h618705f816d9b249cbe2004d6243e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2023d9955a4318c91569b896ecb16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h730e9a464645c511af3a2fa2987dd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76b2e271833ae90d1d1abc764f5db1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10106265a25a7a3e3f9bfa38c14747b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18589ac1eef97d7c59b098466752bbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e0554afad67bd75c5ffd6978d4adf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b50560a51c0fb6acfc7c83151692bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4dd44a70b94c297885e7d84459073;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28e927ad3a701d2ad070034869db3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2fd5c6efac0f933eda6e54797153e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a3631458c205f55967e2af85ceb3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dad029c2cf3a06b7b8aca037357e64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41a952fe5568b674c8ec0bcb2267bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc612a722c75f4761f7fed8cd94730a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f21331631d3c72dbcfa8ec4211abe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7e1a73fb40690c30069d17609f802;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad69b4583dac65ac06988c94ad0cc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9fb7ddbf2c2b4f150d82fa1781a5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89e7a1daa6afa9c5eb34af560c67b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed8a7fcbf33680982a43df99b7b86f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b2ad68e4d6461c3f92ae25801a207b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f3b4a783b768dbcfb61c86f50bba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9b7f4b69529b1101c20d60ba87258;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4abf4153ee9bb863c4f51ced7ad78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d9bb222e28f225179083325f4ae4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ace0be186e7a2403a3a06a2fa3301b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h571b4eec7a61932d5a40cfbddaf843;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8159be94fbbe3dda7b45da97f7a2ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c83383d017699a2ea94e34c07b6a61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c500814f01f6672f32eb2be15ab06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d385dd5b179cd26e4f1a5946cf992;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21ecf49afc701c056b1a732a634b8f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ff70c6d18586f3634d8faa8c2609f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2999d77eeb684e817cbd2e709038c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145a0f8e1f6d673e6952a5455cc1291;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dcd490a7745be3d7fc4514d952ae73;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1433838d3d68050eebf3652471ce0e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc364092a469c95c6ebac782b293f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d002c24eef754ed45c4ee37c89503;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a090569bf457e283749e37744cbc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27a292d2b511efd86384b85f313583;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b40ecce843922c9a825cf6a77b5c90;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45e83a80eb4089bbeb8e99cdd996bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ca72f966c4e2bd8cccf2949531bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1970bf8665ab5d44c842a70b26d71e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1a8bc832e2feecc81776bd7fe1c39;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha26e6b2c4cfdd70f17c4f9fdce55dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1103dae91e69072be98b206da63d9c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd408dcbae6eeea2142e2abd596d236;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bde1cc1f09a97979b7694db341e6d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a384605a964a509968de410789e63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0b3c87b25048eb23f99b8613697b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32f1fd49586f00ee3fceb54c40edcc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77fd76e8f052c27019a51978e643e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32ed64bc23b29ed2dd2c13c1ee10c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4decca3bf4988a7dfa4090bf064662;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a659b301cbef8b9b7e78bd107e38f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc67df6a22ef983ea5533e77b4a38a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf497e10bc13aef5ef449248e22542;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1410f87bab41837b1dbb0fba8d78ace;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1adc8b6c267bbec55d0038db344dc6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd17d4708db272b566d89059ca9c5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdcaa53633a29d0055fec6f90e415ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58731d42af0ae51401b7aea72810df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e6b39dff4f90a19f2be38bbc7677e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7773495aef81626209922167905e49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffaeaacb5eabd5ea0e9b93f1a04903;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90c9df8c8aa7a2014b9298d9a70535;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7ad9614047b281b22415c11f347e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha412f73e071e30360c737dc604002f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd60b23d2db529d133285d39ca7a6e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73c19fffd1e00669dbe5588f7d4c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd503b8531cd9b7fccb5d41455c69d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa35c7eb17df4a31facddc69f46a5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5aa0f68ea6471b66bca2238eda5fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb8107fba9029cbbea87235c483a09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47238314a12b02742acce52e378363;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144ed34849054da1c2ce1203a251ecd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ed782119fdc4b334f214a027a6c2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c6c8ba04dbcf1fb08dd51efceda8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1635e31862f503f16a505a8ad6aef03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112c4eb4cb7b51c2831e45e6b40ea9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h548fec1d99d5b6698ae289f8d031c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1c3c453edf1ff6c40bc03c9d36293;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42d3f17b526865de16169595cf4664;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1baef6009b5336e6f2e88e0ba6562a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h415028a5f2c4e3788eeb24d6b5fcfb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c02dc09952baa59b0c6d51e2111b58;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7230284282b3d5ebd9e51c6848837;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd34b51e8eda6b81b238586d377449;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdaa89b57494b152b75e5598d972cbd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e4ea34e204a6d5f8ec65fddaa42ffd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf0c293d08fb6c52746ad6e88ef2bc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43b5aa3bb12e5da3192f682c4a1315;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0c143a5cc7998b2856c965d98ff26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19dc86fa95df22946df8a8880152c07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h452b97963d62f59767d80a2e684b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1590d3f6533070596284b54179d7eb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19349960cb6c9a13d911ee3706c352b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f8391b62df0df3b679863ea5ccee1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc798d1e87f9019508fb407407c006d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5ce78ed39b2e28ef8122a45951f5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd7032b52c0e6506f6bffb89a38893;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbaf2b80ade94608cfb95c7aed1343;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d23285c4c5ad57a352102ccfebc69;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95e2666b1d6741bc24a780a1d8d9fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9e644367c620d1d1f7c07c98a69b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1352242bfd077326358aff5715bc71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd60c6e416a2ec47aeb4b03cf6684aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af87ceff6954d60db2863382cbdb74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dc22413f12746ec086cc3d380a4f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d27631dcd6a9c2b75399bcdda72edb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe1d74f4da66f84a6357bc0886017a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h578fcfa748fc020d7e19443b643afc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e6eb2498346e605eb4eb7553f0345;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbda1ed6020cfb92c66f22f24261efb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ee862b6e7e9f5e73ec33c95a6f14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf9556313f5703911021cc4d5721f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c285c2a10f9b6b00fc89290b2593a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ce062db6d18267cb60b02305a86e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34526f8dfe6091692e6e13236e66c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f179406fd26810208d628079c6948;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1851955c47d30601dfb13bf432d4aae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2a501d9dfa3e2b10184a6609eed7c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f2c21d1adc6a22034e6b4269f34f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d224444860a32131d86b325a95e38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1beb43014ddd1fe5f64375e44e6db8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10bad47e8ceb27885567e4549f0e6f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h442c2c84f3a3293946a8bf2095fab6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d5aa3a628a9997cfbcdc7503f89b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5c95b492831481c6f9da20598e45a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2e3f26a22af1e20fd5ffa4f6be1a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e9f784641dda9e8acf9c88fe9889a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h88a8e789cd0827caf34359265d6679;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h727b078674380b034ee539b2d51a02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f06141bac43cab32be3a4df0a0ed4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe7b6ebad5607d5538b937a1c1c592;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d895458286dd0979f65a1f4ffbb512;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1031d42baef3935f08f5ca2b1bf30ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf117e4ee13a401616b6e214ccffc22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3c13a3138d19d8d3c7dec588e49f16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f25e930bc326524aca8a91bdaba02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f6e55b6e1ec8e33a751596a2da809;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13834080b94ba2d2a4017a1a79e6e47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34bea279c361ee10c2e09d1479f27e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cec8a15c7a484d00a3b145ecb9c9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5f079885ba1d85527e8e65dfc3da8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a2ac29ab6328dd4b54b885d64f1e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h230ecb09e13c2faf54709b503fa4d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1064ac399072542222489ca1515fcdf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12329971392f2a311e33ae00fbfc977;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e63e179859faacb5aa4c6ed8ee5c36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f46628e1bbb16c855d8a593ca8f3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bad5482bbe04aa3ad1e4d910b88f90;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c4f3b81a53901425c0fcdab5246ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18110f73c8995e072c743a8a58d07a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8f0131ae9b02f249143e82cd33306;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e169a97eb27d0560fa44dd76bc8ae8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bcc5639de043260ed9f12f24b4e62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed3354b0243d33eec8fc3896722539;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b34e912da0dd67d6e18ba1b594c8f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7198a91e113079496cba5490a7a1b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34358a067d585bbaa248101bd4f91a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d8fd3c69b9fd28d873244edf43876;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ae8e7a78f8c6cc13b43fa28cc88ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0b14d2dc71b750474c072249c1eea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cafb17bce3f0d3c8a21fbbc2320629;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf01e21474679c7e60e50d74843f8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c011c6e4c51e02aa0c40f46c79bd9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35f19e9488e5b001c8382d2bb8f699;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he555d859aba5ee4de9cccdac3bc9a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h287d4e2c670eddbc88beef00268be9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d61166d6d218d4d1336a9f0d4232b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d77911fda1d1544366e9864890719;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea28586779f16cf9035cba998aa996;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bdee63d93de5bc04f4d210976d42b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90734747de54f7cfcaa990e25284ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h483fb3526714ab2730b7cd13fad5f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f457618da78464e39699f47f583b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14aae59d3f10fa2cb2713c7f620a40e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1409df819b20527923db27b31bb3a51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he350cbb3a7bf3f696f79ff759e1e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee27d1bf827ca478d89aa88b5f4cb3;
        #1
        $finish();
    end
endmodule
