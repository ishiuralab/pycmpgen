module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [17:0] src19;
    reg [16:0] src20;
    reg [15:0] src21;
    reg [14:0] src22;
    reg [13:0] src23;
    reg [12:0] src24;
    reg [11:0] src25;
    reg [10:0] src26;
    reg [9:0] src27;
    reg [8:0] src28;
    reg [7:0] src29;
    reg [6:0] src30;
    reg [5:0] src31;
    reg [4:0] src32;
    reg [3:0] src33;
    reg [2:0] src34;
    reg [1:0] src35;
    reg [0:0] src36;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3])<<33) + ((src34[0] + src34[1] + src34[2])<<34) + ((src35[0] + src35[1])<<35) + ((src36[0])<<36);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17eca17ef23226eeaa2385125366774c33875643a3728a49a2d7b802bbc41d146f0a9b481ee182e21cc7974f5ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14aa0b4c355029cfcc06794a7088af4c6e8905c999722c6889b574a41617ddac0d6fdeab9241eb3f1c4c39e98ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9d763a98ae3449d19d0494687ee044aabc70eec5cc961e93cd2c5db7e4f286cee4ec1cc9ff2ab112519bd8519;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99e8d3d3694f5a2afd107c6bc52121cd36ff9f589e1ce577b5d8ee306e1b62c40b7b1644ae02fc7f76f4b7d877;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138e7718e976fe62a85557da9628b72d2970e7cdf1c295cd601a147a29aafb28a17a6247a099461d8dfb68e7111;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h484938671d7d4392504b53ea8dace693898156be8d349184bc03faabc7cb0cc57ee7ac2c152d3215c6c2be49e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c135bb5fac3dde14a1fdca8fe342dad738684e21b23c9c710e24122235d994bc6f45ac9aa84bb213e83fa5b04e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153129ac7178ed851ead2c2b7d0cc276820294afa6839fa53033961f1b2f401b335970a0b83b045b34230717ca8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c08e87a7ca280c5ada490395bad175cb8c455307c0b2f94d464a5378f77b8e7ebd2f56dfa8d956642ad6f56ddc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h870d47cb02ad2d66603ed234c9f735af987ef6b49ca5ef85b3f15da6f316a7f190eb10d82c13529476eb371c61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce75943fd23f3c4103e3e046822e53fc80fa74fa7c309e987aaa348c18bbe5436968253a0164e7350f01809873;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd9a2ef0547607e61b8dfb40c26765da0bbe94f6ed857bcf38604c4c50f126e8e374d899c95a477f40ffcec0f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c85955d851b0b89514cefa1d3c42543a93b65bffb0d1885dded1143246201b6c78abe1fe2ebf1fb5c56f17b5c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h428e31f931af9a93e66bb452b0eb39f7d1476cec644cc2292f7c6a7a45fc5cf5212d19b6cf522f230364656821;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20d0672590c9db5770a9dd3f113ad73993e26ff5d082570345e3e8218036063774a235ded3ce006d3d5c6524ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed6d038b79934892669a36756c7bd9f39e26e24875bfe99cfb9592978497007b5dfef0172a67e17976c2d44c5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e6ccaad8b16a20fbaff5d971fb9cd50ab536c5ec0b3290e67f71845f983b704428e1954f0ed31511ee0ef3118;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0e83030c538a724b54a6ee193214764ee905a3ab649073da25636075a03552892ed00dcfd7c7b87889ff71da7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93e193ae6ba65730cc58ee6a5e3914fe0e7437c68f3bd41f841e6733299682b3d84482b34d3887e1595af4e448;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1847f41e927b5241e14f371f1185fd58046c4ae46f4636f1fb7e975a7ebf027a2f386f2d315294fc3deddf5fbea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16eb3a362c73dd062a90068b4ed912767da631aaf555fc2efe039fb858fa9331b14d8531c632e5eeb7c57e69675;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1275952b7f559aaee84df4399536fc6020d3820280d64bd64965080815c2b9a32e25e664d4edc75f22748873fad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f6a587eea93ef86b769a40b373a8dd1d60b9e3bd788d20124522474aa2b5c5063a7ba75c3480b156bcd28c4e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d46d0af62101c6394904622a754283fc59bfb5047d02df5799de8aa842536e9fe5fb1ad8badd60442fbbe7fd2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2d1ecb4929e9d4bb707182930b7dbec7d369f036ae9a38e357ea289b76b29c4d2a5afae1fb785098950187c1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdc70bfaad40614e769b4fad534da976460ca2d0a8a3862cf49d5c91f2a7dc0d4aaaa7a20e8d49d11a0c3ff43d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1495eb6874783e34afa6bf4f3e6ba80cb5686cebfb14c1944d7e74b3714636da21540625bdea3759d4124da47;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb7a32f48a8a4e9d96798dc9356ca82fe94157d74ed1a54ee9ce762e329ba6fbf2688f828b0155598f657a5c8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h399c9798c1b80f7600174d3c81e5d2d3692d734ff033d29dbdbe4fa8c5cc008c63dc3dc4f2365eb97e168f7286;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h913baf2cd841723de987e9264dd453e54d04d39e1a85240c9d99af31a2aa1b93ab44b9f49df69d590903c47548;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h745d6ef3327a5e7269b6dd818218967af4b1c8b5c59a229c43f1b841c3046e03c27e2a7fc15c8cd7a049d493b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1566acbc1b4307dfbf01b448dda2a2d703cf36060ab9cb38b948072e0495b2a5a2e15ae704944b80f75406bcdb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c5c43af1ab2eae0343bac0d5576d1a90c4d7e5e172ce16e97233e1967d87cca7ba28ebf0579fa5bbe5c6ad21b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc3f75d5195c2557588b33875f32aae607240a18ac75354727f1fe47e5fda8ee035da39864f15d0884bad35982;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8de93e13bb3a0b31e545b31dfa248baf49fd2369e714e7492b17bc86f05d676800d2b91d59b978122e4f9cfbb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8e1d5c9baa2e4679928fec66193145362a3205eb7afc8cd1b5499fcdf78484fb0d60b3c68ab99759cb2840769;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5bd3abf91a1778a10c4a140dda3e00df391236544434ec913f848554753ffcf0bfc7dd82d63ab3289036ab476;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1e6e6fa2e84c194f016a4c28aa6177edbc55fc11252452efc64c0f3966032b4482518ba6765111b15d2d42655;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5da3c34f5f6adf5216a6d07795717f8f36060e3474af498f5e9eda91cc61def008962d07689f9775a898f863fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea32231ed08b4523a4188784e89d788583584d4e4082c63ef34b91c310300783344a94ab50aa0d0dc7c66cd9ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he18a632a2563a4eefb791c50338154e490770f729ad2a4fa80417a1199286ea4819521a02e26522f9edbb5e15c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7b7b980004fab2c1475d9168912d105790e6ed4982499d524e7b3f1d0501553f1dd285b14c1d63b69e93da9b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1781e19ae6156c4c0cdbbef345f927ef91a4140c235e59f043f7dee1c70917eedcb714ee1cdf0b2b8e576154cc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a1589ab8eb7bd47c8489061c16dad482c41e3b4f05a1dd225dc898887c0f2e852bd36eb0511c622e7df320270;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb4055c0f402b3bbd0548c96800584de2544790e1b94b155237124f48efd976d32dd2e38913b68a3de045d11cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c2e3a1852e11aa24ae1b8872890416ad5ca8fb553a95df5e14a4b5ea45dbac8cb1f20295b443f5830948bae2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c6312d980ca84baa225a03033d3c804e3b2f3c7daca7a3463ea32b09bbce92a82d903e24ca7535caf865a1569;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1730cc30e6db4a979772ec7fab7dcf42bb7c34ef1eac2ac6b7318e0ad4b32a0ccc042130b0672539a2af8a3c9e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ecb0977742744e979dcd90d7e88442db4ea32045f17f2e46b68671367064250bf181fbb75c8b95f40ace8bad0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20b77f1b80a9ddd26e15b7cd4beec7af3ffb33986f6db82eee331015b0cf4c57712d643cbf958bf08dadc6aa7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a41333f72b30a50cb591938c43af29edc41d27d896b452e383cddc2d0cd4c70c7f34702b0f492e525a896a0ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f6506a48ce7ebbed02746ecc25180f955c967d845bb1f8f8ae3da60b3dee6e54aefe3d585caf33aebdbfa4f4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba6cf4c7396694f00ec4d3be573927ec207528c17559511475ed27643e468e900da6ac231d5e763e58f7355a4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12975de092f81529d58611f21b95ecba8da9de1b69445cad5a3fd564e3630ac6daf00957657cbd75bd9d42ed73d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e81b916391048bb265b22a1f01155b679bc4da519e69649575c646ce58f5c076214b85d94ae7964b3de3b0c67c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42ea568e2284cc00893d7e4de8ca6ab9d9fc80a62eae08d1edbc0b85e6c20c01cba2a129e3d9ac43b6a3ccb3ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1311f57162fe67676631c8f89b453c8c87859cc5018cefce6a46ec40ef84ab9d10e49673a291d998300c95dc7f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f978e6758ea98956764598cc5f91362b10c4f1db7432b18bdb80639bae77dd0f38aadc850819caef61b5cddf71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h162b37b8c27843e53ccb72d283ddbd56fdf336069a0aeae4793067713840cc1f6c333f95d9fd2bfba3d87486625;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d45f3e4502a59ae681ec79771c13087e908bb82c63827c194e70e832037299161535833fa7c3ceb8cc565cdd6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb550f4049f02860fbd60d40439dc7b7d33ddd5541561ec5f0ce8bc79fd45f284dd51f80d667f9abcfc0229414b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e65b3442625f85becc7f20618167472aa78b01ebc4814e0e8c130fb63947cde84ca7fff1c723a3c9b8beb46b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ffc62a280b218993e52f09ed748a4fded58e867f96b83598efc10cded5a3dd15f520bade9c2e743a9d8a391c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1132ba4c7839890d5c6bcb8fc17efc92cd121992ad8a132c81d8db763e4d42b8665be6df9851a1a9405e11cb3e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b3e67f44572ed355ce898376c2b23e04d38f1f17df96998ced4d61659f6b4abdeefbf68985708df90a6c961ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dde86de70f4b1c096f2b8113638f29a018dd65dc869671f95ffd53dec2911182a89212348b5dfe956d4aafd9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7df06c8bcbf464996aa8ee2e5d235fc0c3d074e54cc7c773491aff2e83eae9bd934e9e23c5e2c612a9d2fb6fe0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1667d703e325e5025ee5c26e956c0373477aaab3bc38422fadba3a490241fac7082eef0c349246b4fa73a2a68fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159099c4a2b4775a2b7eaee8b496eeb007e664e4eefb86ddb21545c770e14eab54b194f5883d1b1f64a5d5e43e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e89b135abb5fe3d87a313c811caaeae2fa4c105a76e95065abc058e4a1fc7865cd804d5aaa71e7c780d3ac974;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd76323f2a4e8c350b1757e57af8de18819b2ababc04ddceaabf549c7f52bdff6e4fee45a713cf40da26c7e7c42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153fd966b9b7f6e746e890922d4fc1c629a3c0741c30ea88e6ca28f7641c18a2e8bd840ef3eb25e07cf52bb35f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a100acd5819fba058cda970a7414b8d447ece90a53a7cec2025272a4fe675fe1f7d99156f7276335d7c98dbcc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16dd2662b472fa66ff0ba3fc2daa5078d025133bc8c6c2d86924dd0c3b16804217223dfc6d46e58c60f4895ba8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h758a6a30f8cd9f5424e1d62d6ad1853a10b6e8c81c2f5590d11201cf2bd1af705cfb3795cba575f92e0561d311;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e68abc321b1c406101b07f6480ff77ffe36521443ba901a60c4871fb9a45afc398b259e05a07c5055e30dfb791;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf62378cc437394dac227a41e1b03bed3e453ebd54d8f148341c7a8e93abe1ae64d12cfd8c1505f668c32e9a81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa58717f1e4a3ea15febdb5171e7a0754a2a3d044871194d8e35c421354893d1f664da4afe51a2d75c02a80e7d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf760027665c02de8d996e368970be26ca617f3d1d5ba8fbc2db977c5b5d2abceedc7e04acf4fb70b546d5674ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11dc9a02f63b6f502694b64b810892dcc3713fd8d393495f396c80247a94417f57eb5ee70408c205ed4c78a6630;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1526e5612c009a0f6e54434b2d0e9f30a7e16271e8d950559c4b361d611e583b8abb675d1579ea63aa4589176ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11898db757ef9019dfc764253b7eff33c71246fed498c17ea22c54dae77a83a7eb19aaa1967ac6ff6c22e8822b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e54b235029ece6d88345b58ea3c70cc6d40997056d406f27796f870853b177f7f26404c4356839719da5b3a760;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9cb6348954d348f3eefff6b8065ba1977c503aa50a13d9e05b95ebaeb73ce9213b132e20f248a1b7ab1ce3f699;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47e2083d2ed113ed18c698978dd3ff6658e6e9eb59983b52cd159257c0c77f0ae1728e0141d5a4eb631d3246c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1060f994ba9f32ccdb75c7a5a4238c7eb7d250668b753ae48b2d96c9c4c79d2d367b2c0b7e231b98ec47ef98ce8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h788d20755f7d19887cc20217b3ee76c56845183b58a7764af5c3863761623cc53b61ef16f0f32cb9b93bd55c95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h599f0e0885a3cb89c810650cd3e6233effee683eb2d12594728275ec3c8abffa063ee69fc045711858a3beea07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15750f719a52e673f58b19d38b905bb1507b0f2ed34efb76a0fcbd18aae4dfe620dc70f0d21dae25fd23ecbe3c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e411b82a482e84e49086c7a435fdeadf59fb2ef817c3b2d0f767196dbd7361946aff22af9afda657d0f5b51103;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82610691535b2d2332de887a0c082718d6dc900520aac5cd87bdc74a73307fa2d69348a665178af342d416e83f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2256ccc18ce25207b1c2fb347526af9ae078080962e95457c7cf1f74dd484cf5af5802feaab6e96513531bd14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8edde4944adf609d7c0f4d050e8c8316140159fb28a78bac4f3a082ecbb645bf58cd46161419f84aa93c68c2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53bb4c3840d148e3d4d0d98c859352cc2881351e6606104edf12ed9848afb1c0e9838b239562d7854b2c42cd28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a657df238a97b567b2002d80b3d818f77ef1e037973169ef7b8a9521d8de8bc8ce7b994ff8ffa4534227d1a4ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f6d99e7acfcd3829a63327bed591029d4f703bfd2b85a7dfe8fac8c543492027fe41364a0d2586f446ef65347;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18dec47bc5f8fd50185c1296a72c2b4ea8990abd149f1ece19bd8f0ea825921370c4dbac9c8a78815b1b00f5465;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3294ae6ec1efa8ebd4e0c6fc67cc288486afae0538c20875f57bcca58c8e5cd020e9e0b2126e1edfa7acfc07a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a337b7a12fa195e0a0884b7ad59beae7e37c01891f2840db10090588237a359f5383d90d8a815dc25414072297;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117a4f48237f2f4dfda2dd3b36704550ce1c7ac9654a0dfc86fe54eca4c647d7fd73f1a8f83b42b5e564d9eaf16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b71f0b6fa55433b1b9ca3d4d095684006fd41ed97223bcb018ceb446ef1695a6c3212695335156fea908bbb32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a979625541bf60a1fdf44e910f88445669a6258bcbb504f150d571b26c60d6156977e459fc35bf096ea6e26928;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a870249999c76d3d027cf7b5db6ef2d91258c111763ad55ede1a6e571cac48c4a79f99dd0499ab79e1ed443e5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he81ddcf374a4357a041fd242d179de711d8ceb5ab7c38f3d237a79760fd24bcfb02abe810b7c35cfaba52ee40a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9653722e52144886515921eb25b558c7071289d28143382945633790f3d0319780df15483dd205ab84d1266425;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107466eabac2f3e9b2d0da70ee0cee31c716b3138c9c7b9a3c853957812368d7c38828c7f8130745e41eabae7f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1feacb1c1c1962524d38dac9020cf0bf165055863968331ffe2ff5963cb783c10d79eb28ac1d9145322877a867c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a1202a2facb4908cb8c60c186e37d2f150d6ee660eeb20da7e2a04e01a9a95d80e2280e771d2a32dfea77b24e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169c68b904727b25fa29278b445b75525bb06380c298e8492d4bbd89e14f1147b204376dc2072a79f23bdedc5d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1accc1c478f133645a9f7163e0c86a3df92758ce4974e269ad92a14d0c14b635d212343e43bcca1a3bc2a2e1ca7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5002ff8206c7f247e5ce01ccd5e0197d6d725267a30b046d9906afdf9c6b5f37b10f1b50ad61c4979c60e6fb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1516a4b59b34753d632f5f09303e392f418f1ce3c1e6ac50d05f3be1726edbfe642bcaa1a7ba92201ef96679b71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefb48de9218aa3424a596904e1cf3fab2356266b392b052b72f9a5827e9303f866a61b7d6573c91d12c2c2e3c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha95b397962069156e9d8b19bc0c0090ed337c1853a7b929129b679381aa56e8e55a2ece2ea2e7b08911fdd7b96;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc75ff0ad67cb247c83e8092d035a0d1fa79cefbd44d344b0b0fa7fef70823922bdea31e8a9e8ec9c70d05986c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27bd995e07d87ec34cf606f34622c7c0c2f46d40159d51dac68fb32671a62fad6f93f991f02e608680bff00ac5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4e81dbe462a9c65d076844bff8680637e2988684dcb7808d9c131c9389e316c336930acf337f2cb0c4fa6c7ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9903c60678e315f9fb983e8bd2b60f108aa0263c91292844b911d07fffce9887e52621b17202aceeef9a2053c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72f8b485b219cec7e523989090e5c8f6bc7b34ccc164ee0cef50ca4727f9e369b8f9f0855d23259707521497c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36a6f61bac043a3a33c2462653a9ba3546e444e75d2e265a6b3ff1518ca760391f9234f63b1ac623985788593a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53c449e7105d796ba23479a2853e039571426e650ea6e471def5d8246cd34bdd8f58be6d7436d9bd97f7486b2e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5853847450f36eee2dfc3e3fcd1f833d3c9193e6e2a7178c063eb21f2cf9d4cd86ac0a170469d21b9046966aed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h959f1e83bbf6a90b6404525c6ba96ead378fbfd871ee40edaa97353eccd664232cf62a8c31c75b4732fec9cf6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d68ac03d86f64331b2ae0058416acdc124bf79d77b3e3f30a03f14c8836d98ea46dff7dd383f2ae7e3ee1265e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17da1d42c09d00d04270a7d1b5a59e0aa0809b01d287aacfe3243ace8964ee1350641b152466a112bd539669124;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3e028a736c49a675317226cf9cdbc65567bacdf3122b820e1239a54128eaa7411fc70179ccc0f83d8996570f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1fb0444b8d13459f17988cd50cffae8b5d277f411c8b4152a19d977f84b6a3b565215d2345bd32958e1b27948;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c85a293487d18c97563737feb2d8c72fa6c3779b57348c546e9cbf03160679e888eb87f144d16966fc40424a36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3665658838204b6d4584a9a8c6785f698c5e3fc32e57104c7cda62dc3f79055b674f1131376b3d5cc4d902d36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h814d46e586d9cae68110cac40cdcdf3834cbf381cb0296555d0554f16fd7c18d3935043cb46514c9a0b529bf8c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3dcba54c19c9e6a783290a3e07f2438c44c2549e83e7df7f8c44238cebb8557f83ed53914bc3d4c084fbe8b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f17603efa4672a7b681ef66cf3e55859d3753da79af900b2427e00d166359034dbd8780cb4835ca3bcd0609c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13040430d50b1207194f7c09a8e4c7c759c79b527c10fd4e5641c37176a01c1a414b6f8e1ed385bd100095dfc9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ef69703ce18174e12d898a864482cd3b01b1d9bf4545b4b9bb3370b08b2a417c5120aa6cd1b92f25223495c8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14873b3366b299f002539a9af36eba319916afbea947f73399ac2479938f8694e906182f9b32f780728db98fabe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c6c94bf8654e51a6ed4834b77f0936d3598e9b4f960d6df28c1f32c82c2c02a02a8321d113d2d08e9f8021f39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f6a47819de674861ef86b65eea06f8b56d298f78fefa0d8384e9120ff34e3839dcd12838fc695ccc41bc81561;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a58df850f4a98ffa6638ec264341cafdcfbff01bc19b6ac1dc3a6ac456d1196169b7634776cfc3e2f99bb4ccb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11daa04c26a66ad5c0c4277ba8914d55f791363a3e7a3a49923260ed2d48c43596ae2f3060b8262e4428994604a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105cd457f5dcddc2f282cd7994bf332e4d3b53b5b03b3646f311a2f3cf9387c72fb5de9a821daf3b20f40571939;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce9e5b7189c078244824e48472c78da10920dbf2436e4ebbfcea78b37f35f1068ddb8349faecf1b878f4c81527;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae607cc068d3f375fc6c90585958140498d000868517800f4b062b1bd9e4f3ee383efb516aa3ade3f6f542ef38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf12f049d02f73e248dbb162ca93f87af0cfe9e3fba680f4aae962b928d9a0775b763541eef79dfeaa7dcef9cf5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h210572058c0fde73b8c2ad3922daf55688a9d0208f99ec0efe624215050db7d5a76d3d555dac82ce4ad0950b05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9866ee1566d48909b65917940fc69abaac1869c434112b153838d63c6ffec2c5b0e0c6cad2158a71acf0c84de1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfb676dff442bc6151a10b165a1edc064c2f854d4420deb5727b3ebca6825fb389aadba1fec9a3f7f9c027bb06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h415cfbfcf2bc218028eae283437cfe2010ef6a316f4d603991bffd07ae70d87d93d8304b2eba2ff6eb72ac4049;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h463643e9b4f4c06adcf4fc9ae6671106407ff2052cccac9d2245aea39f02644a32ebc3b2b390fbf8d9814a59ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b64d3a5e34cde852e7efb59b8ff26f1022bd119725b99dfd1855f69339c2c12b57e5a0d871877511790ae1e7ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10752d5b3ddd204268130f4dc2f45858fbea3ca78570544383fa2ca561576da469b4efe7a640973f51d8c26d1b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he087f7254080d2f0889247ef5bcce4385436cadb3380638a0f39dfed3b1acfbc588ee2934c384565470c314dbc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c8344295774fe5c677328db2a2f9ad523b49bf1c19dcbb1315ec71ebbbfb1c2747d3919935c552b8ea88c374d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17fa38416879a57577277823c024bc7679be8ccf00a738e1a21025ed6cb8e7e293225cb41369580cb92aca39c58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d93d55f9f8a016bce5b8db88de57db63be8637b4799ccfd704a4020c9b3730681b5117d756611f3cc897be28e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7685b35563801666408830d69babb60f7f9592d48ebdabe824c666aa8bf837911ffbeae3096bfbcc4431fb689b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcba6ce82abb97676e0812d20a500c92cdbcf61cceb089dedc31a63299c97f31e26fbd44d50774cf2f3230b82f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a1e1218d65cf1246fde4fa8d0fc492e93890cf51d7aea5f58c8cf53f08165d84f96a5e2cdc109791ca5edcb4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bbe2d0b9d7e614ff345fd30ab7f7735de4436d36f8c7dc7c6f80079eadb3595a3180bc21248e58e7253dfe9c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147ed5a4760f7a3d767972cc59db40c0789f02d3cafd4e92f0243036db979cc5a95400f9a1bd1cb60c57eeead8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159627eedc333ef099f829c051e48da12d854b2887d09a75762a11611b27be6a05f91893bf4f4c3a206317bd065;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1552b043455cf1f3aff534baae792d750a594963017782cbcd8bd1ebdea498ee75d45abcf27028b8400f6a40d1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ca8c54d938d9dfd05e4a2d2a794db660ec4da847febf371f6c3c0a3611ee9f9ad0eb56ce82ecf502f4d0d4ac9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2767d3edb0cab38f3285e282aa9d24a0b8df95c9801a268040e5aba9956bf4e875f75dcbe5ad7e2c7d79f2bf82;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h96adc09700756d31e3b64a9b76991d6c3962f858cbaebfbe5bcbe4f8d6bf0c31d70ddad14f55bc7f417f7a9e5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181ed59771d1f3e0e3809a838587b219f6f58d24859c9268f65ae6df657ddfc291370bcb2db143411c41b96511;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf160036fc1e0cf47b043a9d3b5dd08f504a48a283f5eac64f1c998433aec0fd2fd5bd834ab325e0a28f67c4aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c4e918a9af28c74dd7f799cb7198d35415705b6b317a32328575f8edee9981826fea1e5ad403d617137ba86f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1bb88883b5651cd1119e761b44c309a399a70357a073377fa43794894e29bec7ad145392061e6d409106d4067;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1deab028aba27fb3ad159b5abc2a708dce86f18856ef98d03ed4a0dbee45de35851ed720af64ecdf586fe9863;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76bacd19706d38d4e070c4c097b1d0c22dee8a737718c78ed440e3e8a8047014ab07938bcae5b5ccb942b5403c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8da38067267b094690842c48c79a3fec29043b14ac327f1b2778862d5e49cdf0c8ac8e9551442cc19a70c659a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d83f7e67e5742dc6bd8f8b0ab7fe660e2134728aaff7570a85ac72ee860d54ff8f3fdbf652882175c8ace08409;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f5afe492d76079d79715944279d451469074fc69d6b24234716a6c0cfaf5630f207fbe6993fadc0ef6a2b233f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h534332f904681f5ea34199112165dd83abb509abea48f2766936b05c1bd7447746389a39396bc0933ee4deb4f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1884f301b3050c7b9cb5d28a8c977e352b6a2d45567dd77390e8055c9583bb5515b4e5fadbec01a11b445ecbf6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0952f2bd002f06830129a41ac2eb68986060282882b1c1fcfc359a6e45cbb9489742ba3e4d4b2b794d785528c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64bf548bea4395f00a540ab6053dbc6455d0ac389ea5ca895ac357898f5a02152b7b440a4612defdee846adb6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecbf3d51011bbf83767b1e69c6ea2b8d57f4daa95845eda19e027b5040e4711d2907a38dd4c831e7c56c470a4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef55a24c535f7a7426cde4b50bb16a8104e0e76b32564fd4d5a37d239dfcf64016efa6bb56a4a31ffb3c32c54d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9e10d14295907458c793db6add856eb1e9747a3ed1eb2bf1d3692a1d63c0d490d05bfa5fb9c6f483a04a3f87b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10782f834190b38a83dfcc5470dd61e47b5d0aa603e1fc7c73ca06ce7abc8b22c3f387499811a9de9c45989f69e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94ea4b405ae8af5fb5db5774f25ead93f3bfacdc52a5dbf35d473f86a54ae4f92a2257ddd941c7c2b3747bfe7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfd22eb5946698a83733153c5b969b443960900a8354144b547ad7dac9e32dea95726ec1b5fbae6f65e0eb69d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144bafc784d10c0794438ed1a62f7720063e3e64286782f3ceef67a5b4148b6f7f143dc49e87e24d3060a912f45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104df6952f5ad1a803882ed599665b4750af589aed1d6cab0dec07a7432e811c60d3f06fad96fe8914bddb44832;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50d366cc79cd77b3a65cd492d03bd821d48e25bc6b7cf9a2196a8957dbee5998cc94765f318048244ef2f69a63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32a4f6bf519171fdc4e324e6c57f4dbd2231d5fc7b768b063a5f23e001c881ef267d5ac3f8280e076a20b46428;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a772e5a20144bb962de57c3b92fb82c619f535e930938590e5ef928c474e6076cbc5b32de39ae3e40ec70f3a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10eee5d5fda75d64914e2c9bb9c30d6a2334501b8cf43cddba255b4ba433bfe358d276a2150c935b1cbfe4b6b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123e13a0eae68b40b43c76d5c1184e36d8ed10dd9c9eff8b88f6983f1e8fa9c82a73637d8332bb8f0fd99b46bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d0d13644ac5aa7dd3edda18f9f56354169acf59becdab423b936c940380bc6794dc022d4857d5577d4f0ce23a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6694c91e032ea8f890d3ac9a58a09ea26f4b7e42c20979b8c5aa58cfab2dae253f739bc7e8e15740412d498108;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd40a14dd36eca09b30481e9a29d18aacd2bc0c84368ae5a65cf29d85f5d8a6eaf93ff3bb58dfaa53a058ff01a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123a8e5d39948bc0b4cdaccbd9f32c99514aa2c26e3b105e81ef3088ab1d861c1cb96f8a90a45a54d9457f7c32f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1091c208f385680ec768cec89f8d66b004ef407354a80b58c8b2431357893e19444531528653fc7d96cc1df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff6e49951e000cebc0dc1915de288ab2ab50cbc81ff09085704a48e632bdb08ca584576fd47205eab3d6ad9ba0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8e5c8b152b76c0c4afc8f44e805471b26de7f1eea0e99ec5d7f075f3e9094118ad0b373e3e476eb1e69184e02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2e61e5afa631f1f91ecc84d1a052ef32c81a43f07d5500f370cdbbab2fac33b6ed0ac70e7174da5bd9cb923a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ee90fd1b337b271ef7890d53b01175e61304f721fd3841a5e288de959a2b07eb4f5ef4fffe2eb7aa26ea0b5c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b0db07a8986b0d8a1fece2b45d943a96ad59ac97e2362d918237443365291a72a4b84d1f59b55d17e57b1fa45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dd56ebf7f597a49cd5bfbda1c0f88c187e4ec24a91eada2f6fd1354f4f2998a33edc7e36e86fb7b6d437a5cff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b2d52f3dbf5c79840b7a8f7e55891fda66aaf9036d8b7015e0790c638daf2e8b23041935e1087555cb62d2654;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b20fa88bc954187ec74429ce9c36b170c22fa045990b32f383123e67aaec72d20b07bb6dcdf4dd7409f690373;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdd337c1d6a4e9aa8c2f38cd0cb4d312b197117992622fb30da654313f5bfa2c79bde4df0c0c12ac8772e3443d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fe0b0daebe79fc56139e257c299bf285be4facffc05d6d24dc2dbe9d4516ab6ecc4dff711281a5c7a48850ac6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4532722650b25670fbdad87e0c071b1775f4ba62e4032d657d9a5e2d71accf9d734c8856a72f1495b2d151323;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6cbf99c040558f1c49393c3e4ca40d9b44c65ed638d2126a5c9f3fbccbf35c54ffaad16b4c212a7d1db656bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89808cdb365b4c00085285cf9dd3bb78f39dd530f2fd68a351b1b2c94109d6e7a18d4af94a9bb0b948a2e157e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a993feb671992a9357762d821a3af1bd9f9e24482382155602cc5b8459ec21aa07c3d6b4750431a7b9aa12d43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1873a19ca0c5d617810f493c42118280267bda4a817ca68e90900ecfd383c4e75b089528160d8f6f48ba438231b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb91053c346c361da2af94fa5f2177fefd4663fbb77c720955f3a6541dd224886aa54c37750e948dcd1d7124315;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he22501fc3a121ffea24fa86696d11453555c341e12e7dab9d5dd39543f764455e4746e1e9b3e548f304710103f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f267d1d95d9a3614f6980d6d25608bcf72d359ef02ee9eb732d20f9581a3fc0792bec5bd8bdf103512932069c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c80361c5c88b6febf8497603e58a371c1106d2495c0d6a27c57d4233f328dd1340e1e04ac7248ea078d6da51d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a408288358fa50fde20e51e8ec557437bb880c4caba64dad09c0aa2ed2dff0add7ed002f88c95e62c5db5b69d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a0318325247cfc90becfaa43492c7a298d9c5fa56d6e6561f52fdbab05a5b4d00f40464c097a630d5ec84e3f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd3d12c57d47c84903e068694e2517343cebe21387c57b319dcaa4186716fe49ce2d5818908059378f4e818ba0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c8f6769c5d952a6f8ba383bbaafbf6c5b3076cc1faaa944303a3c62ba1969bfc503c0df7e2d96ef3c382dcf71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fac2dbc737d89ff85ea02e0947e965803464bf546c0cd24a5b7f7da77cb964ab11e3b40f4c14d1aa1a297c52a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ec1bb5d54d24db579967e71b365e0bf252a5d66f6977e05eb7e8232f270f355d2bf226f8c66da055cb2931ce9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9b100150ccd922c2a8ff73339bc97fba25d46a8f135b79aab286325c8a4ad7435fb5579c85a2124987d1f020;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da1ef1e84949cf3075e4fde2a9bb168ccffec12437f285c320ab10e7e9ec794ecaf5c88bdb8365119a841d5977;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a67c0a876b3e4820900cdfbd7a8f6b8b7555a512f9b687ec57a78318c5998ac56026ad89fe6497ee8d99ba582;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df779448517b09ba33a4d863d71b12fd8d4c4f397be7d9030e05d8f95fc7e0beddf6b9965639137bed769c57d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128a9d279db43871da8c47a9dfdc2537ba57cf31d007d865b500ae973e10c69fdf305287046fe55e50fb3e05438;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc065d2ecd10b1bba51cc3044f742c14dcfcf3598101c955a8afc7229b32f10e4c0435f6727c3a3dc70a8d783d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15072ece9c738853182fc86864ecf6d6fefe3fc3b9e385713299a23483f13d4d7905f2d853020f0704153c0488b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f197e0eb3aff68074a61ff5b6249beddf2e851784ef9dbae1c1362c31a1cccbc61d2d27b7d6333d9fd72a38565;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13181d2d140e751d1075bcb39052d16329adba3f911eada8ad8b569e5cdc22dab70d218098c1b829369fc46761a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0fd11b0b40a0608a48821b5c8297d5fbf3aa81082e065f1865214b615ea820564dbae59b7bd603f30194c3cc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51b5b9c85bdb788c179ca3e585f0e4e3617e2f61367f6e484def059bb91293926c25f8455120d3d77f07760fd3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5421a5dee167b3b11c9215206df9f631c9f35c780538152acf3b2a8c93ece04a2a6a67f442b56c932d24c12ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92f374648a129e35ccb441960ad96c5a330cb7d0ee25228702b4a96b1eb5045fc0021914de5589909178b1a62a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcff7c71c689676d031ab5ec68ae448aba2134e16926ccf401c5620d91e1cc11440c2e837c9b7618372dba1301d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125edd5c337fac2309b8d5e993f2d820b6b8d56e571b173102b752f78d9f6a21df22bfc7c901ae8c2f6d5e030b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197fe37b3fe86373210afebb554fb0c4ed575c499857a5abc264c13d1bc2c42402e9b7eea8e05c1d76be600ce44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1269145dac06c4a8b21661c5d8acd6e7432900c3423311e341f414994ada3ffd304a848a9f99f702557cea88e48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61fbad38bba5045e428939cb94976617f7b536fc7ffe91cf3664a6d54821f1ac1ef7266cd841f3fe9c11d70081;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he61716ef13cc8dde95a5d8dc311c64cba1f637e2f774e801116806bcb187cc81dba0bafca1db3ecd38983b78a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdf0ca7bd50ec6012b313b463968d706a0f36aa6206c12665c1068f99b131f6722642d10852f4e44af52698353;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6025ec74fa645deda64ee860a7b1369eafc582e44a2bcdbc65edc119816f01c500288f63bc56389e630dae9a45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d5cdad82472dc103ef8c188c529b0ec34b2f65f454be9bcebd76a83837075b4ce2cbf6545e1562c6c7df0fcba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182cfb4b5a919909530a930de2f85e68b1ed7dc0ca400b7f7e11307e32400483e27852ff1ac8076616e4fe120b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12aac76a7b2ece6624acad94de1df1bf991d4dfff1cfe1d7d9c8a0e857e249630c95d5ff3d5c5dc966849940f62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b924b07a56ad448ed09b4aed96d5993d7f8ec16c5b012f77819089fab676bcbdd0a6f35d9d7fad35b44d89ff1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h769f4057a3e8d14d901f9978da70107654e9d4bbb15e7ce8fa3f5da3c655ce1c7fa10e657083af5f6c285f54c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a53525c8d85adcd001100e3192a401944844909ea047ad86ea609f33809cc549db7b7bd2b3cd39676eda3f3ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd063a8ab85dd3994c47657c01b85667cfd6d79351a898e412f262a50491c2f855cbca240315e67bb7586a1c09a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb74376c98834eeead227fe6a3388222fe5a2322f8ad4361a3f7128f2dfd379d205b5e4d7932d11d9c491b6f834;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ee90fc82510d255b62feb5c58fcb4b2c1ce17cb01ec79c1b58ad61a0ded0a43c36df2188e2cbc4f4336ec7e8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he79d01565beb104c5136b9d6900a5e11b7afd4b48cad318d229a27589429e2dc28201733b3ffd4dbdcb12b4754;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d9d1c4db8fb751d7ca71e3476bf320f1026ee53a27f54ad7b9d3c6a76b9147bf97b9ac93db5117fc1ad49f69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18dd71b1595c5fa336ff8fc395d0e3a5f0db54e8c8277735e5b99b6909ac6442d6d033ab9ddd9cfab1a2a49c270;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6add89950bb3e1c5ba99c106b786665ef4a00ed95c5ac0f27f4c20ea9a2204afb786fad7b4b919496a440c86d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf75cbd524d4baf761abf5ac1af645cb42b2f961da98c46c6c0727d7b1bdaeac3435ec89b18d819a6a190d8eaa3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60968fe7862e13afd62a073d8daf3a6b82df7cc4b1b46d60dfa082bdc2e8b7e1d94db68a23d1af5d29b6eb1e47;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1dcddb140e4b207f100af6f58d5de3d187fd14010c381fd5b95ada8c71347b990e1cb574b11af999b076307e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7e3cb89386146b1019073f8803fa21b4d478436926401e935f2e72f5f9b2bd4f6d34226664bc9bbad2129ec62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb048e2409bb7fe42e8bb82384457232cb1597e17601aa48765de8cbf65778dc0575c442b6666cfef9c779f10d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c80a50cc17f82e25814592945ec0916794c7e61425ec02c53d5f627d9260da45bee460e08f36a6e849e6b02d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bffad8d62dcc74ff9ade677367140f2fa9c3b3210f92cc21e0c28027d9ccefe98439bbb3f7bd42c1cfe29d3854;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1722764142dd7bd0c69941822462df4a28a11d195ffdde25e8b8c2d98c7fec330aeb1be8ec04e3d62299350fcd0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ef88e6eb9bfe858ec980b84be6d1847ba32a4d752f992c372a600cef9f957c3c742d76ebfbc430b4900dd9012;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c995fdff595e475ec64c274d61ceee8cc9c465d9e4a7af1e17a490cb01f15a7484296339e1716e22c12676edc8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d0d84c365fa7aa2f2d0f8f3a03e3535faa27a6f76b29a2cc58f17356ba9b8978cdb447b465748ab98800221fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136a69018e7b01ba7a8862cbd1d0d35a588ed01d17e146ab0e487a2d0495a49167e1722adb51cd88c138d22535b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194f202047a52e37a7322e154c6ff87862b6bc24ba90d854b1fba2c48a84469469273be82d9c8fa5a186d99e273;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38c003cbf8b76d697c7815692255cd6d2d1664cdfd3ba921c6677ded10de2213c75419e00e41e8e3a9376cb7e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a847c9a7ce84d50c5b59ee92691aa0e2df850c3f7405cf0a8b27097953c4981be6fd2a218327c61516d7520c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7f986bfd5e21241a2f09d25f884eb5fa5658adc3cedc3944e778b164a22d89e5ce4757783e0894a5b250b64be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h995539877e8d95f3fae0d1848ce2baa9b5b685f09a6b663dfda2c891a8cec83fbf460eb8b4a197a85e5c8a4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115836829b8ea3fadb1f71c6e7e3b7eb31bcf669da404b4bdd0f15eb0cdcb7875d1c690f2bd4ad95b8eeb0e7a54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a51b9c2ea4a4d377db67c74362876660ce7ef0f5da24c2fe833f5806600bac2ef8542085e6df692eb0ea609d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c23f486d44cd977cb3775838faae77bb65c363209576f6311685af1737e63f28f15967fe54f8f06d20a7ca042d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d1dfea755fd6511b7e8b5a3280f87662752cb2c8690426da73c46c4358e29dfc7f7c017ec1bec30e691702b02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7034dac0fd4992e28a5359a116ab3df4d56bcb60159ae78b98c1cf7a3d5bf92de532737a48d487db35f0d19b63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc2f5e4201d8b44aa008d7aa940fe8f7e9a5f025424ecae17bfa4a98c1ae66061dc12014c7c63118ef8c98525b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcd0d8204c6d7ab2750f5f282b1271c980b51ece40ded98348ef4be905199ba6171d651a63648f39cfbb7e56ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h799e872ac967f26e9134c1e6cb1a5545c989ed495a3ed0467118501eee89a64af427913b9a02d14c43d2696af3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28597f46b31dcc79353bf9aaddf0a52acdacbf7d8206d58163afd7fbf22532739866ce85e85547801793ffd510;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a431b9f69874005e4eeeadb9ead37b714008f3d3a7a79b6bf5c79b45dad4f94803cc84c164f32d32e0a8e65bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d62d6a175af03ea747af58273a21f7eac4167590c65708810fad6c5beb433a699eee607bde8569f844efa949b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c1664635d15b471e70d491e7842ea536bcc6cdf1f443552719b9de97fb7f38f3cdfa580a180aa3d7872be54e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7569bd9f84ead6e9c4aef55f101fbea835cccf205dc066da872229c67d36b65d176ab1ca440e69b24f5ebeb126;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf97621b90fa41ec0d654beca501609956a3a378cbf66ee6a8468da535e411479cacad09cf21c9db9470096722b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35a3e66a943ece7a63fd4dd6d2b4b3f190895c48e8f9aab02a8248faa896f781ddd9a31b8dc67b00beec579e3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198e8e6c920aa8e39957ffe75614cf9b86a960f4eb3c6dff01b0329192b1ab1764bb4bdda667304cc85113a34ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb8380004f5e45a0bcc0dd93dd7a467d49c6432d3ddda438ecf1c3b1edc18739e4ebe86cd721dc226df270a707;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196a28112efb15a3639b20911d22c6a408a1a4df0f4f2a7541b4277072dcd0a3cb15173c10d3c35de2621f5bf2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ba74927eb44d9207e143fcc1395ea027510a22dd129547c906f90a0b373b33f6fdf1b5d66d26431f3ed0b84ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33c44517462682fb30818793aad90fd8101ccd37d5b9b5b92da6b94031d8c52ecea42817122ae34a302cafe67c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14086dd60a401f1a942cd00f41553c2bba24d9c4dbaec58779140b3229da7dcacb0f82474930d38407af9fd9c7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78a363254c36157086ab286859fdb9c90668aa99bc76ac7bed1d4f9a2eb061bfc5bfee0974606109db55280d46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b6cc368ae31291cd8b97645f71420c0b17257d11d2cb12d07da6715d01e692346280190fc2e3b1724e361d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc77ad279dd253c6ffa6a70ed913492921119e72e5b3770c052eaa21f2c7234d95a870a130e359524bb53157504;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42229c85f4e76177e9c2588ff7eebf3afa5f627eae866f677d2d3fed9c2868236b3eacc63a3f9b91d172c4356e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a69951575b9ea7e43150941adeb306b68cde6c46797806b4c2027b5d82ed761f3826e01323e95d7a6a2f06b608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db95f0af124953c2c30093e2ab7f253b0a31484b690f31395099488101e85e5f0725273bd3c60d97117116a471;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec354075f3b65dbd43f5054e883e56fe809e35f1edb1e50c0efe7117ca3068a7baebe684c32d5f623becbc8488;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b31f0425602772defe683c893854981bf1756d6a4172b1a4dad617bef9f3b2b474ef6a493e497ab9f0d5d32ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'habc67cceb6b993be5788605d6a2129d5563f0ed6e0c3e3b33b062c6ced98eeea08f51382313535f650b637139f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16be0a71cfd1bd3ed6275ae8b45910dcec80b632119136cdbe5147ad8e128e6d87dfd234e684bb48c9df64d1ecc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ed986afbe2f05e88afccab3c8e499123b790adfbe1b502569bb125f27077b43b3f32b5b96bafb0ff5f1d7f9da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7cd6097a26d2b55edd7b992c3d8d7b4e341b8b2b5c0939c586856bb0c7ad0d1851886166183502b58e7f2dbf4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159793f94a66904c826167d553a10b4460d763a7475a6464ca1e88e17a065cc945af0773bf53fa962ad93613c54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2e4c60a4fd686cb75bf0ee0ee28cf070a272bacef08a47a568b382d8384868ba5afeda2f84a12fcb12298e762;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198f3f3fe06a3e633e143e6eecd4117081ba0d96bcee5aedc460306cfb6494a7cc2bf6042a2772980f4add0c38c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec2f558121e8bcc529aead48c35d634e454c47079194b0dd1af36b06da5177b5065de5174b82bb66e88276c9d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b61c71e32cd651f5c29323221ac791f1e92b95e01bae8574a47ad577dc633e8a31b28547792a6a859faa3082e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a10c684ed5f8bbeebb61ddad95231a137e73e4f86544bb5a46a4487dd5308cf7640fbeae405c586849357fb16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1677c018dc4ea325a595a96c899b5b1ea25e2880ae905e4ef867805bc1f3f2b4601522ca0528e0b8743ce7d5f2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdcba0fb819732e04beafd24077bc73fd068250a5bbc56f432ce0e75e3cbbb9ff16fde54b29671bf49f31744cb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7b3ba447187790c7e84326dbbe4a9e6fa62b90a2a154822142a671cd3dc7a12d3302ee0021e118664a6117a59;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2bf640cb7e2115f356199fad1ac4417dc66bf15071a534a82b334a5364589ae91b66974e5152c2c921c9f3fc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65501f13dd94f7f583ceb9538f88c8111e34131ca6e3d8a9e390df4910557da2396f016ca33b05583fb1f53608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'habbbf874768612d57884f7eeb7d34210b2e19808017452e91a1f429d8bfa313b6460f54415d250ae2cd244d6aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159d615654155b66d0740382e52ab31d311972da00657a29817dce9af6e793b872d28995b24750f49f6177f9a3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b4389155063d7c98fbffec19da9893f37f7e61b6fe37b4b05f96cf65f84e4a9b190c5f5ebb30a1ae6d3450ea7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3287a383f89619abccc275444aae9a47d88d6175b3414b7720163a71f0fff313ee3cf8cf2e10135e95a622b3ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67df331c456d0e599877035597212887bdbff02c18e28a73af1d77c3f8bf6162f78433224dd408909f2ab305ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135631924b69c153c443e0a0e6f837e524b5bcd7a853833b39e8a1d29616c41ad3e0a2c43ec51d07c4249e590ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d271b94dddc57814a7ecb68fa27f5db2affdd697819218103fc44bd0467c3e20b18a2947beb7207c8a50aa3df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b113717a0b34f89d84698b9c98305fdfc436ce4d3e4228bfed2384d9602b35058a4be292b32f3c7b16bc7b4bb8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac6789d0ba9e29c7b17e9a328c9f900a3e422367c99e5e98f6d8054edbb6a3b6e5f0459aaeb6df024c90bfdf57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11883cfd7c64d5f1afaa131bfd2af4665467f51f2e237299888784be0618c24f0e59278ba464a000c64829ee390;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff43cdcdd25885ec0835593a626a2236cb7e745f36fae972630c05dfffd4965750a0a3bca9217758afe7879d66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd6a4836778425f9220dc4bbfbf58e9c79d20e93ad54f634910527ffed07ee96e4c2506138dd740d7f851366ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188275d0fcefd162bfabaca4651f6d076b66b61b2cbe4d7956a22bdf476778efc5960c98e193632c26173a865af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98b5e600d89d47b578a3a9dead01518ee2b7ab520c07692033a8507bb72c7de79021df9129af7b54294a065134;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4866c75a930ec83a3e667cd268a35fc7e7f78d3834c2d6b44271791e65ae543b25009f59c9eaa9f494f0edff7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h425e18cfa5799dd359e93b67ab71b485a41242e57faef7527ce7f59f26dfa4b924fd093f805d4026e86092245d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd20a1ad68bc079a69fc22a43aa9acfbbc05c1466b1db43930bc8ecf8b23a4dfb463042c89b96e5b634272fbeec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53b6cf5e942649182d67d7bd64300ea428366142930db1999d26cd162a7a32a0550327a6c46723bc9f26856fbc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h643292eb54d36efb337b5f7bd35e46d251a0f05b087be8a72c429e0ffb24ebb2e8fdfb7c4eb2527b4973543e6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41917050cee1f284361052a53e8eedc678a863870c5ba35234b58ec66c6e56706edf33a71b96d40704cc89db35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9323e1571266a67077992e80e5974743539c2614bafc97a49c205678a0811539b315fa33ef336c81248c1fb44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdef57c6de91e2fc11c1c8fc90764731d92537e468244ca8a1bedcf3e506ca6bb0fe08ec1fc45a5037283e29b37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15713e75052d84dc95b1e238b9f47a1f22df00c5b84982d764977012353cc794e25f16f142a80fb4512a297f122;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5c0d6a74cb9f4622a3741bd931b753f3ff7442e07bbc700c16dfc5659a38a82fa8a4634a6fbb0db651dd90dde;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b78c6af6e10a7df387a450b8b32288c232265de46bb94e5481241fe6347c4bfbcdc07a6100bdb614fcf8185272;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117caf84d6cc67f1ab54fa4ec1c5d8c9634467146190ef201efcb6f3a5602826179a9c16fa7a1e0e7832dbe7621;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bccca28a55911b5bad0c70c73b8b4d67def4cb6188e4beca83b42e0109cb3869c026b4dff01a3a672adc30ad5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c06a583f10ed1df5edc3a54c55c5e1854d9966484f936ee0a297af321e37e5c658bfb189ad6671d14d663fe0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e055177a82509ced0137ddbe5c0249c4e587a0fa36569798bd8ceeec5f7e8301a6b5b5f9d44f50997303685177;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d799f12d95ae251695eeec263f87a626492b8e048e094a0b6c8a827a3f650145184c0e2089553abb462956dc4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7e8d124c263c4a0f353256f7b33a42d5004acfa32189505a4dc087a624e11a21b64391bc3d3702378f1ca5c60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc20bdb47787b7a0e04b289d0d1227ef29304c172b2817c16e348d031d8d71d439ee067a0f74d99a8581711a993;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d74040f638985a1dcc7ad4b5f73859b5651886e1966da4414aa8185677d8366b1cef593d3388089b539a4e91fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f91a11174a41b5860257442ec4ab955fc9522a7b752f5916940b90fffbfd69d5f60c6b495fd340db26205b24b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49be1adc82e95ec76fbb9c87ae5e418e255dca028a8c363f1286ada36c3557a27629aa3e831e0299f9887e222d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he18a1993d727d74d3763ff52a1d4a1a56c99c28d84367f6cd1f22406be35ea60f5fb7dee0b9deffec1f6ece052;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aafcc49b52c5df5d026ee266bf42a0ae6d7040a7ebd19c0e215c50dec8aaee21062f0fc244826347846d1206a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa45596072ef01b955b4aac46d7874ec3d8912e275e85f10047af08a3d0ec7c495e41a47a29fe5393481661f5a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2b0f54da33dc4b0031fdfab170225a38e8261f4fe11fa6df5d78eda80ae27c41bbb1f31f8e24f971350078325;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6df074ac78dd0e6184fb48e16e653a08b1b2daadcf0e113a996f086d73a34e969834ac8b7cdbc9733defa9135;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119e430d325342e9b979c56cd566be29bd40f20da2fe045d83c607174694fbc17f76b76034db71c6540114dd034;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he17f0f0d43419e16a1a6fcee2c41d6e5b5081fcf1f235aa90db9bc5450f618e3c699e106524f10fab601e8a763;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf051df5a65e5f852f23e089fb01e56538ef1d144b4e91c7ecb0ef69b949a7e8c16f2b379810bce3778db7ee61b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71a3bcdab18c880e928fa25035b103a9d010dcd08b16ce979dd0e23eba3dae42f008b1b2785b41ddceb3eeed1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17086173398b5ff8c0823df9a34f25ad690e981b49548ffc0024b1e3ca50ab05da119cf5f3257af4c40741671ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18792f8b73ac2410d776f57382794587e6dcc86fea196328062fa59e53fb6c6b45e678afd7b55b72e5b76eb74fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h942d0e16ae0bdb6139efc3b03902ea501d6ceaf54df4b302b12c0a66b4b3d49bd97ce991e3701e29c9f1655054;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha795778b497b9a99f0b901b4785e21c895b70a14cd9aba80689ce53b60c4738ced48263ec9584a31761d993ded;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6189a54e948c02a29c81b66800a0fe6aad3eb7fee8c9b40968f8bf33cad6146f9688248514c8fa37131fd1d19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17aef0bb875c24a025aaa4109e964f4196895ec31ccaeeb9b0c35f9b84bed57ef66d3aff3b31f68e78ae8846fd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a1cf6dc25df18e0791d0f9b324b66d96f4f67740889f5c3c4517ae38090bbcdad26322e34e7a08f8fa0e3f635;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ded5cc15411316ba0351854b63a59d577bdf9b8a365cd36270b5d83c4e0bc63ce71260f8e875befdc54edac2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1460c7e4672e6d772e29593cde360f0a752f85d6dd1c3f8ddc993bef8da95ed74d6618b72e9232bc047088a4ab8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95761df084a0c5e798b17d83ef4a0d3acbb8ae7ab4b5dd9df43a9d95853437dfa91eb137c43daffa26c90fe9a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9312af3f2068e82ad17ce0a3340a86ceace58ba0b503addd6adf2d89cddc8deb4e8bfa6b255d003abc88f649a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19374a96751472b26b0b707466d6161d9f17ad99dedfcf7469f228d2fb8f2abd5470ff66ba97a7c2bcc3f8d5da4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2e9a1b127794793102c14d22fee9706bb130f17c3c0b727864ef4c7e7aa66f4a6be5233e028edf251e4788df3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185a75c856f4159b2ef5513501aa5270597eb172851d88eac41ce84e6762637ce8834bd93ab4089eaf0a60ecaf0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bbe72d9808a59ab58f47fdc14e8a14bf2c426310784b1cc12578584bd9c32a88e533afa805f143e8538afbf61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb399e1f2aced8ac8b41e4bd06ab1223a00963e44d069187e053340b10be23ff7a61e89ee5b1770708b11e6dfc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b74c40009af1d5ce0310ff663fee165b016dbdeca5d6bfa1c4c2ecb2c8c3e0bf7c4a90584afdc7a7420a04720a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1411a4805393e8f7c1babbcb020d5aac5d3ae62500186cf021c73ffe7824b4c3645233eabfbef07ab3167fe0e1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h237977500527e575a4f256288e11960d923b6746ee4e19e87dc6716d8c38049af7248debd348fd277cb52d1521;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h687eacbcff443cf4d06a021f215624be3a9e0c42817053046e85ef291651980b62624fe33fa0f5a47b64f83908;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefd59eb21d02fc576284512c4a98275cd51f527d7a5dccab35580d6bf5687f6839c7393e94720ff27b10578e07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f825ebbc3fc6539de83ee1882c9c71a2c38bf1fe3485664158ea3a7c6de84dd01b44cbff6ea6deb6ff0a3c144;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff4c541826ed159369f8b62ae9f2feec374b6d42aae0469c685061c74ca9bea0c0036927027003b71928083323;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0951d429c37bbfc5e3531c6152c7f9521e7f02c6577e1aa2a06301780c5f48b36f61da9c09c8e595e9ae2277;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb120db3a1817f8cda67a413ae5e986cc6174a7760bad8ef034c47bb3b8f30f722c25524b5212feb64b305e6eb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192d71c10e8504d23d2b09638af2a73e72b54dc4cbe201ed5443ae3f8b488d5b6adad6b4b2f9546552e5d9e871;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7513251049dacb3461dad26ba2487a248af8040225373c208faaa1bf82f3766070e585721c333c81171ef5193;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec287a4a9f15a4394ca8557a09700665dfea61e3747d406f2e1b3939431c63f6844d2c21b5dc5291f27fa68d9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c47643363b382a27e00c3171345b9fe5128c2a2573c10136df54ef9bee21a31f1353a13a8a35ba4bc010d4e3c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27f116f67559d35e0b1fd1e6287dbe16c7df3fa80facd9124e3aaa14303ed2220649007772254bf37c7b272445;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3fb9bbf8bd9349caa347733b5ccba0034a439f9a0fb89b7c256982fb51f4bc9b2d4f44b11e443e1745b1d2f51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e9bec457a110805bcca8c32100372f0047e7fa6917e2acde9d9d77ca3f3b77c7f0b82f4da31d986f6287f109d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acdf05a815b5850746f05e69b0ed8553d6ba490339c0f2794404b64b57ac87de335254514b730c1562e2311fc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ad93bcc4b901adca42307e83cd38f11885237b9091f4bbab3045fd77f98976d1253c83f2966e782d9c96c8e52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hedc2a892c86cc6b5bcc4e3c82520bc8f48ff387d0a8a1fa6e279e2c2b4a17f3260877fc3476cdc7ee03bc8249a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1778774b63abb0f499015811dcd9fcfa52425c9cee18f6f320d2d9276d1dcd42f9380f99613f456bbf431f76cf2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84d65a94dcec0c52a90c137421060e0ed43d0fa8595fb9d472cdb53f4f06fcde565d89bbe211bf2ca83df7ec25;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18284f745db4a532bfcd1d791c0a79ac80fd778c30ea43cef61776f11e9b25bdb9417f65d98070c65a472197b38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac348259be2861c6844a112ed6297a32387819269d7ba17d9d4c309835bad90263ec02be5d19a501f329f3eb0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e14af133034f3ddc3a3de4be5d8137609d3b0d3895bf40d2b07da799a666fee2953cad18f23c300ee30896665a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b7fefb560792a2e8b20ba2a5c650abbca28e1c160e4e86d9298c8efb28aa157f974a2bfb11c11ac98540ed54b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef4cf87e504db65b735f6d1d97f4b6437b43e40cfb30f371b3dcd66938a1957639fd8e9554533aa50f7071eacb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbab6412f8fb54feff5d7827d15e557a78d51c6af52eaf7006f6f887b1d9e82ce1b21a33ed542506f4f139ef9be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebdeb1497f90e0d4586a799408b16deec8f502973e810d4f48c6561d88f96d93e6af769173923d5874de5ff092;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52b2fe2e6ce80ebc65049c733f156ce203af8ad040fc93c7eaea8a304169dfd53ca0ce9bcc0c9feacf4fbf1f56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1042750f070c7da873f15ce99be26897db9a6fa6d9f4e361e22806af2ccd3e783ccf2e1bdc749f88bde3786842e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1f85d46410dbd3827d2cba476fe9bd93d9f5a2dfaabd53b2c0406c2f503b8f2bc339615f34bd7371e24edba79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c408668d8c249fe937dfff3a1fafa43fa716cadff75476cca07bc8e88392759bf99422c35188c7df4012991f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1334a8e54277d6b3c46627e3416c104c0f3b5dabe63de14ca74a3be79e8da5cf62b509e6fffc8398ec6827b82a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39bc2c8d5fcb61f62a7d5fa578d8d4cb91cc26b27473c379237d1508a16aeb83ab7c75ac0695e4d980c86196f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed1d0f5be41621ade0a71d8438c132ff3625c5c115c0cacc3bb3be0cb92ed615f5043e8addfc9001219916a50d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8961b5c1374eda2d344ee977a8058b6369c883fa9e56d8e27e81cd92b035ce48c7e38fa613cde822c782b9ea3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d87b7d2f3c4678328b4e65a128a44f5d6ace1fd97b690ca5335ccb792d07826296fe133f95f123026502a2a6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14179535a42b9c4fa10da938206501916a03aee3e52a66d6454444084758c3b8f415691e584c0b5627b8872a2bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3321e46dcf4cf3550c4af3c17628032bd4b2f98a16a178b56ad064c5bdc0c346cabb771092e2e99097c9d1bfa3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e1907a170e7ff49881a7636e43f6eb96ba09562895920a88b89a704cd331b400cdfae3ec58d00626d530ec14c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62b62b53b8f4081ac94e24488a401baab90c19dc8cedf799e65979f00f18e0c8720be581c55f95dea92355bb3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b23f8bd2b89915e0779bb760c7a86e112f148008e0c11cd7141f3f1ea61c64af5680d1c26628b985418a9dffc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha418f61836a650edfc207677a94e9abf9376b2d931aa6a39313362c8fa3a69e47bf388708ba2b12f923168620;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ad01f2f11dd1bcb28e9f2a5b3173f9f1cc52ead2bc4947c2552fb91f386ac9c58f5e343cd83d10c43fb0a1bd3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a520364d7679f29f055fabdbb55616fe087791e6785c001fe39eb282eb009931e08db6988b6c56d39c2fe94e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd406d0868b06bf3a4de9363ea8bf3c2942fe307672113147b80ec73a922b4edf66d1471f0c840bd731d3e86588;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e48f864f26683a30f7f87fbd600af3b8749fc2a0267cb0a7644b1d8e069212a862f8f6c4274d2e079a29ebd27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6109cc89d35386139b3d78f106d0f6370a2000238842f52cdec651cd0449905320345846bd9bea35a6ad536bee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6fd45ec202c07a25f62dc3720f977300f907b42f594c048966fce307554459dd20f6c1e163b6cbff0daa358463;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd32b1d94774cec4a87c2ad6d01a5526051ca7e966de85eb04d5ca1e02146dc28926139f5bca653931876fd86d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14711b4b19d27814746563976e354e96b841f22d2b5b6d6d1c16aac466a7d8e34e4ce998fb998b22a2e6d1f2cb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e4b73d0fdd8b47ae672e4b54cb5fe3ac6552975f8380d2ee321e8d85ffe3f93589635f8db852d5db8a98aa632;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2e3fa56e4cee7121d3f99c2df01b9b7e9a06192cd1df6828a214c97a151b34ee3e753509fcc57ec20d50501a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h412a293b2f7957f5ead093a4695c2b6716ac86a8c030cbff8d59403423c367ff95336602cf211954a925c761c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54d5efe21cf248e9efbcb8c80a908199e90d507a81e6e5057cb843cf253a8f0727feb3b0a7b1fe6aaf4261c168;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd98a120f383e5a38633d94403e31994815c36ee71b3fbb340b748e4aa32edbfb23e5c3b76a3cfc029a11065a0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a7c55e7e6de4c1768a8cb9013ffdb9284dc16431d8f900fc4ad87f66cd8239fe444252bd793d63ed799a6f50c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b92c759aa6add43ded82e8a8e2f1c358ddbefe0411d9daf904856367460075c6de5bfab3282617a3050cc2b98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119a7eed061e8b82eda108b775131e1c76d2f761846ad0eb6348a6b48ab5131319c389c4001afbff143f5a51674;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aaf59555744c23d4f7a5e58c65cd00c4c8effe5d8b4635c175967d27d313aba017c574e55e91f2f45ac00299f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h716083c62c082ee43f124b21d1e2fc9746cae3dcfc2eaefbe88dc8402eaf7197dae1d559ae137e2b82736e6fef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a6cd24fd3fc489057ccbc956ce753f3e1926477ac71a7b5042661229cdad9fa7b137de7d23b6420f7b86bc23e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf462d5dee28a377049cfbcb50767ffc6a30bf93bd235838c8041ba38e814cb6aee89bcce63da7194c47ea85ea1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16d9c62fa7293aa7e22f378ed47650c229c4516b85a517d248382e92902b737ddde9e363f26447d192b3f48dc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h351cd481f035cf488ee15c587936388fb5b00ca439c22aba1c02dbc64024dce266f7521b2e10381b4dd28cffcf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h786e67ef4248d237d47bfb09ad998f884bdffac198056b7255998a0cb6595884e7417afccc054d9e0b0c106fdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71177fe3afc0a70879672077b52dbb6682c2dd0f59f1a0bcc9ad2ee341c859f6add33a9962fb372cfbece55033;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d3055906051b2534188689014663372aba7ba1ac514075e977ef6beb0157b3dc5f9bc581fd548231633ea9dc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h414128f8787642045a62250a7950ac8ce82ddbfc6807b5d429713c2cb36a08f959de346899418202ad035cb2ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8008e49c178a8b32a167e98be10e71201cdebd9db10695498bcee4f00902fedd508b4ce16fc8350da1a5db045;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ab484f89721bb27cfce84cea7aab9a684ed591b7f5b708ea0dceecfdc2a36bc5cfbfa1dbf2d049ced24070121;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f094cdad87012ab16bf04ad4ca007cc018b922c25f7786922dd79840be65ee016aad626ce6743c4c7cd0329d17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb685b6f68ece9c8b30a1f60ae12d53c6af9d2a24e315e828db69204ed2ab9c661c73e58ac2b8ac3acd8d767e32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54e67d116c88c8930839949eaaa77890855f4d3d71fa68d567e88c1b58304df661134c95506ce3f9d305f6dc69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h177bac0848052260148500ca28087a2522ae53713374c7eee46e87cd9846edd38d476ea584b3a0158e3083bc3f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da56d1d1aded0568d3bcdd6f5133e01b2d4163bd3f672ed003f251801742aab70243aded99c49394910f565478;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf45d143b3e2d8d78374372ff855e10994fd6fd7caf4652a567a29cd3a4473424f93fbd37562163a05fdf4ab15;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3351757964ef9180f85491a143eadbdc297d3356297f24e862e50d51b6f188db795b9d51390b82199d4dedd04f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e85c4399291c7787289ff1f07eb5e905318eed6ace5aa6fe6c4d1ed3af06c4b7d3db705cfc8f93d6d60b58594;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182ca7f57f9f590431ffa67f67b71438acd65c623820db292c7a71cb38fa285ceb2516479536a5150718a99d8bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159c4864dc8bbf877d84456182b292dcebc35f4707414e9f09deca9d5b0ef6463782deea5cce21e7db2d05c079a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161056803c640a055b81e95a8cc879b39e8298e9c756eb571aee0b99aad5da4de294060b921ac4e1a6dfdff3cf1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bd91c4846d1090199b38851b9416b1ec9eeded8bd8bb0399353a1df514dcf30d12924a067a28c304fc896c8d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115210b71bae4fa9c0a36dd19cb1e0f3b4b2bf9a3d05c04faa62a68eb319bcfef188447b944b41f41d15184121f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d495554d4001e099d9fb620609ee34659d3f01660a2d7648e53547399df3b8b3637682aab4be6af5feda21544;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d781e8371091854307033d90aaf6c7dddb8a3c30b59f9b93983044ac2bc63f60a795326cce3944e5fcd359f97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c31bc28d57a0dce4853fe720f4be66842e01ade6f42e2c4b939c1671119e7772710558774156ab2e100efa18f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf8a0f341d4fc94bad21e6d68fc1cf5448aa56489c3cc7138dede773d55fb1942be957b38bfba3da84b4d005d5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d68b528a99b57d20cdb9f381bbc880cdb184006e1f59fe183ca1cdae7a609d7411332d5efc1ded561195c3501;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf46a3db8d5861c5c93a459266a33935a4cbe0b583ad59a31a99f473a9459d2ae9999720ea4cb606c099ec26b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132973eacc1fa33ae8824add6aa026b4a63bdeed904c19f248dfd5243fdc28ce90e118108d702b2376e296414e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7f2d65a314fb017cf2ee8adb6998870c2743544d267bd3d8a8486b763679e256aa85475393f2c0559b2b97de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9cff72b0d992ad016a2c7beafe90b17fc0a0263779c49afcacf6e3ba3620f742aef0bd57066038418c57fa7da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0484e6e598ac5b62293fe27bcfc18d2c17542676dbc4cb5dbd54028556ff019035bace53b7c05599093ea6ec3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f99f5e1cc85202bad7bb757c4d6f664ea8965f9bf9be11843d7f653261790396042521ef37754456c96a263b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e1c22d2402392e515125d764c3c0194e6bc391ee358f2e83fd50fff9eb1a10c964ecdf4cb68957db8e7984538;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172bbbe3dfefa9b78347c5d0db95f5b917ff4ba5d70081bd34b4c4afe005094d40a73b0f83d3ccadc378628128a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdf2a305f65fb69810d04c6e900de42c311d7248254a9d8d53bb7e9d81f469df41656716ce68f64d23f77ef088;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4224b78dc5cf989e59cd5bee24f49ea7c74657cf1334ac912468d7e9bec503ddfa7ef66b620e84fb88e41bc3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4156bcc4729c418856dc6b8feac63dbcee86d2404263c5ba5ee0fd726f0867bcfe63d8699d9adcccf9659ea38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41c5e978d72c7c9bc54ab5673362dfa32a8bea387882b85e0b72e877c2692e926d1f1efbd2d1f6cc151bf92bdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c4034ad9992ae706d0b518e69757ede5f6e873ac95e23dc5ceb54cb1fbeb96b1b027c7dce232a87d559272aeeb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4038a1bf7081546c66f453748de08722cb133f7dba46714e8d4e90c1d9cec75f4a434d7001b02f54c776f99884;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148af791505714a04334af782279799f5b8b876ce8c32dfafd6113d8d05b95644cec7053c73e8cf0798fc656615;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10fee51b7a682122a3f8a148ad3a6aecbe6fd5f1df1a4f4d5fc67a2f5ae8aa2b924f0b33c016c6226ffe88dfe03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58ba1e8fb816fb1167e3ff9773a9330cf893e59216819f8f60fdaee6a804b6ef3c87ca92e40bc4dcd2924275a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d5d5ff976d6cf5abd83197030b75ffe6d6a1260a3936da17f5ccda28c71d40f986347e74bc689f7312e9d7953;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a1344ac0442087ae6e9e1117880bb83800093b4ef917e9110e2d9f02d7f7afebb370c958ebd6a480718580343;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h802770fb1e6ebb0bbfe1d4009b1cf689357eca875d8d7a817c722bc6d34335fdfc53e44365eb2cd0d584142ee7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70c97aa8cbe474718f80b35800358ddf7f14cfe894debbe37158e5eacc6211262142559872aea549e35f70c86d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d212cab0dc5f0089eb0cc9c1393ab5a2adc7b21eff3f7cb9319ec5edc0b9d30d90cb3abfff33b4a62ab8ce7e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a4c2c050673a4752b9bf1c47c0c7c9a586fd8f2c4f39454809413dd16e00e5230af74d2d2453a4de6aadea7b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0078cf11efbaddfd2a1b219b2f86c2c338fc68c0047c4fa2610b82f9d68014f3f2263a9fc335dd9e25fefc85e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b06b6fa753ccd2b0e25eadc465ec923ed631e1b4d598f486d5339e1490081a1c5e3a62d4a5b6c302ed8804760a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d27fee9e5a9ad08187c7c18f0147486507616cd43769e58fd1bea56786d1af113aa61c532bf6d52c65c738239;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80d63088b57f44055399337d29f8b3483507d79ff6105ee8ab1f64a34e0210068ec262925a7d1f69de99037c31;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ecd6f00de8c0d249aa1978dc5ef6ba3e839e8104a8260c5a7d350d14d57ff40e1b84d669285d09c43ade626af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173afa0d852652c867f59aecada4ca5e0505e497eb5ed0110a7dc423f3008422a4664e394429df7b26ce4b984b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8c73b93a02ea809be653facdcf549a09cac716536b29175f71a99e4bc21a3df30e4400da3ec56044dbf9bcc49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h769aecf757778b5632daed1a45c626db8ece1480281ad51def31971b9b4e92a0ef90b301e1fe16afdd6adc8d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1742ebce0e18cf08db03492366667a65bbe5cce90290458cd8b30af28e1dbc8fce9e0b2ce81d4b0aa0b7ff64b97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc2e9a034f1423fec15e532518686b5f0e115e42a878f1adaf71bfa6f742f7c883ee24144b9617ff5141cbd3ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1276f5382e16543296cf4dc45783c1124774c67bbb8e24ba369d830a07c1bc573e447c995230ff82095de14f470;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c81a12fa5fbda87f74d0b8cb156d0dc28b367290e08f7963fba80469b2ecf44af686f9a73c6f429aa75b825d89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbea91434fef02e153dd9d37f3af171df5273a346e3ff38f14537aac6503cc1ecafb266f626186667fa874c39f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3284fb1b8af441a444137d55f55a4ae801502c6acfac76148acf7d9009d9602c5f485919632a82a8160abe3d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d795c8f4798bd9e07d5add3cbc4387863bfd24a6904d0be45eabf76604e3bb77b94a241bbafb989369e5d4cb5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8cd6964b008dcc047fb5319c9a7a18f861702d5fb2600f7acb891f397a90a2230f535c9b56f7b480305cd9c94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf44dc9944ef541744876280c7ae38e9d0cc02dfd00eb62272170153ef2a492d374fa8134d2cfcfa57dc9e8761;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13fa44dc3b317857068e883c2ead85c2687360120a5cd8a3a313ff20b463959842c5f729fc15a2cb0ee7bb00159;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc576c170ba2878ce59a55d6d0d86b885bf6ffdcfb849eff54854b2a9ab4d8ac553c8f01bfc605aa5491b429a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7a6b857b728e45d633f785fe996dd9c47eea89fa0c2053f3ddff275af501106d2257d70182fb99f9fca18f6a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88dc3ffc013f0886e1c8b5e91d5e3d12ba58b4e30a56655dbd466468c4caf27af4f4e046f4492ce19318af0566;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce7c389109678df9458a6741dc674a7d2ab7acb693eeca628ad117617ab9657fbe0918add604db1a94b3bd4a93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e902b3881dd725b010e3e064000b37d76a1522f78826e1c3c016aa051bcceff2d32923980dfcabacb0b2571de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d15ab8ae3de7521dd635263fed28987d20a690478bf66a7ddaa35704a12e67e7ea3d012dc6952ba2e88e5f37dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h723d13d8a9e07e1b13e32c71306b474eba17f5cbf7e71ab451f8add469c93b97a36525ecd7fee5f3e20f3a5212;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d8145a4c824d42503323859dfa42d797d5c6fe58732d6500089f56013ebfe60b36ebc3ba238adf536ad25ec7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a9965e4ceb15da9ef1d7eec4216a6cb2fcc6b31dd45f0feb4a2eb163afb228b229df43a9e45b4b5caebf42d87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc81c40623c0befd74873d235f078af3de49d3b6ed4f110f77820f9f35765aae3ede50643deb0589beabd84eca5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a784c428323a4b0d2b6c51963d85ee6442b655428e8cd67987b66bbdd79254a845e79fce03f63b85924a81aad4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6ff9e7d0d0baa6413e04f0b219a8d4966da71456ffcf1677db2de9b9a5700068b48e6d2ac07e4f51d08135fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ceadc6a738a754c438ad6a5fd1727ef917a248c2a941007181d6f2e4c74a26d447625ac95f7b7792e31fded7bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f79b8ee80e836020defff1534ba65c6485f856486e40cf3fbd66928b42525173ca50c47b6f6edf72254b00f6d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da0447182d714c9e75a3be2ce31ea89123b5abf504906dab3522bc94c9afc5ef942703170555e49925cea033ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28e271d674b51900b6891834789b3c115bcf0503843207beff572b76f9e03fac904b76c6dacc6e010299216c0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3de4f31d5a4b075df906e52c8a6e5d6835b5a67adc7f041d51740e6d68187a22404b4a6fa3ca6f75c763ebbb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d50556c6bc3e7d428c9b83423602adf68f7316e473746384b18fc21af4e6760af45c061da450698679f9581b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32ff4d18d6734b83255f81df9dc9ea06c7a522c5b85e7d4f72466dc3154b78993a4491df684b8db39a212ff4d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h833dc718ef6c70004a0cbe87ca0437e40988b9b15e52a0b4a80a391bf766d845d88eba597e9d590c3c39eb9af8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf6ed5992f1aad60cebc6ead16c8a4b06fc195eab61b073a76af17456b504f96831d5553d4ac8c772660b05856;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a00cde30078f6d3f8930ea8e0edace0acaf64929b321e6ff293a52e43945acb8eb6a0782ecdfe419213dbc965;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bdfece448b5beaae4d00ec339f31283168bb79492675066a96a4790cfedab591904830c3423e70d2513b968c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a72b803dd02c54d0a1e431863371b2f10e4afed71b7584b754ab6426105b3f2f49e642f033600a6148e8d49718;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac68a66743979ee5bd9fec3c126b97dbf2e1662ff1aaefa0c80552a50698683ff50a1c1a3b6ffe054671a7421c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4aea80d24766cff2fb138762b5561c9bf129c7a7ea807f8929ef4184629754311ac733e378a5379097bda164a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcda5935ef738b4cecd4482bf3518ff18b7b9f108c464b469ab738f86880aa7c6be09b9f705e6c1fc8b8070b652;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h390daba99c301a533a56915038af56a990a2cf078c40ba6b8130acceb5977383f76ff210c2205bcaea09e8a7a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35faf3d7d520fe4b67889d1ddf755c3e26915d676cea8a488f87b1d6bd33753870e3ada3af78c3c3a446b7d649;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f543406eb9c939a18a162cba4b9aa7b01b741ce575cbcdcd2f98c76649b2cd702cc4a54199c0d016dd89eb173a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9c88463a77ccd2c1db052b3c5da65892825fdcc6c39030bd09959058641c0d3dba39392d0cb443748993493db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148767850f5ba9d8241463c8e5394d4f7c9202bb68643ea570b22fad20128f29a056d738d5d4a600217221c1ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14714ba9202d86953a82a30e1ea6279e7a77fa2a752c84f09dd7bc2877096bda70f888a43031d8a9456160637db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56d6f68a265f2b5bad5b6db0c409d10e13f1cf4822fb94d14a8a5bf4389f192b9b8695f7bfda9929aaf9b48850;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf99ce658c3dceee78d878dc1779246ced3d41963939a671ea6b9e52c72100614c4335cf982414e8d25f9e93e6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5497d5fe090f865004592b7eeb5b4966752ee706d0ac5a9be61d4a6df9aab621203493f8d5eb76df0af25f84a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf371299db782cbc9ba70b86719a6f349647355e01eb8db1d6e85ca8492d4fd7abe8d6579881487e44f19298892;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6417be7403b5cad9a6b3e86caae74c3b1848453e68e60451663af25536b41801f9cd47380ed982ad22b57d0d94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffef7f62aab9f4b9eb2b039fb4a867db9a951c0413459d5ba5783822667f27e2f1e6387612f5cf8ac2d2386e32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d39fd94e9355af6455ad15a4b5ceae85d3f6941eca669cce78c22a690bddbdf3d02d47afeda8b9ad866cb0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10cade509881b527fcdbb90b6e319e3a46e932a3b78b3f32dae0b614340f1434b1d9bfa7e99d85b35765d50fb8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c17cbafc34195adddbb390113cd5c70e728c9a2d03b90feb2289f0fa577afb33f05e66475fde93b1855529775;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75e5b8310bb23f4f9ac21ad8ac3cb0fba5828e14f52c0ed9b685a5097af1796b441b704a6ec91416360977344e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be10cbebf82dd09143fe2eb006cf03b3123b7db43e42126af1379c730aa58db5bffdbdcae210518e08470b83f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h451134fe6871cbb0b467a311b24937e3009a817039c3b704c51b1309fa74dfc65ddf075263a88e5ceaa334f9e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fab8983a4fc651e5888e49eb405d40d79581ecc6cf98de82d3c89510fb7a26d0cb6ef6230c38acdff7f62b2a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77b93b0295572d4c8b2a7cb1b359b9244a7fd716bb72bad29f8064febc417959e05bac2f565eee0f0a73960035;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6ab93f0d199cd98889dcfecbfe894bb239f8421d165f3c64d904a835914247a5cc28e383dc5d19cbd40514f2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf25428410362f7a990eb12a80e566bd1767dd939e322deb270140e8e443f23f23cdd113a90fd9389eeab06de37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa49cdc7750f16480a7deeadabace29339389b087c566bd774f73a9cdb6f146fbade2822a577753b1191706769;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3166367e4ee95ef8b3d58babee2f78043e704d732c6380021309e3a16829e027b85fe103994b264055874cf87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7da9ae4f1e0d2accbc615aeee4f65ab7dc75d09948adee0b394b6a9e71bad783403b9a610dd795692d465c1ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h204dad8e2db8c0d683a3935a7bbb57dff5eab28d74ff8619a57cf4123bbfffd948500ef370995dce6c82ee52e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1282fcbfb2cf527944ff1400e00978a0fe5b6c48a3c2239930eeb829d35e19234d041d553b11d5f616e8af68a46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4edf69d2134d81f3e447146977efc5fbadeda804932db9e81532ee091bfc84195af5fae06396a24c4e9d554891;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13777a5ef85b721623483e17a69e7ebf8ddf25abf2c6f8bce2337a8ee77d598322c975f9fa944a7ce2d681de8b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e47f34d329cd5348fb0103c2102a5bd54052279857a4ec592a9e0c55146724dcc02f2ace459ae66bbafe398893;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5750b3c9d491f2dbbe814240fafc43daa3a62a15188df4232b93460d9b56e309795edad2ea9f72afb2a808c21c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0aa2c8acb0d27d591641876efa9e31024d0668b473dbc7c59fe71385de411a4532d49d94eaa8763f03198cce7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he436ef0788fe7a42e5662afc7aef3a4f4c4dfb0ada9df041b81eb5eb52f5187fa5856763abdbafecdae1eaa3b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf241b70d93f0124875382d312099d146db67c5bf7cdb3585e80ccfb97d70e119fd7039ddcd2a4bb47edc78e1ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bcd62a49fc57f77f4802664277810d8d429097ff4e769e5ccc464276f2329792e13af71a446ee029c43067ea5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f1410e2d1182cf11089dbb3e6f74ae6c8d81d59256525786ef27cd0f70b6a198de84906081851eca753faa18a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he18cb27166c1457cd7ec326ae1fe523c31bc62d870eb0d19a3b49a2f9f63f206ca48a8a79b955af992b8e45a1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186f92273a62d9ab299eff6622b1fc19cd088dc650dd43f0794c898a0454c310d98469d70fe6f2154185f823917;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1516b1c68c37220a130d239598f19af131a4346d14f51cb48d2b013ce1fc47af07227ace57689533ff3fc905a3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24e585e61ab4006bd392a1cf6ae810e19a1c62a4458fe1a9bfafe27effe05d3ef0a1a72b80e834829af82b3e71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h977a0f740b5a2075e19ef040d3be60b34403e20a2e9224cf6c3263de5318c041b265882838aea6b406ce66bfd5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5604893fe587d723eef9b304d6086da00b4adc6ef397df05de51c21ce4881cbaf18054856b22868199e0540c2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2154af8c56c79b64965931dd48032e4468052cfbdec681baa94f6e46eebd93dfe0411b5e35d10d1815fc0b553;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4459148b1424a38f7c8b507a44629dbfd8add03db49e9b6624fa612b7262ef7c44365aed440b26971ebb5c855d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1826c95f3db2b4d3c091c81fcda359b550fb1cdf08558bec3644f2eae35d39b1884061941139757c09bdeb3bec8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175a349b1bf83d9fd5239bab9a2b3de527348f27390690bb3d734f5e889331a95ed0ef44c928089c02ea8a91262;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1824fed9361fdc9d54f911166a38bafc4ad2ba539d0ea0c15977398aad91a56c7c4ff9b83470c9bfca50228ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1500d4876ae85e2f0951b0f4be96f683cf7b047c38be2573223c88b92edb94830fd310a579d3aa9aab4d18d7668;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18aa62d3d2f499f0c4099d8070e384e66a661ee8644b9f2c874e58889cea1e46117bfa89e72f1ee0e3b0f70dcbf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65e7c69cfab4d960452442cab5beeca78b9fc25446c8138b64008f8d326c37650e2569e0c6947b9ab5afb539a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28e4dced2a9a038ad4b4d77d0addf50ecf2d6fb6f200df65fa460123fdab3f36ed74f1c3faf9be07c625f71a8b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h968e0f7860f981eb2f1feb2277b733a6e402779bd108caee5f4b9c8a8abd530e988ab9a7c84a4648004206e0e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d292304d55877fbc5c52380e9d276b4c20a94da466b52799021e18e617ba03b449f7847c1247344ff72dc131db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a256d7152db4adbf1b41b44770d05a38233f75e82cf2bde1ba87c72ef63486c5d2a7200a8743153376fe655b29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a49960e15f4172fedcd387ed4e90568300749643c6749fea7eb62cdc2a8c3aac6a77937e7b2c319aa46c33b673;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7ebb3bbd37b522e091f85ecaee432d42aeeb4a04534ba1e4f42ae8522317063254304ef06301a8d867aff62dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c1be00b1732f77ebc41b40facc905ecd291a2ebf8fcfdd24eb7b5778040839377136066b988511cde10bc8758;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1734b249a1fa2036e611baf70976b9e520d65974b87e18cbf0323f7add27a6068c04bec90f98cbe1f0e68e47e27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d00eb45cfeafcc6d7182b15c279ae3fda1a0dac07ed31fa978166298551c14742b9977a3879071c146eb9bed2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1837be07688fe2d70f8cb9a6561b4419bcb7a30727bc78e958ec66b89cb26148620faf6095619eedd05524ab331;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb46f03e805d098df74f33507db5f2703ce691e3a1f4126d4ae7dced25664de0a6fdae14571c26f2ff864fa8d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6708b282eb1ffd37a467ccdc3c5993e094f829744a7f07250f1479811cf56c2f079297dd157c5d029c97364e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76845eb9bb1b9c0e3b75a8376b2a06b745df6a676be7e0ec3242cd6e1c83d5338616e3e34af359e0ab325fb1c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c08d1b68d8d5f5717f2d79ed6de47b9e35b8efa8e85f0abec4aa2f1c54832e9597d92c4dfd6b7a193f98029c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e538d2324f43289a6917f92d425264cea025d5bcbdb1caab7d6bf2e5620c73daa4f6132e56dd40c90c823242c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92f2b97d35ae921d40cf2b37e9dd56538594e4890fef11cbc0c0fde116162a4b8ef8f8aba40129a198aac06658;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h721234d5efcb9080da7af78e7635bea612023a3352b94f47d176be8fc737bf5ab5a37d2471000dc6e8f0e81f30;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a4279280b17c854fe8a56d43cd4341f51600376eef2e9a63fe7039938e3a01cdeaacbbc3248c173d50bdea26c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a52f7f8d1791eb0130e28496520ff0ef9b8275ca2701ddf3255eac92b3e611af826ebe6cc8a331e78fa672dacf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d068c2ed271cbdb22a30e621efc75d0d87d535b3a47a30bc20bce3d8ea236dee616a8acc7aa7dce864d2f283ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164f8ecb03965bbd8bdb883d1d47d020de2e1fed3abe9fcb99a1d03d3d3c4eca000c240fbe807f9590e86fe77e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10500f1f884cdb580cb5fb3f82cb155686414f885d9e3e7528d690c52f09400bcb91ec7ae26f1f3343a9f547460;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd700b4c83b52060b08e08ae8d03cb18a90dd25f8c742e536dc2c79121148fa8c676e980c7867e1d5d5644d2739;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1385c4ccb08f8aa56ebfb590907f7cfeda1705d9aec9a706fe5e7a8f762642b681f34f73c5e78ff7d84f249d0d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103d49b3131c7734fe9af7e05d0f288ef69198299fee2a3efa12e11cd0b645233281a9c01bdba00d969ffeee62e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h527ee177a65a71eac8d3c743cd3fa2818bcf984b6577df734cf66f8b9b8bee3ca75fa074e90f1826326ead84a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h458acd0174185f5120c0af2e51171e220880c775953638f45277f76ae90ad14f0f248e875d71a2b2ccb6a8d615;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a45a71a17d13c08980b0bdf322601cc7677865ea38d80d67fe5415b02c401384745ab43af63c7de5a6c692a695;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116af85cbb742364cc2a5e4f77b5a6241b0ea03bc23862939e9cce940efe5219d09c5b5136ddbedef720601e8e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2fe5adbff19330ea6087730df78e5df492c4f9b3c946119ff64cb180a7f1cfcddc04683edf80065d25c1b3609;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cda64b521447a69562164fa2d0d40bebafbc66f5b40e530bd6f7a9941deeaa8e22f7306031fe8abcca7eaea575;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1646929972f5cc0a39092ff79138b8f23cfd7fd1bc3500504fa8b18a75ab28c8b7ff1a85639becb355a90814e24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30c74f7f862eb1fcf29f5399083e585881608280b5e2666a4c0cc6a6fed3dfff196c12fb2efb5e8722f194aad4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1207df4152d3f71b621c9bf96d6bdc859be049c986e9891ad12db0b0b170773a3848e4947ae26998ab02b2cf0b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8595a2b3cb3cf927edf373505dd333b1164a09ffd5e48611c00728f4f6f236959408eb0114150f76fdac1c6185;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c55ec52ec06bcaad8b3502c80afa24947a474b73ce0d290a65ad1570f88253d8663b4305f74a7848f516f68a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1efc6a921ffa29fb77e129052adf581886e05e7c4fd3a9d047445ecfeb9de01af885f85584a39b8b4491d7dddd9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdd96ed076538ff4630d6dcc5bfe46e3fcda94167f77a9795cd71fac1a6035a69320a0ac72a6d08144eb642f5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2069449a33960a18f8483997c0a3314020e81f14c91663daf51cbd0db1710d2f48083a50ab2a1daf2db5d731aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b82e510dde07e09cff59de51732e8a5e9bdf86b4b023b0cfbaac4180277ab9a05af1fa75954f6e2ff46f6cc1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146ab30516e2e73aaff5e34e34a74f5b1046249f4fe31c1b018c5736f67e42979d15791e63f2dd94b7121132a6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h793eeb5fb494b2112825d222c937645999dab8f783f8a805508d925a090793c7a24b3115121a9a82502c348849;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e30959a38f3182be871c611c63298a5a32222c7dbbd6a147e771c09f2bc412f08f87c669be8838115ac03dc2da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f3f3a3e493544debfa4957784ac528f3a3a01d1803e0c2a11de3321baeb6f7ce619c6bd22c236c13bfb3e0387;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183c2a659e474b286884e4f467578d84522a6a1e1abb49fb5fd6ba6117ed745608295072a0a399d6d52f865d1f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a34de65cb3f1c33feada8599d6ac513c2491dad8396e33b2daa857bb90cc51a05b5138a5b1bd89aef5b029ef5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc1928cf746f1f853e1c8c02ed282efd1f760b4cf50ffe45f93ee0fba001f6f927dd286d03b6cbf8098d758b21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14285cade42742066eea902fe034731eef2d7698c689b9bd45a12f6e343894c8cfeafb1d90d40e17acf36575302;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197c827b082d54ac103d844691a334fa5bd32d8f84f8bfeb673d5fbb07158e3a3c4274228f994f7e7846ee35069;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64b2f3cca66452d7bf78c0af3223e8cbd85e7b2167c596628c56e7a4164b0578e5e3f9e6c64a39745d6084f05e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53ac88f9b2a598b1f516a6f5e7a18b821384ad03e3ad310a6ccfa0d670e5a75d2eda7c52670bee3a87fcc376e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1816e7f49506d3cd4c5d5caf01f84c5106db9e053d8964dee4ae7018f0ffc440138b594e3a0e09adf89668eb501;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79d00070fb17025c78958459b34182856a614f08396dadbb6697acc99599fbee34dfd8e228115a1da99de3e9df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3d4bf2d386a762ebcf90aec159b005194cd883b44df156840efd6cc45582949703f8ef7a6a1a081082ae8f1be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1122c9429e8200b1d67d50531405b48c4565e05a045c82231c4b872338a1f1740588d257ca326bf2739a40e193a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77a7433aad62a05bf2d3898b11a89a1e20cf7c2a9f3bb0580e443c7c148b26188b6fac9a2cb24cc4e291e5e354;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c8237775a1c4ded05bb15a5af1ff83a5bd691dd902a4511e6f9a6f0d66bbd0d9232cc3e1d142e810e9062ed97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1918cbdc920cc65a650917ba57a596247b9183bb806cb7c8e57a9aa465b878810a661b4c09a3c330e806f49c245;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188799da9e54e75c61b5dcc5e48fbc7ebfde1ff63fc0b8ebe5dd18d488ef39a5ac958d590b24677cef72db68b5d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a1a026f6d8f19ec07a57ad1b8ac408320b9607c92d84c52c6c5537f15dee7725f90b42c142fbb7f404a0a2931;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90583711b8768d7cff7b118b083506bf407792ac448a6e1634925cfe2206db2bbe0db2743d460e5337ba4a0112;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a2cb89b58c864a29458c53c38c73ee0fdf47d1a224d1be5169e56930638705da4144f54be5669f55320c00cdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3311b309d1cf787b7e9cc30eabe55d2e0cd8497d726f8bdef7b0a46599d0143601b7234d2e73e5b6a0a06dc576;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef59eefb9cd04d8b62a6651d5225f339f826d3ce9ec1542958fd6201fa0b1ccf0ecbdedb1da67a5a448a23bee8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167481910ab6d43b770070f9e5a160075868a7314b3b042508cf929f9234c64dac54bc5d0cf927b412c0848be83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118bd1e532335b7ba8f15dbe4ce6cbd91a8cb74a8fa6a9482c01ff78f2ba6b15bd8daa71c3a54963fca277b3d62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fc274117709a7456fb52b02f84fee8979ba0fefa5978533fb7132f1d464adb4e08d3283392dfc6977eff7d8ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179ef14a567a23c8c9ff4658194f5b8c8f7938c703ede728e5d006bdd45c6375a7b0fff13ce45b0324ddd0f27c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdeddb3ea6df30e7a00fb65ada308f9ebf0c53d38abe8f6a234adf52b68dc3fc041418ef9bf6da43af12799bdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1313fe7f273178abe08c06de5e11f8aa2f2d73358053431c59c4df2f25aaa3e73d304511055510b0c1b9e2a6aac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6d3e9bdc460364eb44e01f0deeb7823f620d0aa078416bb66b4cb59b9270961794d914b838bdf077eeda4efa1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b23bf22e3c66223265085b6e9e494d113170838fd3116934d72f7c67d7ea3bd45fbd165e490e2e9f7aae461a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1494889520350ea3770c59f7b21cb330b5aa9d41144371a3bd3482c88d3646d95030a4ee410e99d03267aaef8ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1029fa04959ef68e05860154b05adb09a1b06ad9e9a670f0681c4b08f89770a2bfbf6bed63d465905c1e743c461;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104071ac8704a41a0a247973232133e5b7dc5a04bfed83fa50bfc8837eaff15edfa87ee9bb25d37dcd0933ae33a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1022e1f0d0976b5c3d20b3ef9cd529bafc5428b47701aa6a493bb8b36f8c4dc01ea02b193735c161fdf577dcebe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60486beea2182eb7ae5f64a31757456e7ed44798bfa7d0e6c4b51000afe805a8ce73ed3f53d354a18697ad6c55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d319d5e1a57c9f197caaa1888c879ba01fbc65d0e258de769160c4576a9b4613efb3c1a11a1b50c8284ee0aea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153f8acbc0816d9d5c034b1a30c1f1203ccb8b9a3edd37f73c1886d74b747eedd7a45bc1cfd3610abdc37ea151f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb24a4d65c4c2debdb4d3186aac8814a553cf7ae6653172b86fab08cf3ac6c4ee219903ed6debba2f416ad01239;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a349d7fb9aafbb571fbdc0462bd70577576c41d1f2496ce2594097d57eaca753ec714a5a2a9f2df57776107b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac069b997c6421e30177d831aa5bd9fc14c9abf979ee806af5824ba59528094fa6d2435dc4d8c37085cb2a1955;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee04b96860a34b1340ceb5ef14185e3eb08c1c6b2b19311bd973d64fa9168df4e70a475ffa9ab438da571e062a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180c8d7bc90d62c529c863ef39d6700b06ed390832ca6fbd0ae0280551538912831e3872937d146c8473721ec90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc91485ac7b85297ce1a9e64db8dd26a4164580efd02d4c89e0139b1c1f6f629a92d9871079fa069ca17649640;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14aa97808a47544040e52ad12eb642fda7569d1e3ed4f772b672d62ccb47e6a881d5c57071b4abfce48217baac4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a57ce4409d9020ae22173695c069adb2117228afb36b2a14e525492bf71096eec53a700c658880196fbb88c494;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c70bbe9e9a9e9c569d8e0d7ca7a91d31a35b81590654fe2e31bc1b605c75944d3acbacd71b4c2ce215c488ca6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdf40fea2da7d750afea0b49e9a460487f29083862181eae731c7c6da37782a408971be85c8854e7d3fc2bd41;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h847e45f7e372438308800b07a807e05e9534230bb0165bbfcaefddc563c2d12cbd7558b69357a1ae829279e45d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb65f9d01b6dc95715885cc6c5061789b0b041680e0c61207f47017b91ffa028f4486863308a4f5ad6afa656d83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1add673f29dcf858c187e35b98ee15d4996203cc4068b933324cb88d78e14c47a2ae45df078163240b56bfcb43f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca73165fb77d37214f6cef620e18c33c55c7a971c0a15978f6668467942e8bc2ee9bb409dc43e3b5ef09a3473c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb223709a9ab0fc3b78e1e1298f30f31d7b2c8bb90546b9dfcee40ce2056c50e22bf65c1b7b5e498f72311584b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc645f25315f3e45b2075a27aa438feefacc912c7d7b153cd3c0aba24942df2ebe6a79030e0e0fe1f229f15b88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5995d825ccc4f1703fbe915cfb2b00f6644b3b7a865771e187b5e5eb585dbb0f64b0d05ea40fcde0ade18e9691;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d060232b91be39ad88135e11ac4619400bb9d0c2d91d7e8b456b19b6ea053672fac9ffaa54271725bd3d2df72;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18cdbf91f6b1bd81a241c8e74b252a1e847155be125443083101f8f4025f3d33cbdd329d4d958136bc7e3bd29e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hedc3d64bfc043b8cbbf772392670e5b0f498933610f304fd644fcd1bc8f0629707fb2731d1a4655e462ba57cc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1fd251d6f38fe0007257b6461b47e5fb77caa83e9b75230006f92a27e966fa0f7712a7530b7d35937516ee981;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f436bcb3fd9577da75154914819c383461201ea1f17c09e764ac9ac2932d994ab769ea064b9ec60bf3f84a49e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c7860032ba0fc49e078a88aa8063ea4e46fcf3dd73528868fc7ad5a06d183ccbee0de5194be9ba1205108a0f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159ea82ea3bb4a7d2c3c4b92fde470a62ae96ca1dd3de2034ca16a4664f3493f147dbe699b5491c5f3f1bc7e4ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138dc072c4ae054f75a820d3aff0757d2369c603c27da3e52f9522eeab4225f2692bb36ebdfc54753e9f3d0ca6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h700b6dfb8490b834f98cd94fbd1af3ff417c7db51ea95dc72031054454f8b1c5c020f5db49ba6cc99d699f9671;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcff08089b8542f596ae61347a448a994e878b816e3b8308c9ae97e619a6021bba571ac04063caf1f22c78a3716;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eaf3ccf73464ea4dde8cd372acd958e2e187396c4bc13f8f6efa1a841cc5ef8ac8b7f74a16164f9c1fb5cf6f99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb3ac6deccde7734f36114355d2e8920d786bf91efa7129ac5e777e4cf4c81182d09a9a21fed032ccc951e5c9a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f9054c17458b58ee70125d1f4c89f62ac679cbd92dfae47408fa19cc70a3e8916703aa12b70ac769f66881e00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb71f00d8385491071b6c200fa983bf4bc983fc1c12acb0fde0c40e5114196c28765526f92844f7be0a5e82f0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106c50e9e5f25b132cd9666b1af42a41bbb7fe2c442faea327a2c22995c807bc21c8a032e590320f624e49cec3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba8f34d14e72dc924316ddbd6622a152d819cf10a2fb000a1992ae50e744f7f55b19afe1727194cc3133f6987c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c78ff4b50dd88703cacb68afd87a51b809f100f9eea95f5251aa7215a43cfcc2ead7d30ec3c9e71d45785106c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2b2187fb4d9436ce53b6557a6a401902037216348cf384d47f4a55e8d269d9cbd3174e08bbbf303262a5b973b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2e80e244101754ae5650dd66404ff748c86374ffb58054f3624a37e55bbab73af8f7ce21345dde2f96c6dcfb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30cfded98914c249918107ba1a30e6726e92b64c915e992fa187d76680909236964eb6d30b88b0bf06c0271a76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ce3de9ade44aab1a787278e1b9f756d06cfd4dc3dda7678f912f9f48d00cf25a6afd4ee8ba1885d08a2dc5271;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee265ec5abc896b1e46789e20206f48cad9e277bc9f27a9649903ee622b5f8747a94fb9ef08a4733009a2ca101;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98098129f6bbb1aa21072ca6c3ab2711f9d8192d7640ed96df9c2b121159280d488b1d96d816c25aadf04062f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1689b56abd38fef00f28ed942e2b326e990753575c35186cc491c357fda0c17706360864c2312c8e22bc0f0db00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4115a1432f0efa819edf2d3a86af09edd83568e7d9e2584ab28e3894786e715a0bb9e188532e40a58416946f1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47448f976316bb8803f518d97866d3330531b4237c6efd0927f91d16342fdb4b98c71db422752a11b3986fe107;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e11a1e73d027243c7a910587f82e21abed881848e67540ef0bac1c0626545faab593e84a528754037b6de72eb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h405fbcfe34efd65f30689d6dbca2b9be0099899c4772bcd561d10881756da9f2a30b12ac5d570e5e76da1049f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152e22b2bc4ce3be70d0ff5debcaf129c1bfcc623c627f3b10667f76c837f4572c7a37877b1264f52bb1be229a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1940ae7e89d48b07c77874cdb6b9903999cfc061789f5c7f951ff9a6d985e7173a2d3076e9b14f65a5dc4a4be92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1498f2c39d5c7e9d5d887d7cb262dfeed88bd716940e3d8192dd0388b6c0cdf596c4a9b4e53f9e9aebdb76de6c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h311d29eff86feb9141061dd665a7d6163f3b3ae969fce86765556eff5656225db69e0541097d093cfa86fb8739;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2e6ccf6c51227eef7625a7b680adbb8d8021ac1ad8b80d65e76db1d792f581c52b56260f48e77cd03ef524702;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf26c3cf848fb4bb8212f53c0007a6537baa4fa37df70de8532d9c95f54557bcf119b39f28d12eec2bbe9b708b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0dee1b272000a689614576ca08f6896fa2707f2724585b74113de6b0dc15197dce6b3c3735618243423e567ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62c93ab14600e8945b2f4243105cb7fa60d63cf29de0a10e641048d9e635cec56d287cec7b084c06b3d6572862;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h368566dd4419ab471ecff8153f26c866c7ec4729a6d2286ca17b655b52cbcf661fda661822c07c60cbd3776efc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38266002c58c7b684fe612093f06da8f4b49aebd90cba8b5e8fc91a7b2e7546e51f97b8ab7fa34fad61ff5a2f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ca43b49b589b42e0e0a1deb10e1f8c7607d3b6445d96cda1678af59ecefbe2241fd1aff8e3a8c9413e91eb597;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b0d3385ec1a6e92aa442bfdcaf6ea97f17a65114ac6513453de94cb518c2d3d8270cfdfb956002d81cb1e5352;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaf188dd79b6969fd0091964a0f50db9064216cd5d941ed267fde1cc860d470a725580a8c9f0f85a5c710d58fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfec35f69b5deccab0f6fea65d012e4e81150def6625a621e906aac9239f78aef93b93e484b2677a48e5212ccf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e01b7d3af0a3ab16fa2302b86b511e8dd86140bac0fa0ded38abce45035a3178f409642bbab55eb8ae76e429f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13674fcd9328471f674e0e55b6cd699f02ac0ad3b7568afa0fbdad2ec890ae9e8a3eb097472d5f2fff56c6e2fa1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdff882be78f7e95719a2540618a00ad2f1d97263c3bcfdc83aeead06d74c8d04e7f01e54dc37deb6ca1ad714b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a01a0c371807343738b6a830cb891d8ad5e3d474d0411c7d02086d9b6b24265f35ef99b0e8e3d107a95ed3df27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6e4f7791e718776bb30843ed300dfd29ec9a975f3d2d5b7d9550d235bbfd46866de58368e430f99f2ecf6567c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed6d0879977b6fa27a5aa04e2f0f2070d3364058725c59c6476d01dc8e3c1b42177c35ccba3b22014617e8064c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c3c7f5ddca135e947f72435a180ae3b0db01a61c03f8375b247f3f160974a2a1437f72336b347148e9e074d8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7da4f09596d86f042077dff55d6ce802438fc23eadf0d29224255c537b83397bc929ec6fa68b0f04d86e54b282;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed551b4a079db333532721f5967a86d0d1deaef4b1b238b68167e495f9ac333a50d7f84269da793f53a23dba39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h233c0bfc6404679b20094e57a86dd9411198688577c53185f1ab8c77e98655e91dccf56a9035e13f8ac0581ffa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b23670fb93a3396ede15866467b9d365cb2f27ac1f440ea0e415da0cae32c918700edf30b16f122709d361d20e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef7de0aea91bfee2c1c20b37369fad13ac83ee1f77ae6f99bd8c039c1eb00353527e8531b025c942dbd6170888;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1f7d45aa1efe835dbc58c7727720866b13ece747ab924d4e4a0ea3cf5d1679606858af187e9785786c0d0c07b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd07fe88bdfeab2b19c35695ca78d648b4bb71daaa973dba2beb4bebe25866b70428368b97c86803492ae778514;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4391de04fe2835f82fb386728a5f69f727c0ba58b1e237200082467b05a27ca96c70340b0de96642d14d40298;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5e29026264b16b2575e1e527192c9911ee4433c414dcb8085eeb481d2ab690c14f207fd0dbeaed50498fd5491;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1eda43c87d7e6dd180a2869f31f909f19f710075926e865d65982a6cd649707006e6bedaa0b84b6e5e649a5ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c437aba9dce7199c46449cd2b46471b83ae841213209a9925bc2e0df769d5c679d0c365269b61d6bdab2af870;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f90500efd95ceed3c7c851822b5729b2fd16029955001c9ae97239aa2e84d72a2bd82eb7a3e1e125febd57711;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1125985ab49806f01322f6b08d605b613632ddd1f5739e7717e6faff35cd17d72bd1374ba68205838caf21d24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c286861b5e4f46ab926a8b0ba045b25d3e89e1046863c1950ce43490a81711ba36e0a0eef5f766bcd136f852a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72623f9b012694495c5ecbeac7e6795c8d77ec1ca804d6c4f2a17a87900395273f1761e447227799a6afb1df7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173e752154ef88b80532c8d29b9b80d9b1eb953aff1568635af827b41df8f33931257f8e526455122a1c53bde9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14345200657e0f46aa8680b43d168fe279bbf75a3ddfe545859cb21d56fdf82a07a9e039ec8cc99c77b53ce2623;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65f3a2e69f6b10952c85291d3dc0753bdeeab3ad11c32052b9495ceba86a9c2ca8dc3b3792b7331e24a7f036c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5da5ca593ab9d1be9a14f7a03913b02d7664230466efffd9313dcaefe4d2da828bbd269e9072dc08d9695af03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd51b05143414c0be0837de45782de665f820ee34e89228e95d78d06a5cb25866d06c72282c510a19e86ffcf5cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de2e9daa41556714eb3f3291bff1ad6fca4c0e0a84555001d73f0b5f2a128cad4c2c190cdabd700a170bb871b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ecf65cee9b4c77889a6be519a222bf9a0c5c33e128c799d0ec04510439029027b116c3aeab57f319cea851b8c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1729a8574900b372d1f8715481722ea7d3312ff343dd1ec77e52b8c0be178ac8ae59a4c1babc55a5c1148962e0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5675d0b9527d658bebf79e088b5c9b1e216024b40888387d61c5ece32b0b8c859b0c3698af3ce4de6a25e6d66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1191f38c5c18b3a2ab666746365d5624e237a79e55108696e015a2cf37a2d61104c57ca55bf72e562c28bd0139b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29915dbe37dabf48cbf318cba2c18432b322e58cbc21ad88ebde3ffe8ba295bb0343b2505e936a29db5194cd8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31d9b052e18bdf929a2fdf52e55698a8cc2cfe26bc6488b3990004992603dd6fe330ab83a5edf57d0e74fddbbd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1108c89fbc97c18bf096ce49ba79d9a28d1e7822b2cf63f6fec4797bb7dc06170cbd9306c635cd3ec120e4b3ffd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5c551e1ada81a1aca133e6b1dda8e93b7a991d593d84e0edc7c06a942a04bc6a7c50218d4e1ef04325fdb53e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1697b65dd1e4a0ddb40ae1dbd81965d06c4bd2de1cdf89364d07b31f9d30b180d6a1831078effeb75ad9c983c0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c288a06dcb2f589791a016e648fb9f89ce2887f5d48da83f4ab88a74e8f671c4a90987fcc5925b8396ee2441c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6d2083d36ba4aa9680923e28bc9f519de7e0ba0151cf21036cea7b34ecaab7eb67e748082957162bfb1fc679c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db28bad87ceb88907368e5c11005b6d2c2b5d376a21cb5fd2b14a83364f22ced33493bdb454f692f852acbc9be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1dab1a175a7ae599780a6f4ead5ea09dbeae835f40eef3b74cbc27ee3c7aa4e7400505f158b59fb56322efd41;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h523786b67445672cdae716c90e050c442713b42bab1eb7bf857c34fb896c7bb2c4627d5e0f97d634c09dd5f7be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a775a9fba6ad044670f65359dcd166075d3a3af182e3410e58df0674ec6f6caf3c9fb19aaa56dc77abfc0e1a7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b57aa95b455560c17d3ec97ef398dfb979677d253cc5c26caa2eaa5c19b2314c9c700c9c118688966fa46cae1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haac3272bbde09cff901615e93f865a526f5ede1f4fe155e41bc49aba7abe018a97f3c93514658568aa982422b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a904b6181a812f85a81e67474c08acdcd9546cf5c4ef024261c849f84cbbf5b61c540399b3f82e3cabcbc1e248;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c63ae0f6731aa1ceeb64962a56100df4128973b8d933a51ec5dfcb616679971cf5489af33f3703cd256232af1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h735b4dba549d7f5627b40c092416f3310dc8f7bd56a73b60d29c6b25d7a202fc4f1e09bcd2f827f06b188e82ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71a33920597466472e626a4bbc16ba227cbe5766befadca04648566f814963fc96963d110186f9962bf0a976d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h731534cfb067e33527fc7eb620a1c2d1d3f5b1a356e570f012c1ec4a520403f700e320bd52d36c323740afd38c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3943e38cb86e7ddfb9df801eee780fe864b60a19e47bc7267efd84707574377607fe33dedddae24ea982b201bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15092d7c06bac2856f462f13bc3b95a3febd02edbb96fdc715274c9065732705af006b85b2f5e065381734ca95e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13dd56f81c13aa2ee10e39be220f985da7694beb06b78c88d2136e0634248f2abddabe4d8db79a90a7829cf18f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ccf1087d1e2a8aaf41e4a479d66578c63880ee5acf90e696d7c1418364aa732da156ecee50b9c860f0a6570b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6349cc244256a1660150f9265e0bad4268ff010f2b36a2f70f2891389b0ec548f1b0c4c497dde008ccf76b252e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18637bc0f2246f403d32424a1abf83af5c5afe678014eb5d24339931083ecf85ec21653e166023c627c3d7a07f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5b73f6cbb73df47934c895bc30082fd3c426de89baa340c459d31285c89e75b8bd337c6563d047b0d611a4582;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7c42baf2a70d5e5cef4b5f0848d4f4265167b2f418924ea7277ed58616195471fedf23ff6f721eb1c28d29321;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182bea2c85ab9fcaefd6a04494e2b31c1f510783b3b1f2a14982e5f93a1d0d9668306db97fb3e99f4a524b79bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb39f44c2a715527d0497c1334a2d262783e1d9fb2764692c3116dd20aaaebb32922c1c46877cbe90341f10080;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c4e04a68dd4d3435235a7345ff6e7039f96118d36e6bc3ff5ad80be78cf75c0085f9719b91e645b0681e53720;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdaf7ae16b61995c06d9d2da948d22501b0ae60a36f6db0d61ad00a665d003f73290fca0275005f0a90bddd772;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb85be9328d3994a8f2150f4f100e5784103840e46e4db421d14dc5ee417a37201dc4c0e290684489180a24abb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdaa20f089dc681d690e03b1a6895e57a27633c0aced468ce3c11b37e66dc3d8c030b1a5737010dc78d1af988c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24de0d9ef544ae4735a04a8871c2bc34199619e0d7d5b13619199194106392da6a4306c58b54db100ed33c938;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1194fe71a43aeeca70c7b869b8479d23e307b1d986911636f32525a330350bd9d34a19324b2b32d5918c57220ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6977d98ea14cf23c8d96beadac6d8cdb962cbc5acc3bc6210156dca8f84ad4b250e626b71ef2801c7e85fa10f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78c29254fffeba924b53a0073d56a66f27399bb84facba6d042c6c76399a0be41d4044a8df175a3804f1c29de6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee5b91ae964c7f54bb264e1c0d4f38c8782ad4f08ce45b44160d9f7392a1183bf0a509d2d388c1c6d26379040a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab8bc516f34f9331f5f8afca57b8c5f4502b41ee5f9514f734bbc27649d4e68740341be2cc7d70318b138c7c49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a50513c6d22f71e5f7598bb8a5cca8b515c19f0390009cf066a9f6475a31778fb9cc799b098a75db93349e0c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed82d4da3f29512d37f129bbf7c79da44d37cf06877126a5bbf749b4417a0f00a07bdbf62c32d2d8bee6b46f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae227456a3b784b3b4d6291179377f06831d15712e1b17a78c4c334c03b7829e444cd42cb38dc808a8e6a3ee38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15096ff1da99ff768580639c5a1147a9510d4fa3d049cfda7474f0201ff031c156377980c888ba601fd995fb0e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160c8df6f01d6f7c71b254d092199c1222bb3246d1069f2b54874804a8b1793574ea35d4deb7572665c0243a405;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84700a37abaa5ee5d5ebb1001181cf9f2e6f876ad90bdb71b212a0a5150a3b68bff6206b2fa2e633a1142ad254;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf07ad901e34ab300dd7246079aeea22ff117ce693ece0ae3ac2e0d14946c5ed1f23f0065c622e62e3e6b80513f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b2c5af6536d8d46dd4ff10e07ce3d2a41bbb95f67fe7b47c40b25b58d65278c899bebc77119983f871260dad2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154633be9be169ebc9beb176aaf1c92d9a43bab70a9cedef10c854a22deb18e08aef87614a195aa8877f159ff7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h463e5e64a010480a106dba5347bc04e2e0ecbd1135423acc7e82ac5385bd2bf86a8b07f9790b19b16765d9134e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdce3e417f3a389209a8dca69568b54e164a83e7f7d3a192e0209959a83948c011aa7c36f4139da4b0e058b725;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15809402a3f7c27991b65e9c3beeefbd6bc7e18341b3e7837298ca7a29bac7d89475f22f71a62f25bbc8bbe1489;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9c329841f098cd5c2db01b72540b71c6ee6d3ec0bf075501896af439a421806d021175d8b3eb3ff1cf1d42c68;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1089511934286d368aa379ee1e8b52319541a39d0188a28ebd8e327f4f4d8ebc0c981fcb5fd71234e6dca677f05;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd176687ec7085e1778afb7dac024570d8123cc5456a7a8fd5cc8cc16c5ccfed16500ef4a3bb214b697f44d076e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9ed317540d5e0373eeb01871528d4bc8c9669728bb986b472d4fc0558ebc8088c57a931c629ce197a33eb84f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130513478b26760eb3116627d877d8f6f70a6e1117f1f5ed6a91da80a7236f0fbd32c9f8e8227fb90ab749fd8b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ceb52a30ba9a7f1a2f2a6ff71d5712205237c245e8d249b9d3a1fc4628a96db6142a29cf2f98e3e0feda81b297;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179cad1723fff4fe9bccd30baca15ee3641f802e7672c2a02e87d5b65c6ce248c6cddef3788388d39970c466e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcb717c2f2cbf9394298cd28c13444cef21766cf94cfa525d055d7b717a133ac3108a29e55e70295d231569054;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5c6145b8b1da390da91ee7cec90c063c3804376869500e57941bf08433b00e9da5552b40d41c663e1c10aa2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c48b5bd1d87b3026b43ce556aa8f71c0e08fbf65338f5ea602a32504e73c25234e17467579f2e678484d017441;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1e6f71ba40e3e7bbf558e64892f858c8b2896439ca00db433568a649428f603056f4e8d1e9a5c5c808264fd7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130e486704616372e3c4082b86d52efae377b1a53d028cbfceff18fae08730d4760d349246828b6458da40acf21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11830797a61980adf1a54321ec03ca9252eb754582bb2fee1f283567a4e0d30885f6cf91fc623557f9b9ffb5a53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db7f6c07d00875f854661b2b9a5fb29d85b2a928cf88b5f90c03fc751944f0e9e04c88fadbd0881e33222865bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb843e0c42835aef393023f998490d6eccb58c6fb0d241cef794949a8e8d64e60ecb5cfd10bb85a01895f1be0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ec3c7ce2bc3682f650b3daa80fa30e6406215625655ae13f655f4cb8f4e08fb9769e34b1a288fbd372fe696aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5625cf12fa3b9fb866e860879ae7bebcef38c9e9ed31ca9fd58448d31090a5e3a867580ef01a4d51884577940;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39e8b1bdd14182d15ea644a7e03c31216c6b995c55a1964980d2e93984c85ce6959b6e1d127a0d6737080dc6a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70da5df95a2bdad61c29d3f7735d7deaffe7f3c89abdacf85dd0a71b61cc9d5f304a2819f22c2700f115413111;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44c84428287b81df2fb5d7e20a66a6611f9302afa3253f0310a909998f0ea0e15589dd7dad3cc87905220788c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fe741afe2bd0721cc5fedee1e5cdb0b1a6e81de3a8cf1c97b21da68004591d0b4f375750f4b06865ee733e1d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdea799c06f955fd8543b50b9341882937722886b93dc578816a98a9ea76bfef89d651a9ad73e6f2ed3946ca8c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d57000445353e1bb8dd616903934da80718c78d9ec7aca3c69c2897a458751d5798f196622924a9a92921f66d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd35db523ac2b047865499c8e6220a147cf0103b79f9f1e9c4a9858810cdae59a527b8a500b4d2da618ff4697d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5bc00c0fffcd23dda1208ab5cc4457c8d4d5784ffedd05e8122b5935d21c55d91e7d88093731032c91d884e51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fddbf2ffc08e0edf27fa496ef7fb4e6c8b1eeee3330b4f48ae4a71ffa205de65e810d4d3a86153fb19203dfb91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haff1c8f8be83d6382aefed7bcb89c2296fae05d9b7163a32d1e050f2d794f5c0cb76a96e9350718f9f15959335;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c73c06faf86d2b7fe03cd7dbdc88d13db8a0fc0396320bea3b3f87c0a3274be2e5212ff7a3a47009b2ba206a69;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7bcf8fc7874954ae9734a472688ef17d260b865dac4aa2dbbc16e82badd532664e5056f6b2f95d390c8217b1e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54a097d4fc1cdf04589e246d4c88724ab83606abf0709a57ae119f1258264f99c5a30413f39680dc62edb5a79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dc0cbdc4e68803f5984cc0d941828201b32a113ede7b2312371c665e03835a6c7433b4e1b19524df328a36844;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d8bd46995a4fcbd3d105d7ea6b9343143f8c45c91c77b5a906e2bb0f37639bba13c252cebdfa99b8bab955d7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c1b86aee2c2dd6b3341f173423d89d86f84ad99d6b3915ae0f91492b2de0cd49a1ef29d574d90cb60765cc440;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9f78a84fe0591507e2b7145569a50e5a6caa9df6d236c9f429d4a4f8f9e44025d7876f8f609f1ea796fe62aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bb7691846f4c5846e33ccbc5f4438a7ffe7ed9c22304a022fcb0392f9f4fb40da156696923715e0b963a764f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1349979d436e8e7d053f7e898dec65b0813a90f14a77373e9d941af355102e7b4f2f1d55d11dcf8dde596edef72;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0b9db609aeeb142301934fb824639badfcd44f5d8e87df466c4887644e3d0772468df8cb80b2f9d9266df48ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de0a3370896f720ad5a4ed9fa82b6969829fd923ea5d4c0d5af01db98476f8118bfbdc29e0001e32f065cd5bdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a6c313dc456284e12c3d36dc74607092f0602100f4abe0fda5c3f00704f81fa9120941892fabbb11e6c9a367a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120e95e45fd1f6a687890777d204050aa4d573ce63bdc7b9d98ad5abffa781bcdbc00f8c13eefc1b766e6809ece;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b31b72c55b4ca9df3132b105b0f6e607f053a5ce80930fc305603609721b3808304c6d874d0873f676cb1fd2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11869be323d77db6e44f7194aeb026bfcfa12c19c6f8712a5036589e096b1b79034a27e4af075ef4c464f3d598d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b16622ed50f815c283afa132c50e0bed89d9cb31ca15019892b0688cd49c442e50db4230f22318c518196c134b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f73be8d1aed246279899ee24fb27c9504218ab54679c3bce0cd052cdfa256241f9dc0c726c682e01ae4acbf0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16154ee720ea8ae5eeea737047d2eacda1e5615b73ef831227d1234bba9aa0fb743c8eaeae6641f6fd4b0043d88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed93518566ab48f4b33ec36c594bdf979046e38e0e75ec20f8e42b09c23a122c50a64e7c837158fe10f1fe1ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd5adbad7a9a7d56b1aa57a11ced201185dedf751d30d169e659548cac7b6a5524d9cc346972a02a434c5ff973;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75ae26173bb3697c922f6a30595bd90ede7122ea7fc2a78ac0520fdcf4caabf37c9dfb39e44a61a16ff4c53ce2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182364a390470a0788e2f4dfde9d24a2b79929ac721c53c45cada4c99d01f23d01cc3fb51620c1a276b983e3041;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f95097cf8f2c852a658f51c376be0cbb45b5fb2a588063d4694dd0c84134c34f156c23a1a6603573dc495771d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9040d3464e015e4422742cb45fe8207bbbfd7c24e70bab9809c5a133e840c5051b3fafc99a361449367c65e17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20edd245cbfd71d9548daa8ca3b64c910cb6e544a477504968688d965b5cc74f0d6e175365a6092a80125686c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ad29bb554bb64cba19c4c50fed880904dd30663411c92e70f67b215e78f8d261e3de6e173b8d9b4483c2c801d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd108f762da053ad6973f4b67c96c7ecdb6e43d42d3c438e10ca88bea292aa1c452d6087215a34dcdfc48700c09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12feefb87e5f5b23d716775735030e0a93f5254f93f91215b22081d28844ddabd096f56ab40676483ed7b088d6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3971d9c614ed5019ff142176a9321f58f4a8636c5ebc684e217ad8e7287e2ecd319f69cbbb4e6cb51d55328ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193847fc8876ccaef8be5746faf3d1077ac11bd5d495ee18268f87c3c7b96de27b2fb62d904f95cc145bbfa3374;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf47db600691fd202709a78b4b5cbcf995f9b1405db5222759f71be579340a6c5569eac566194270682f6b9d9ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aaa3efbc997ef13bb68b49d30e0ce5b82baaae60a97815a3270d68f83a8576a1121fb61851853732df4cedb3f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c9b2006134c8d069097aef19f842a10bf93689139d2f7b501e67b6235d2ca6bfc8402bc91ee8e0653deb65555;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bb52decdee8eb304452abeb29be98a9396336fbdddf2b4aa0f481d39ebad73c3f357a95e76dac063ea96d9112;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191e67761cbf829bc70c8c9f0cb7ca1c2b99199f19b8659d531c62fd35c7e5b459bb260034b716993ae21b9e419;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h190f4d74fbebc76b03434b8a6d16cbc02629a6eb70a09502a6db01503103e21e6965de8cb3bc8ecb9c0b767b601;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6cd26b3cdabeccc7a689ea3d6fb68796e2c96842544c7db531bcd982c0a7dc67962987f2ef0815f992fee785c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d47d30c4adcffcc2afb59345bd00d8607b3ed79a57722aa36750029367875b89541b2e56a7a5e5f7a7768e832c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h594e453761239fdb5817977bcb5024036e188b99997faa163deac34704de2635c5a2066d954e6cd02868bc4e37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1152fcf2079923f8fbb79a66fd90d8eecdfb0d2953c79086c62212ae3517e685330de1f94972eb708cdc0015fb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd2c3100226c7320b061599b7246136b51da06a0afa82cb7774bf82b6c299d869a4b4b412c52d5e44faceee59;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he53b5e1a5887550a01e832cdad2bf878ba0ff87125ee4a143ad3704f427196a455a71b530be9416a1049fed5a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed6ffdd3024b77f02a768d93653c36ddd0e9b0b60c5523b613919bb7020e939fe09242da581a825d4af488dab2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0063cad81d44fb7a501f3364ca0296b546d1a2e41276e56fef55d9adee77c5b8b9499a16ed157def3a166c303;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d37ecadf63343d223deb82fde771be23fcc88d1a5a6b2a6985504fe86799844703c9a487f41c8084bc127b3f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4f4f60ccc71a7a7e488502c3bcd533cde583983af6ab92a9db2cb5639f6ce4d8af817cc320f99fd8054be26aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160457b492d1cc7f79b3cac0e06e0564270ca20f46a1f40d0cda2b9193afb64b1d689e45a48ed69500de02dbde2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55ff5abc858d73312f8158dad5c7c2f01b9e31afec568becf18ff3be664c70e9790da8a989e8b188e111ca0cfa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1488f451e34f58f9e97251fc26f2d9e36f246f1debf6c9b8a022d551e4d0238a016d5a333c27fba79b1385cd159;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1ab4bd60cffabf83d816274a8d44bcc8506dee91c2a1da12db6619c3ce8c01afc4ae5d02467d026284bd8eaf3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3318f0ac9528f9a5a7578f231355c9c07d839f6b1db47cd90875efaf6a1d1fbdaa3138c68fd23198d730dedc59;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc3d41c0871801b7314229246500db669cd6e2c40e36d6c595228e5b18c2ee353c0b451107fe93934c42e253fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb55289efe29450d832b201f8e01c8510c5ce132e083aa610f26d367d7745089ddd0eaf38656cbf0ec2f2cb92f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9178dec14a93ec722af7c06d40cf42780b19c005786d9808a82fe23e83b4b344ac23af0302f24880f4250b74d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbfdfadd914ac00f0621a0a42e215e9f6b1b108de82072fe2d10991943a6ed44ce7b1ede37ea44615a1fa4d344;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb461c1b2ed053bcdf89dd35fcdffb5a865e269a317499d229d785af8db1986cdceb7ee64840c1032ddc548f806;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df2ab14bcbf4acaadfb2b5cd33b16274aa6e12c41e462cbc253784680859c9e1f33f5bcd156b2d976e59a481e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9549f9ba63005d1de189a97195d1722288baf450ac8a3ad43618246ffcf919c2a92792a6a9c7d84f293bb95eb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fdd64ec626f130256f0b591e7bf8a59509e9eebc0998191da24bd06d2ee68ac0cbf328ea5e68bf4c9b5eac45e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dd6b45fae6e4f251a852f0ad11a728fef6878627090e5830d70bce7e6b24be0b1f86c4ecf2a381d8880f3e125;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e85293e85ba743a34118148760f03bc52656fd98e940aa97232f090a28d429c28acc472322b545f1a634cbe55b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107e2a8941188a0526792bed1b852a2d326ac70e6913c94a1a636a0934b7bf6be0e6df356711964ffc9f486a8db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16877a05d5955a2e6cab422c9bdcb80c32702497b6d4eb1044e3ced4074a30ea8f621f8b84738ab024eac505534;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h278ceef9379901ef5dd005a6d8d52cee6b0e8bf303dc8567f6b9cf578583dd04e3bee469267a6d8b5f5d9f3b67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd8af24494cf765867d3aaac175fb00475233de1b7e890eb0c3527e6c23f4d6e60c5a990e763746a05c299c11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a9141c8c5f1fcc78d938053a629c3da74e2be83d0f264c667937ae27a31234a04c1a8e81561156903401034f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4aa8b561fee3ff858199a2e2f96cd45f2adcb3860065aa8ece18e0ce6846285827471d5bf945fcbdee838ffc38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10381d0e8923f940795f11d57b944d36a9038f0061ed16d71dc1b87a70a76115b04577264f0225db52625761fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23bcb984be1b960dbfd093feb389c4e262bb850dfefa11ee744b5e50a615f3347ecbac32384c11f0acc54b9047;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ac3e6837a78c5403fc7fa8c20a3c0d267be6036efa149893c94a56ae06e5c44a0c11f7a7356232cf84af00ed1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h759b3f6cd6f14b5a2bd1bd23fdcf98c72d435fdee478cadf101757435fb8c1e3824066179fb27d48fe2e77aa1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87f9b2749a793359a55a2b48475422919f111c85e80f74b9bcbbe7860a651abba2684b3d76b8ff40e97ef6e9f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193b5e163240914096abb8fa1d4d0bc351fad9479b1a53841fdba028de88d7729d873ff9752a8065c63777d96e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec0112f9ca477862b3b76aaa472b1a9ca9374c811fb8c4c33d12b4ad6635d9890fed5387f7ef570c1e9e658f79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcdf29a3b1d945bae65010acaa63074b105a459fb5b57c057197cd5e218a91abca2086391e8f214e7c105400cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb89b8bf8cb9afc0b90c15d9844217e92ebf110e07d16dd4d996251a749d2e9713c8db65722df87fe9a7863764;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb235fdca319eaa903263f7d8e2fcded134854cf9f7a68e38a10ae02004da5ee9507fb3385a97fc3a4debcb7eff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38704cb7ef4fc333862439c14353c519f3cd6e8315d964b9b89f91127c117325e173b0bdefe0198dffa8e7d055;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8119e16f994a3e6e60e16c9f2acc11c82df3a0a9fe9046790985b816c1473c7a79c44ab229b5998e39f688aa78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7363168bcdf5c9e5ed7e3b02bf41826de31ab34087281564ae2beddb94bb19e457b6911166296bc8550da107d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28e4d478635fdfaa62f26c11ad8435626423dda19fb7dd690125d820b452461a1643c0ba3958772ec98426678d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d66d703bc4e365e6e820e8a1af1d6fdffe8205244dd2ea4bc9d4d1c5b93b348c2b8a51afe990b300847134c2b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0cfa7f26f296e7580a7981a903b10b3db61bb1f843a04694282973642883e8eaf081537362e51bd849c0b1895;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c5d01623ca68d419c816831e3703e80959fee8601671da0c961cc3976592c6195dbd22c0979d8ebd921cffb6e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b55e4f870582f8c1abdb75e08189ad61b3585b73937bc92c31ec48862280be79e4c7a59d5c992f10ca5030678;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4908d8a827c3f89865dfd6ebaee589bcb70d3c4e2f6cf4a3d47d0f502c693faa6ac1eae995fa439d7662680bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51c7cd0613619a6a8ffa8869448f8051df76dd8a20ca111f23f82cde6df65615c8eb057f16c667ff400c8ed201;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25176993d1bb6603fb9b6bce33c4e0c6d9e7117bc913664861417ed1de2e174edbee180d907068f90c66cf5a23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h503701d9a1f546de7f9aba12092db2ad7bccf9daf2c6bc789ddc5dd18e49ae40ff27e66ee1b1f5761d390443fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h623afc852999c7995b6b3a2e42cf49d6f302d1810e364b2bfdf83dfd83bacc6e2563ac2ee08705952695e60759;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc6bb8353aa97165466db53267e0c93a0baf6a5268eb1f37710848d36712bcb3e6471e83056bbf3abcdb99b65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4beb1df209602e2b5cf8f9b0ee7e60c7583f449ef75e71745b7171b0adc250a5f9c07ca400ee03f1e2efcfc45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b4eb31d8e415eb26b8eb8c8e225f1906e47ecbfab104135f1d81d6d62e39deb3935425502390d736bf26d3f50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c8917cae01173d0a447c63c1c46e2a1a9b79672f4bcab364e3b12451f8895da4b411f91a6c7db2a939109ccff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7947f65e7113924ed58fe0273ac8cd0152b76798d7101cad1c7ceca23e81676fff1aa96e9c9165c4b3b8f9f00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74d970ecb7d713ddfdfd2927597a7998f8139361498befb10b8ff14e9517cbba41db3385353a5fd196255b8b3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5684f47bffee20f3cdd843dd370c33cd42c8351fb3e3fff974e83aa5b845470be39a4cceccfeec636833c99552;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5e8305fe64f1ae9c20e007bd744978b5b22607df3ea3179dc7ce6191457fb41972eba1d9828e65d7fd0e24cd3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8900156e4dbd273ee8bfa84874f7cbb02997026fcdd04b5dd55cabbff5885d60b8e08556964b342f3e352bb9e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8bb86db678eb3f1604618d8d9ee5293b76b663fbde0c956ee8ccab2646802d59ec731c11e9c1eadb2e352ce3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef027efefbef6519c701e643145e525f70f8eca5ad7e36dcc45af2d01d7d8be94bad244553c4429de9e353f090;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2ef7783efd65c35440d4653f759e3f6b3755eddecdb8e745b29cc37782e258b2a733b4fb8f80d43b95368d16e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58d17a3c7e21efbc703fe3fb15e51edd3ac5d943777aad0bdab0c7e4bae91089566322d257559e43ed726badcc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167d0aa4c7822229c76bbe7fef135afd24622c12d1bda176d238d7dcb554f388131b33ae292d320f534c8a8c6d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a4cfa8247410fe91cfbfe1d5d4d727e98224e735d0c9aeb1908128c63cce64270867fd6521b3a1521d0e030e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h272fbf82e83027554cedba3f30be5c782de339d37829903211376d2de9b78da1916f1fb6e5d0367201d669f5ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ee7824c25a4cad410ab16e1019400d459c8103fcf7e1f272ad9f2601760a3e72456cf86aeb8467f8d55ea94f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156eda414c4bdb7526e9d053329d8b375a0b175e6b02cffb57e8a8f311e284f47aa6ca0c25f5257e92713605244;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77c0f10590afcf1228b73cefe05bcffe4b869af7efcd39f3e12a1d50328cef731a162800111634f2d41d2fb842;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dd768b47cc04c292516c825808192c6c3f47000ebf6db17d9c97c360ff577fe1c25f39eb912e0d9379d30dcdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a91b8014fc617218a06bc12c6a3e440f9c1a603790dd6cfd35cd1c6dfb5658e43cf0c6d145c03c7dba3aa1f841;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h972f58388788df3a67933cbf96ce373830df66dbaf919a68695b0dcb80a6cda59003ed86db96d933e46e161a1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db6fc1d0908dd2212ff4bb258f15488ce71fdf0843f6b791594c3e5ac1e848b41a4319839ed819fad93d586509;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h615778499db7be9c12ae6469ff450291a2277891fbaa18b50d708352380fab2dfb69d2048e00630db6d683852f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4d5e08c21703c06252e4717bf49a5d65960375d05eb675f9a76a06e272c16a5f83a091df0bbbd05f8a820883d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1513b066493c937ada16a2317a924e848e75e66a2794bea1b2c7a6d0d73428a896aff54360c147cdb7d6a0a3d20;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124d92d8d78018048be58e21010bc19117a29d0a35a99939fec5a6043a18e0d6f4c37d745f2b9273e417838bd10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e23e41c6da1abd74530e0713fdbcaaf77db2bb7e75a2f075d85580909dd55f4179fd4e195c153f3497a8a6ce85;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a459c260f7db09408a6b1a2d8a81bae399ce9f0f2e7cfed298a81a2f039da05988eedb53afd0594b90c3f7d8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20464cce90ef070186764fcb132f8972ce01817c25b12d568b1625cf1c44f4ebe539fecf2b29c17fb4e2d554bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e2560aba7ffcb90dfdc2bb7cb9d5d7261da99d84955d641e26d06b846b4f32cde9f20b1161a6d0073951ed0db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72e30b8f9a336f7d2a1a0749c9971270f02dd0ecaa3d5ab10156df05b8f76a6c0e36d4d7d88cdfa4e39ab53713;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f39ef17efe6c8b2f5c0f65dec8d91198c2d26f6a28731be575ec4580799929d4240c258354374fbb36439efd6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1789d737f58a5c0e184ae0c9e67329e175744b3ff9cdc83bc3f22847a44524cfd39e8b60260f914231992b8e075;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2a14f1a89d80d4061e109f6092743713f353688f6e94b2ce9d0453edfb9346743685f64c8bd1580e082823d24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2d5c879e64aae24829c68972ba45944eed4cd3280c68d76b61c3f3ec67cb7069508e56907621c55d62ba79f80;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0a4e5796bbb73fdcfa300e842c2b0d053753cfe542f6deede5ff84e8f9f9409f55c18f0d73027789bbd798416;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h436f1581460f0dfac6a33125cb266658f4bfe3b35660c04fcd3c3e20a7ae445b978a01b386b6fa80ec1c32bfa0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6baa79d7aa2d109e769fa446a3d8727cf5fd3d9fcd88e015d25da8b540c06a66ad97c4dd89ce9bdf9034a7a430;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3755b42e78095dc9e30f2aca5d09e24d7ba23568c0493171259aa2c060d8957e22b1d178624b1cbcb85b3ea1d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f6188fe9122c57f652c35825c01114a60e5ddc4bda1e6871714f54b9b05ce12c0db97bc804c94c4146419e2f3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168e9a3911885183ec5fb8087d4ca0d147598fc050fc03db31b20734c4b8ef4c0565999a629630967145fe4f13e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140c43e38c3a049612db176655a639e00ab413a5019415582f02a43f68e4b4937947fec7efe02dbf8c726a59b34;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9edd96e2d8ddd776dfbb2638dceb3eb8b830c95d8ba7686e8997cadcfcbf5e8ad77fe9c44c6b83983fcf8c5bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c49fbeb14ee9ef50aaf921c9ee525e838d117586414ee0a170c9bc47974d6cbe3c3af669b0c39293cecfba68a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3029e82b248356687db02d18add5510b7d0e4743c631b854681f3890bfd8f76139d7181d150dc80dd06fe4552;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc363670baf94799b4ac565e936e3b2856c65cbc83fc367f0fcc48800023982bf6acb0a42002338435f781fc75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7e91095ea14060531f84b064d114cf82ad1cecac5063fe4587c3e9e8023fa92ac360fedfa807ef156e34e3e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c5c8cb7b907dbd70689fd9ff73e6f5780f68407d413e8039e0d79ee7d457f9b8a6a6e847512e9bc31a2d19367;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197e0e386725e2eb1b746fce6628040a3bb5bc293f174fbbd053365dc2847ac3aa9ae418c291605da84d1ce4e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7335317fb0ac74dd5ea3885502c0a25a5747d2e2b62761952bd232f43133fdff865f8d862f212fe872b4ef22e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfed990cee7a85174995440031037dc9b063a24ca8ce393f0c433c02a1adffb66e2c61389b3d1c4636248714888;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16844cd8b925ef108e972fc520b7206308bcbb74df0ca55ac087c56ebb373be4706d415b030bde7adf125bd4f1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c6e6c16779211e9b21d640f8218230be9b4b335a0b8932fa30613e7518c727d1ce578589782ddbb9c85d089ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4fcd1e4229f075c215f5002a4642f132a6ab366bb98d6a9ad1cf886243d6bf034348d5407731bcce7b30d6723;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4eb543737c4ea9ee2d11ec5183e097bf67765259db96242c35f2aa87c4376a9c73e2e602c020f1a9de08fcfd15;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125523a3886fb2b8b816a9bc307e18f5c6916a601d2fe34234951b8269fe3d6555f06273def7ccc456acfe8938d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9227835603073ca47baf9becc50e84d0f52329b3b7fb515b28d5d74452354b9b761da240cc1778d5d13ec04d98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3539993a340b0c3640b6b79844457fd089fac63241fa515b350f282de4014e4dea06363cdf2e448100c440d673;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181d2f92f957d4cf08f25b5dba1df5540a381c93cc54f47d91cc101cf21f8741c85784647cbae1804e520b8e872;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b4a64dbbddeb3dd7756c0da0cc28fd8a7a0cf253714d56147baa7a1a484cb6c9eddda7e64b5d8c3564abec0c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff4f4b90a69ab49467646b61389f7a065c2853aa05a07fdb1fe35be8ffae75ee78bf187d9a8e2cc5a0ad71735a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164ac67a0c0ec55b11cdab4777f9e89233aef5e9e5adfeb3db79c91cbf308f82a9fd32c6631393c9a9b4f7621f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142f4e3b15599f5a32e82084d67d542736579b829962cd4ff5bdce3ee41417ab2ebd59d1e2b80f79ee15f59bb35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99dd8cc8301ee471457120c1b59a3ce1d67530f92d0fbb4420005f5a4ed6430128ea32b911ab5b2104ecfbecfd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db35120ddfaa4e7ea53a1b3e0fd72fe40408acca4cea6b9469f4c481c5751b13e033e2b129d8f67373d02003d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1fbcc5a31b3836908827e189d05cc4d5ac58a38d7aecbefcd42ab9fac6dd5ac355885bdca8c3f38c1d3a42530;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb71cd68317cdc581c7c9927505f5037b4f53ebfed8294a9460a93c4aff672336f93af5e057ecbd115bdebfd5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha29c212e5ed23629bb3eb7629a8d4f4d55c7f1a4c149bb4748256e39521ffe6fc3afa5846da1020a28ae9875fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14adfbbebc703669a292caae8135e3c7b344ed9e2488df5a574bc41f501e3a0f2c23fe3b7a5e1061e85113046e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdd1fba113ee8c9be43b0f206c2cb7c5d7a02174ea8d8dcef6223d7c7695c844b1a1a881f21b95aee29d360c71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57028471cacc7e9d3655e7686533d54491ee91acfacca707df7e7c2cd812d1cd62a3170131c1de2dfc28b3d2e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7d68281e920a3d7ad97cd0d718c1b9ff793967ed5e5b611ad254c7ed93daf48a9a5c810eba83244fe18cf2a73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h113c0bd6b878c3afecde8760dd6eccc0630b783ba878bcd3c87d18816e04d634d46f80630c1dfb90514ca302dc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1336aade0d6650382c3b974a887f39eb1fa19735a477fbc89cc83633e33c6573e84e4bce6a0cdddda16b3e8af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15bd95a771c91c8d846fdaf1d08e9082a12d0c770b8fb84853b9b96b1a9f936d1d332b65985f4824449a4e94afb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111753a859289a6d1b1194d8c38774f4693ccb6e019bb7fe21d91f87e1d770eafdf5e8265da3f516cbe7ef3d261;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4440213b8ef662d2fd7a1a34bcc5a11e26f1ec2cd4be8ab6d169d99630fcc25f4f1797a76cdebda1edd755e70;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h631d57ac7c133747dd15b90dffdd3879a8450bd0723ade016f92bd4d235c6f9911b316cd0995870c11b9f4f3b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b998c6d0af21a62835592cf3836309232e4343504b151f6e71d459d35992f07ae5af0367ea4a5757cef57a29c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf70b373acda5385ed15700d75e1438175efc0a6242a59fd4e8de7c3541e38ebd1c6d992772d006cf28a2dc5e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f9d9f68a7ebfb9fc830aa92bc7d94513733a83b7a01831d43925ba82231c0d46cb92e91036327424187cb004e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d97d4de060768e686e558af284d7567c2b0a3af59e22f6fe5c5a1e36cfabf789d7f9c25a4aacc8baec2a2e1b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19121aa0e782c32509dab5ca623b505d6f35958ff93b1ae14eb1e56f435e900651b479828e6a7cd0973b4a68266;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10725834c54424a18f692e3c01168d9be0f116dd4c27042153f5517bd5dc9e1516af4d1e68c5e7dd941d28f6068;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dcbf44173a84435d58940553416a8a2737e905409aacb725ac4a10dc8b91957971edbdd7ee9996d9185eef26;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fa1a14426430b3fe87c763d0fb65164a0c93130f3c9f22cf43a49ccf56e75219f43952c7d3e4229b11a3d90fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0d47da028937ea9360bc1c8eec16b92fc18a71c83ca9b985cb9ac02fa918ac5ea4b006b19ee38f23c6706f976;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c6c33672ea1c23a86c05d2a639c869a5f64bf74e7c614311c98cede2b569571af9aca72445de783357a517186;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he845ac3b60c69bed07d220a2bd478c4ed0c92507ff703cee21b99bf3aeee11987e065fd69dd8516bd1712c6637;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4199b81f1e8135eed430ca5c4fd60d1866ee66039fde73d94f8f2cecaf8d9923efead65a8044da65cabc46963;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1a7a3f312e69c007e374cf25b272e8000c9d934d8e9e5915bfcc929636e2baf02e3e1cf8de950b8f84a35f2db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbb9c435d8bf1af5887b012722052e56f408a8f8fc4f5bbfba5d0dc1bdb88090b57609cd6dc268d1b2b6c71364;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18501be33292a2596108165e915b7c908561292c43c0cb57208c947e4b71ffbb92e670211674e619a102256fe91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc01f3204070f24073a24c45d1df6a1adddc87e12b0b2ad59bde92edd34e67f9975d65d3425a60f48ffdc29ebed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1324ee5a43b877f56858bcff95d3f08c7ef8d160fbbe32497ad48a060b5626d1b114bf19c7f9a2c31e57990ba2f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee6b586f594916e7c95e4553e726dbbf24f580a3cfa72deb4fa1fde5c469958f628dae8520456126c3a4a2b2d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122c3aa7a384f03a8fcf986d68d5d59e95efe7f73880a6e6eb6e3f8a5bfd91674112a1d2cebeb86d68eaf6a092;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e037d918c6ae34d2ff8211a5b3fb12e758e5a0cd6e171c9957c6cb5d88342ea70fa6c55791e6a1ecca7f4f77f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aab12507bb9370b0f3c33e47f140b165cdae0d9afebf3e04050736cfc4c427c38477e92538574f1f7efc81fe48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha492c09be7742b0a86e67fd60d1fe37eaac1f73243ccb6a8621b0bb020a3f03f046989d9577e38f32facd16c63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20c2e2ed4c33de1cfc8168f73ee5e75a93c7c8b71c4dc37d3f631e9f9dfe6b27d262e0d0d55ae1fa20d42dbcf2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17edc2165b0e61933d2f3a0c9aeb14cb08887413d8c50a9263049306f43c91638a79b263c7dfb6e3d4a0798082e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h881418180cf837a1aff559294ecf8536bb0696797c2363a79d9e3ee844865a06d21031b6f377405a28758e24cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ffb4f9421a7d31e6a5f0c4cbc09017fa58ce027e4ce2e08625d3bca87567c685661831fe022cc1d2c2124dc27;
        #1
        $finish();
    end
endmodule
