module testbench();
    reg [19:0] src0;
    reg [19:0] src1;
    reg [19:0] src2;
    reg [19:0] src3;
    reg [19:0] src4;
    reg [19:0] src5;
    reg [19:0] src6;
    reg [19:0] src7;
    reg [19:0] src8;
    reg [19:0] src9;
    reg [19:0] src10;
    reg [19:0] src11;
    reg [19:0] src12;
    reg [19:0] src13;
    reg [19:0] src14;
    reg [19:0] src15;
    reg [19:0] src16;
    reg [19:0] src17;
    reg [19:0] src18;
    reg [19:0] src19;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5096f3fc94986ae0383affdab903b3a721abe51b2eb26e4a19f68e9bd80c9cd66949f67589cb55abe17c47147d99542d9947;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha36818954c0fe35d4737fe90b3eea05fb8b3f165156b1d1d399337bd8039c712a19c4bbe8b3e6423da49a9daf4fcb32ababf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had1e16812fdbe822fda76ce8c0980cd4cc328df44f6fca1618ef9d63d6d254de38a69c7ef419cfb8c8e3c679f85a989f6a7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4933916214642960d4ca9ff244545f5eaa9522b1bdf7600e01c403061f3046abb08a72b2c2dfae9fef075f1cf63478e50a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4ed4ebee9798fcae27714de9451415fabe50f4f76e3beba648b72c993cb4131b3934cd3ea0da6c502b7c52eac3cd295aaee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7307c9ce579d3f755a5011c979cc8f51a3d1752efd935039d5be69e1e91a19088392e06cbdc4469b75240ab661c25c28a0e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72ce2d30508f3c7503b04b1af4b2ca410ecb23ffd4af4d997efd059e457334347f6876e9085d71db53c0a4acab94b6d3900;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcb1219f0d4644b9598874bc86c81819b9e041b022c76393f7b7ac104db5f4f545ba957bbe92f7b62550bf242fec05054ec6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7053fd80711abf768c1118af5a9cfa61080d18cead2e33e74c38731c2981993f9c1e96663307b90fc90b54ce3cbca9dc7c9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbccfce29532a1ad394dc6cc90590e8f79f6b06a53ae042c6b3a09821dcfa393f63dd1c37e544e62a2eba74bef203d83035f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc55f96f876f15066756295e77fc9e146ef18bb2cdaef3cd435940dca8fc3bff014d7c2b3fa4ae610bddfb6c53e4d33103c75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf717a5c0452db2478e530b9a8594ce82691bb11adb3b1ee2939cb1ab1654001c52517dc573ce7a4d630ea41a65bbcc9c7224;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65a8e86958cb274e6d8fe7c2d5ce05096e819a6b38ee2f4aef1e68466ef60251f64b75ad88db1982e6b64c64fc0d97d3026c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c79258319d68eb2f4d0c1c61ed5a171060ae3dd3b236db048c58d863bf1d409bacb752b14157865a6179e242fe14801d60f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b5be937e64c2b2be4d04a9d0c92552fd5f12bda260003cac58fb729497daa336ce0d5b94df48898c3e3dc2d59aa72db7c85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb83a790da5f5ecfd90f057b5cf4cb86a9a5b080e509fe00eb24a8fbecd365473e0146bd44b380d41144966b72be697bb54ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f8192ece31c33333e98fda7e124d8393faf597fd8ebf05dbca992d550d6bd7c468e163aa11fa6aed10f5e125c5f3232318b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc5d5530cccc0ecc4abdaf3bfcabebba160bc7f098cb9ae75be18138a2de57066a5494975b9fa74c15cc7a351ae84271dcab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc2c4944e3d6d96b754b99f78df47237a39b81a0c64a60bb9de1b2ddf392e8cc557ca980ac1213528eb45829e1ad02c925e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h337a950eb7d1b71ec2853028128d373c3f26a30aa4d0a3c2addaa41839d91e1bb36338c42e3652f7f23ad262a7a9a06c8ae4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0f8c768d15e9a14d1392a24c6dc90b582480133ecc6696154bc781b28367ba37714edea5f6b3b2a582369873ddb19f2a60e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64429b2b46b9d98e2af055c1827412896f5de0359546afecd65157a3a4ba0b05ec16300485fe7fe6307d49aec1693dbbb3fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c4db2c43a02d14060df5e4bd8ce8806fd5526d9af24b8ef4c7159ff2746035ee3aac0caee65d69ac11de32108d2ad15e699;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27953b78d1f6aea89e22c7b7745b824622172035594d157378ff7d024fc10fde2fca24a550dde3e6fcd109522165fc773425;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacba75e3422c5df7850a632ed647bc2720c14e2651db636ca06b4014a116b1cecedf1bac473562de9d21286b7d37543790d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6626d5dea472ac89792baf800c0de0ff5074f681e90a57371e512aa6ba33bf45325239cb15f6d1c55d93bf154f2e37b9977a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bf64accfdce01a5f0f5e968f44b87d144eebe6299aae9c0c83f24f3aa8db0f916831ad3e2901b21dcc16225d0c3a7cb0246;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h287e612b21f58849d382f11a78cf99a7d771378384d738f4af07db7ef397f046a9d189a6b2c06e7506d75c6f801835e3efa5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56a675df9fac1d8ceff32d5d296dda4b6f90de8aadcaef26a7bf0107239af80ee48c2cfa0b9a3fcad0bf97e7cd87d4bb9546;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5728861d95dac6a70484effcb710a0810b63149ef9ea297ea3fa10bbe53440997c839eda08685017ef05a462b3af5becd626;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf9db0ef57e204cd3fcc123171645a9683f495595ace86594cc32c58df9ae162e589da528a05c3da0ea93e9c68d8a4db77c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h558a6a708f0b1950caa26f641df9dd5cc42b2d2fa74fcacb273af273f32960381decb8c2b17a6a6c977ede6fdc7bfeeccce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8bf4e421cb56d52b6e513d9beef35042a9ff8e30408de24e646089344b15c60eed4078282da321f18264e2cb25de636642;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f33e38a11b42c52cab59743096357acfcd34d2e0d70641ca45f9ef400f67966e0496c5af0727c8124f663f368f53bb1124f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h897e8070dcb9af96dae9b8503168b18881a1c7a2bfc74d649c26ecd87056f9eb8bba412c45f38d68ea01ff36074cda36383f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cc5e2c29a876dbddf91dd9e4857d1b86b1f1e4e6c1bc2396f31d08bef055abab8004e7f73aa36adff8c83f2cc888f2baf7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4376f5399b070eeb4eb121c3c23c18ee05e4cc472ac4fbeeb15995bd1488fccdc61b6e4545c6c1a01388c342f0d36e31c070;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8af7d4aa5d776ab3bb17b3841380e3ac93b2cee39fcee9c170bc1a01203aad0b31103e34e3d5ca199b9899a097bb5b97b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b0065ea93b1187d8deb87b03a8fff406e8193042dcf516623854b5981e7d0f6f4bca211e44250acf46a0db47174a70fef46;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb2a3084e260d3aa934bdb02cc16b304e2e1abf5b0d2fa7cc071f54a683c92da8fda9b39ea493217722c57aa40f936cb1cd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcede84f1dd70f4006f2c84c6c6c2417f96def146d33a0f03f47f5ad50567a71936b5c2a756a6f9bbf5c07f2140882c65906b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61d26696b6f5b8aa9a115b2a0378c5e76e912dc7bca2288211b4cf1bf99a8d78dbcf9935964f90749853e4f0a028af704efa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19772a633bdb7bcb0b2f03912a110d5a285d1a794bf1af97b813208f75b1541b1d7f0894ffd7ed45ab8f5311cf9a3b761c7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbeaf350453028afedb63b8c5ca29c0e1870921742fee3c78f7821d59e9b16849d36508d94a149212b83e11993de1b25b31e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h205a098e2d26e48bedc44f1a65af03db83100d282f2d621baa1dd59c03efa212128d65ea019a7b59be333ef1b8bb3e890772;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76fe4a3cae9f13f04389a49044091a84ce0c3a7e0e5a35133ea4d23a5b5af153d2cc9eb0fab9dc84d336875cef4cdeb80f97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa35ec4b91098a95a13468d5882d58d02e831c148656966dcc03a8e0e70afef282e9db06a1832bbfb6f56920d44168c1405a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24bb2a5e693195becc6860261bee3525c4237f4daef53b02136e95963b2340ed3cbc252e1a5d547ad6986930e70b7d456048;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5846d9ecbfd0ee8a04d85a7bd657155f8573618ef0fbf53465ef4fed24ba438bd07c4bc45db4d4e2c61eed0e33dd3a7244c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6210ac12cd99da6e9d13ddf1abb3c46207655b5dafc5edb3aa716854a8bfc661e2b8180ba8618bdaaf9245aeef3f6bda053d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f9c16180f0a9cb5027937f24d6c030694d8f5a656011d2e265651a93d11c1256a05404adde84e0f5e739b2a8023be03f534;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d16f576e415fe84979dbefe57dd13799ebe93dce48bfd85956792af36d15a794502f1c0fd8c39b2298be119cfada3913a71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he92b7ce411012a800bf6c47e576a0a0d293e15de0d42a3f56f9b74251767052307c2e24ed7b55493485b8616160587c9e9d4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e87af08a739c78811390fd0c96940b59b2a6ff9c9d8f8462de4e1e72674fbc4e9cd72a381503016ee4ab1e607175d7d9a01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ee03a895c25a366c3acd69b8a8e5d6b88cda34dfb810f33f8d01c6a276b11a2d6744dccf9627ffa272700ed33851605fba1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a3b6f7a3c7b9b70fb1c5e11f303c1aa22f0b59322074a00c02ba779d3e0a47c201874aaee7345008067c562f06a0f390a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3b64713246a65b224716d3d77e25e0da902f098f888f61643183551252571c9d8b0ff01d3af052ee8c31b56dc236aea8e8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bafaf246c685e9f260dfc7208f528763e77d391a706f71c2727b519c9ac514d38a400686d0779554c961c3a0ca175f42934;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d7c75948eba8ead23c09e9aae8bcf099669c4af0477f4ee0e43cb91bb187826baadd5718bd4e6022a985cdbe8f2247e8d74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5afd4a2c00e62513c8a9d883a825bc29722010da8ca083383a06c93a8e0143f8b6a5abf84f66debd14b347614b6e93e27558;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2c90ef4845fec7eb451a97a1deabd5a27c1f605066eadbbda8273935ccb674bc376b4a5be5dfe2847aa390c16f2cb4f11dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63537dd92f71e0ae1281414717e9edbe44abbb22ef4a56153fd378f10de952bf5967d2dca0f84e2296b7e8ca0d8c0eb89149;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb765c1c1de1efd2e589a3dd95ba17a93697c9f9034478dc79aed3988e81dd24ac59d03e7fe9635378f139dcbe1f808d1a731;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b62dcfb8834f270a9a9dbf4d47b9ed257d7affa470572ad347813f211a7a47e168862360f8dd26a7e12c5820d2ba19e1cea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73b2bb9d68e4684f438e345bbb59c211757331e4ceed1007628fd05354b5949322e67cf93fdc2b4fa94ffd5d88bf1696254a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdac8a60e8fde11c03fbd8b135974c0408603e716f047612b3f0dd24ef260b328a8a527923b3d16ed5ecfb314deb24b33085f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heec6ce1361e9da4b1466ad6c57cd2afb16b9fdf88931a94f0d07418367bc6b3aa006644ddbc07f776fba3460b5256d8ca268;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had664cc2384819927daff9b394efd8748a9440d633ae600e69a3674033497439abb6d7074da2dd6066f4d458df1a03f83c28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h286b0ad2e172b8f46cdf3cb1ac85960222e1c0eda3d86709daa8a73b9377a5fa4deb3fd913b853758141530a36f7bfdf6fad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf9c227bc222638ca1bfe615e6a323913232631b21cdabc8065747d14d83474ab8062cff3dc423a59b9626f34d7eaeb539dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58c2347772db87309876e79780dab27c2cc69d25ca2794abfedae96f6d841f9eadef7f437a9d7566b6dd4435819920a42ba4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd4397acc6d1deb1c06115b3d3265d323ad5e3ae9737a2013c7c19f3cb97c783ef5198e75acc85cf330839cccd7e05f9d39a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf82628ea317c27098c240651ba60c08cde6b6f0eb1ccdce26e7e78ac7b461a6d55b97f0372972c7dacf1dc0b4ea2e5303d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf81ff606358d8456b361c06eb1d1f8213ec08a563b8b3c9050aa4ba552520295694af3e58ef3aea2fd257a680a765304956d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h372c1bc5bfde45484c515beef650092be14556f82cde4ce4c5beab7afbbc1013b5f74765abf74804ed3795bb7ac8a3606f69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6649f07acc11385d518608c5379020b5f3822222d61ce8ce5e865cc32804a66c5d7b986d24adaeae8526822650a9ec015898;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haec94f105ac2f56cd8852446d8377dd69eb5c58fcbc104d6c692849f22c4de7ce01768575501c6e4a5f8f80e97a2ede14d99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8a24fb2152d360d930d0d12063d762a69a54bc011c85a5a176043dd3ba9197188ff983b24f63541b4e95cbad7fe7108e680;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3c73fdba915c2841ff3466fd02ba2c3fca2b167509c7f4b21802d48a13e02a7719e2d1e2407b23ffe1ca7902632f384b5db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h433c0494354930fb540ff323acd10ed8b29bc594c6600693e9895a8547a64d59ad93078bb6e7785ea96a7244ea2bd30ab46c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f4cb8ccdb439215f7e854fedc4430d49d0606ee02915140e752c765ac3aa6902be0de02d4f0ed1525205e47fff0588cb776;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8cd5a6026b9990ee60212fcd7d1c3cc500bcbbfaa3294f6af9c1274091754ded54283ad31b0558fa27fc17465420fc48784;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8229a037aca757b244f249a2c031e10cb096c92b32d4db29ad8a631f8c967862524c96f973820ee37de1ead2a93c29a92fbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf346df5cf09959b334092e30e8864f4dce1733f63c7478d0bad707294de608718b98cee3d1e0cd5332652aab4c892681fbb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1164567816a71005fc425b1105c8acc144a02731205e998e37e558e7fcd2de890f447c1f52ff83464e7911bd313b34f45763;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf694dddd69f26def6daae6178ab5628d093a30e31c640001a32bb53a71f6e8ae51d0cad62f3d0e0b02c01233ce593888eee1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0df8a4bdafa5159e432a10954471e57c55c0079ea9951f8854232059d436f9462d9ba37cb9b1b96d2e4c23d98c6b2e4162c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a221518ed600025bb8e77a7c34ced0acafb8833848fdb4a428f52a3cb0d3897f5bf2a36f99538fc1438dcea06a6198c44eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e923f956301699e3b929cf6db563fe23751461b2e96f00526939e4d7db10df26dba52d9de9cae71f15920aa4db65fc3d71f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb131fe360f88f78fd94d0938cefa601b62e5b275c12628adfbc80748f3c44a1c042ab3dba5e0b527e71ec729f5227c602698;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d17248509812ef5d8ec19f4779b3a50200ea57bba27e8aa354077c1ce90ea4d74df21de923dc46fa9f546cca146efac8dd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9819b92873d11f678381917527e33399c00df754e87a6c35e18d3b61ad52ac39c2fd9f9450d373a66641183e3a14119da70d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h192d9660f7c8b65c39814ffb306041595380f93a0611aa992b6d15785d4dd738587073c1902b6c55f5332c242677c38691da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h223f364aeef29a965b7cd787d4633108ac68af8c643d1b713665f99a3acd72945d5eb3c95ee6e6a03ee2b5d294f742d2137f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf82a750792a141c0394dc38d082b8b132903d0fce4166161ddb9650d10ef7d929635c77a75743b3023075d978326390cf0f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6048e3a4a0d9ff392a8ec0a80908ca12900b9c6a78b528c184b1e7a8c706453569d747849dadd560094b91c7e0894fc4165;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he653f5b7da78de3c4ed0b92dd2ac3ece4226d93b30be43456e3c5d65d861758fe2993b0a042ee022636ba565552df6a6333f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he98011f7dd9fd20750f9091deb487d34f59daf039eb1fbe25acb0a0b3a0d87388c66df41fba09052cb09f6784268fe85b9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e323dcfdab82443274258a7176b4fdf26c5c32fc53073daee7ed7241ba43fe4da84094a62c577e105db84f1bc8d1b432d38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h608777c8ef5c8ded71a07d9483b6332aa0356f9964fb2ca190365f6251460d21c1edaf70c4313ec1947fdd437be6bab07037;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8eb41062d2755951bb2612ab7ac6d2c7baaa9a156929f185c3387f6496b0e6b80a6c60f316eb82b324cb46222f170914a06b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha88fa8dee2c541e1410989e3e0dccded8862d61e5e085afcddc7d476e33db788ee3401c9295d0d17a964d1d8d2387843bc52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4cfe493286977c4e13d186659e422986ac099386bec55dad46ba2e8ec3e2eae7e22bc5c546139e1da6144333dda9aa0f88f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h848945fe0baaae9c8addac11d3fee464713b665d17f91304327fe1d98e21674070691faa59b4048dde363f4ff65a252c0da0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf4edb16f976d3171fb1da201a2fa6a857c9e97b3588d8763068829acef5c29e4c66a22b74649a86fccf24f44e5c7e953873;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h392aec16fe0ad65b00371203b3de7d12f029c83b0636078c4a863dffbb778d67407765af863259e8fe9928309634879a99b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd893511ac26fe1ba893c28cf8906c8cb6f650cee2b426541874aa1da9eafe02a636a6e1481516c224fe0f3c05fe77e83df29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27ee1f6e9a4e8c0c56b6e7aa9e822d6f5ec13049761e3c2a57d55bb78dc190b25059a98aee170f99fbc07e056fed3009a6c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h788ffbdc2a28e6198bb7afa7c7e7bfc6bc7f66e825f92e89e34f1a3bcff3695a55dde5d22cb3642d5f4900edb75734739ff3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3cc0fe52cd49b824cdfb3d3ceb1df17f0fababe12443aad4daf9dddb417b8c433813a699c31f2db9a27122abf804444b304;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5089319b518c4781dd92b54d4d2957a4fd1498e9d0bc20bfba43af020b4c5691288350f7b94ed03606256ec4b13c6e23da4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h982208f8f504891afe2c0e2f9fb7b12f28f7c7318608f2fe72b767bfd2812bf6740b5cc241342ebf5113d2d15f83aeba1eb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd68a6de789bac0c21e3f7f9065f9cfced14e4d7bc291b3ce54964878a4f03861f711376e8f0259faf0a52ca30bcaf94c2db8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h261299aacd632ebcb757fbaaf6a23f009018ecefd86c0fee4cdaa24daadc0a5bd97b39139f212d3d0f5cffb268037bf35a36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ae16b7f1b6a3599ab83a08d80ec46df392ca58f6506ccbd5b49e177dd31c069b4abc48bd86076edc38856cc87fdee13a455;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51510935712bdf1c914b32c955b9578ce3e779e097c469b77471c36863845cb9ce59cce3f063e7e12e319755ca1658e28ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10c37573ae3940477894f1af16d49e0fccbdb0fdf6fd7f4366fdbba9cd650a751d2fa72a184618b90069408e7256a94c4ba3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he887912132561f3386e07250ccb529af69c83dc67991bcfa046c7a70ae290a30542437a6df118e2ca61c1431182d30c4c89c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb83176b7811246458cc6f5669d7f6186892a42fbb16dead11d53f5a0291abb71d0e1cdd5dd7dede48802046ea5b1d35ad9ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h873a9934a84a5d1d0368b685c17687b7e246eb0f017cab68cc69efe7b12dc88116085b9a82816ab5ff998ec2c36ae2149e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fd4107d113e0b41276fddb7c4a1d4798a524f19f60a74c80d1f2be277813202b15d3667936d1cb1515aa51948ec51a3bc77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h837482386f8f0b160d575a1918f642c8f788972fd4c03c5f831849caeb745a0a0a919abbd68f841c270f13833fd3863027bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7948e0898a48b1cf6d09177a4873d96525e9ca4597d79e3b5a7123ddf7a6ca7fa16dd0b88427e80f21c95c20eaf22e523d12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h504d7920dd960476b869afbaaf090132e0f67ffdcad13f4a1386042c2e04347b56deb9e1e3cfc3e1267aedf0b3aa4c03a321;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f45df5c96fbfc464de511ca24d8ea4b7befb9f4fffac05dcaeb52cf4c92d93cb2a063c216e16d721aa1c8e0471650d9ab8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4709f59041e02ad00bb95d1f3a2a82256bdf923c7b6b0a339e57845c58fd91cadef266785fc35c62e180b0bafecd62232931;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha562199753cc5e755abfb394812f1ffb2a3225de60344a3769d1a971249aa7fa9f46b4b58b8a482cab512b1f89e08994fd5c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae3f96fc53f8dde846dc74500ee1142808972c958cc84144597c2a8196a1ae09d4197530ca93a82926ba73f0e503bac080f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h233c1cd0310865fe5bc98471735c075138f446cbfa3831e25eb9945f6082eeab58ab29ff9868cbd1c666d50910d11eeea05a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb1d87ff3cfed4df965e7ab2ddd6282dea6c48d36ad6f9a20153c195f341d1150ca9e91defc165e584634461777d1875ac4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb638c894e1190a1e603da6027f458f5ed56761df32cc72a4364c046746aa276ca8bcc7e4f283f0d59981e71603072f8899e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aafc6902c73bdbe7270612f2dd17f04fd601573d5b6b3ef550b4a318e768715ed46b70b1adf4dac92897abf32535f69910d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf97549d174289700f174ca3c09ea0f65913a22749a8f47ae28553a613a178f0607cb8d85438b76c0a7589c467426e18b04e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e5ac4b152e457809b31bb953801126c25313e9014ee452b93863f68d4adc383ce4b05127d90ffcbfed890ffde98210b15b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d0ba9ae0329e4267b47711e779462a5d6640df36e27b1c4a8097f271407e90b7952777d57ea184c5cdd5f751f6c2f391858;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he026d9c3dcd8b0c1155b36b0c4ee9866e73bda8d133e39860ebed3e4e99f590230563714ede84db8d24d6e0aca9713552e46;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h426cdafcbb8c4ec7048febc28e9d60fd4a922e3af9adaa7d8e3ce1434a01b3ef285ff5967e8408a90474a6b7ef44892a10fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf04e3abefc2e9f1374b87249ed94f4befa3d01b79de3b7cec9301c95cf2306715a9e36ba13d98e7e3509ccdb91c81b8f4aa8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3e5206410d12cbd9f48b2ae93fd0b34cc3bb9ac8d23b7ef889ced264c4ff724a1583ebe944c910bf874812ea87e29b36054;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8ba4780d76c0591ba675d7114cd3e3a03faa03c9325fbea5ff61d8639d2b53aeab0b90703515fbc1404c0babac7fcf3051e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a4443ca8bbddce64b89997fae9b84eb02ab8bec0488d3031ab48a3511eb1353eb07ba9982d3af4638a9781287acb9013f5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc591d1fc8397910e1582abfe7bbf289257c82cdaba5575967709517254dd5d9bcba5bbc65ec5a6f985f1f8e876d0b15647b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a54213d07981d580790de2c41ea8dc82886006ee91108eac1b557242daefa3e72e570b9a23dabae3db49affa93166154c07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39581ba36cca3f4fe3f20a8c9900c3f8022d9d3ac0a80f36fbf3ac8bc4606b2e1c6cdde8423717844b4a952afeb5f9ec0ab0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59fe1e635fe964c7eb2aa61f3091aaa8d741359faabb510c90d7fff8edca20f17fdfe8c5cd06aae5ec67af50187cc1a55f4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b50898abc6519cd9f04e8a0a25efedf625ff7cb3ffd28cd4a42b0c16a22620887403a42488016d095fb577801b214933e37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc26cea51b430dea5f22bc102721b03b55d00917d6b22ee327f6470396458b486b1cea9c11bb25f17759cbfee45189dbda650;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a846cdf8572e8ef63760f734e36e910add12561c80230024e9488a32b850d0addbb8e7229143607d7707c7159288e77b64f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50a11a8f4699b6b7de1247f7e09e892a1d5812f6bd5cb489f38b0b130091dca8dd77eb8473bb2a69a679ed05f737ab626b40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha96012d64ec1d2459a6f3dd95f74833e11f5092ebf6a28a7ce83f5c74069d7f75807fd4c1d7b37f4127bf218171bbdcff802;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ce77969573e77df6d7fd37ed6cd4b39f6416f995a9a4f7ae48ddf93a474e1430bb9ef17c7fa5f1d4ec11390b712d381fbf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82d89505be47eac647b17c50b970847766302bf4af92ade6dee9d12a126e03c70cf4391a7120b1eb345f280e0ae1d5f3bd2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18c1f9f778c30d2cd935725db684216af202a71c7a9654b6c24723c902221c37b4d62970ef3f475cbafbb67f5d928bff1ff1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bfc2f4e432670c6b38b982c1e8ce3da4c509fc007e00b45c323e34f0a90965e82bc2e67e1a723fdd1e3206fd5394e1c0878;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h470fc64d595d3113dc6e16b1ed89cde0292d40d93cd7d5a24876cb5d0da10f59b5dfda12b44a87704f41d10e554a12a39a28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75ab61daa1dce3dde54a589ec71a9803bea8d1847250d9e7e9908a44b29d6030542941752f02cca661b96e4610ee1be036ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h505373743caeb17b0a97546a39786bf138b904099a020952e06d845a68d2ddc8ff3b7ae7d3365faf47ab774c172b314798bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha52476632e9868195beb02a9f7590fb50e13f367b3ec4e4732e048da6fadd188db05daf3a909c3fccd8bae5e4d6a38a907c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h837eef49b3fcfef9bc21343ddd27203222b35ed16e6d9d8157116f62eac61c47e6143fc5edb0e7525fc8a39a59192dd4c740;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb39ad59bf376fab804ce0389ce3a38043dbb9583f92f8be676008b6a562ddcced024c6b26c17e95c794f84cfc37732250b40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb67c14c2bbb2745f8f3813fd2c2bc185bfbd2f028cbb96a5b0a1aeb9275befb9b2577cd1be7ec910702033c50352282c9136;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1918115148d16dcf88b87da4fe92db0c8f3448f758e5097bc832417c2e2a5d650dff556dcfe21d44a4927bcffe7a9c04ee96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf49d067375eb2dd7da83874427faae97f0a468e194e504e39d9828fdba32585b2ce28deb79f08d1de209f5977ab08fb1aef4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f0c3d3a3aa5f5da964ee46067366728075e022481c07cba26a3e3149799eda9ad191e939e6a3e129802b654eaa50f9d3072;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4e03436ef089a182f92bff2cd6e87f16f2ee3dfc0f40b2d4179015a61df1e9d596c1801822eab34d7f208289d15ad7f76db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3edd1a68f97418fea0b570e9b5875e07c3334d1e1a029d7b137321b753be0579ca34ef83d93c7db43c118c12c24bdfa6b7a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f308df9ae564cf781c511abe1dc8652593829ce2ae992ae7776b2a995e1be0e045cdc9dd0bfbbb52913e4b710a237ddf991;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e86f564706ce53a581a2c70d7fc31f6ca3199756cab86b5f4b2937c5cdeedf5fc86c010a7402986e89f2b20c5376028d5a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa77e47d05e836547b891bfb427f13ab8a26dc2baae8e2018189d6275b9df5a4f02c8fb754e31f0bf3bacb7b567eb4925a8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb03a0c602d20aaa99a2eecc19fd67a7046722318498d9a9126b19f0f4859df506df6bdffb5422ab9b284a5f6aaca81f34c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7db7eff92522587aac0a907a16f463105a4a42db9c73683d7a88c6eccfbef14e5490a5edd0dd05c6d41203a78583814044;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefbd424806bc817375603c7674edcb258c4f4b14995865d67cbb49bcd3091d3e27763f94f19b3eddde6e7a3dfb53922f4e1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dbea4207804f071477141e96d470ce0b4e26fabeb0e8105041d386512110399e17ad678d8eaeac574bd5090e301e8811cc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2c491a830b093e5b5072f3d6268fb942c752809692cbe550c78805cd1c53eac6951c81eb28c5e678a3c67a5df9eac04f8b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef701078a4a80ce304b987f8db5039aa6c2ee89a6fef4af4644e78f928799d2e08b25a3dcfbcf5a9d03e96d94b39354461a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d4b3451504318cab98760b9e0f92b7dee4486a27c96d76fbe2eddc9e5e86652cf05d895b5f128639031b149a41f9837fb50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h994d900a4c3221b2b1c6a6738f56621df53d8e97e5ffc2b5c35fde54865cec5393e4f4ec55fd6b0202fa1b1a465e908c00a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45393b3f832ac73a008cee46ef4ad8711615b6d590f03e85fd6cae1748dcbccab11d99aec3cadd550286d552ac345a522f1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd15b961092051f064660b8092505d6c2614cf1919049d15853bb6c09d646611591f92fcf7475bfabb3a6658c3db91a2949aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85ee1b1f34cb45fd790a8f5919d4008f3812fc35640d54575cbed7b16a2add103d396611f1cd874bc616621b713e0c4ca3e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5a42b32fc10ed1ca380f52f8a48414958655b72bec364ef56e9d57406c402a416858b6c2b853f9d51656a3e18aaee1148;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda7f4f4996d0cf17c200b9992dff225281a89079f0a66b6fcf09451076943127e49150367441a483aec0ba28010a0ea90a33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf34d109ff828ba3b794831fe14a8db3e4a7c65fcc22152423e2a5b97a39ed861a93cdc1c0fc9c2ca781caa2f69a527ec698d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habffd0fd5a372b4378951ba342a055ad4edd258ee7ea7123390eb5e5a95e9963e1a8b1634ff633a9e00747cab6fd87c838c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8319d4c5b7ca7e2040403fdfb8e2bbf8c80a4855139ea7281abe860f5ff684ad25ec19fbb02d7e18f6d28d83c7252970be25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2343efbdfac5427d1bda65240c254f519f9a7b5444b3d5284e1e898e2d4c6c760468862f807043afda2efd9f5de53e1221f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96de38a41a7e9e3904ba07199e9748fdfa507e5989a25ac3b3a40fe611a24dd3d0e2b877428a5bd9974126e01183cd5d4103;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb4ae28667c15e64654c46c204c031553b63af50244f01d19679715e8314ca9c6b7956e22f6a08e23e2ca33b43a11a6937fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb24bfa06475285f2195ab8a45a8b984442820d71940066a63dfa653176788177526c9f49a78dc231d209b727709d0d99f293;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ef7788c36fa6334f8894795268c29642f0578fcbd724c4ff120b9ed60efb8f77b213e1f72ff8a4528e36cbf02d188dcd96d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98de60b6b613f091746c01fee083afa63c3bb3890599dc5a634cc88d33252e08bb02d2caf94719b76c25f32158601bde0365;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h439990230021b7ad1bf567571fe2b18e1ede7138b2792c12acc736eda69694cc5797a3a053239e66f086cdf78baa6bf04c34;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e9c38ec644750f3f211201293ee6af4b971378521e9d751be4c58ba2afd41d8096d2416a7c5a87359e8fe64aaeba0e5aae9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d05a47d6a4d27264b0ae244e90665876c8c8eef306b12978934c81992e17c8dc2d6b3a09b410285d546f9da8928558db07b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10fad0cebfb08b091b4416c5cb51bd08e0297341add5c642efd91d27fe569cda597b9807c17dfc275f5257d2f8ce2fa3a69b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f604336dc90c666bf994b511ad11ae8ae1f1cf29290b273c83a3fd1aa5acae816070e289f93acdef1ad93044bb1f198d368;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h249c45f233f34b636209c4a55a315730e13e1e299a4718e8bdd59ab984ca896457e36657fb074a6326bfd7fcd6fe1d519bba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h203eedbdd15d9decb4f81c3c06fecea03058f89f21b25df9d9fc4624d4a84ef2eb0ea3dd0cb2df445744ac8d733b71caee6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39714b24f1bec762705559825720401aabbfef9281a26e0e1ff69fd07713ecb030df4881c080bd26c39543dbc709243023c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h336ba554bb760fe4ed2c5d43ec2b3e8c6cfbb715e349e9b9a41cae9fcf6efc5f8b08b664f3cac7386e401bd827d86826eedd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6e55c9d7769536f3955027fca336698065ab7e867006d1da6e25bbb7d6dba2bfa052f3b28db8aa7b6f449b424612cfc3f6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h648b2fa21eae3610c50109febdeed4671588cfc7b1b2f5801e12f4f913839e46f662f833bca3dac6c600f7c126a4ecc95f22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he68e68df2f6b51f92a332e3b76859fab49e02dd2dee4e09f46ae683004fe2649e90268486315b7836777e58d426cc6a97d77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h839dd7f5eecb3fbec6a60f2f6cd52c6ed964dd6b1a3bcc613c2670c78f84bf1348a05e30a03cc86b64efb72588018cfb9dc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55ce39e674ed3e365cc0bbff6eaef40c8f702cc92326a057c1ef59a75e7e225e7fb3c97c3957984b9a9d328075a982c2377c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h873fe5568ff1817c5d36f7add6a80c749ac2f4045fd9ab614581f6e5e1fcdf24f21779964b460748210f80fda78eda020702;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f45eb471802e9433f7c8435dd876d524b2f48ed31a63658d0726c270a81f0c2e6a996b0ca1a3aec488fd11c6f0eece15140;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc834178e63c62c2987080f8ab25a3236465214d7f09f6964483e1599124490aed91c334824e0a808ec355c55e40de3be00fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a54f3f9f499937e57fcc3dfacf498707e29990e2040702eda760edf55f03782ae0f014cd31b28846f5a42960d12b63907fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26b30b880ddee90849487ca364e4bdbc5c2f2ab912a8dd0f105e4ca3613aa65fa3f15d4663b0d6670395fb663a2f16b68320;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1df44773416ac5236cb833726048982eab04884cbadc03ab07d07855628bdaba0c3bfd2f62965f2f5db5f96eeec81254a835;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbb187855e9cfcf6aecf10bc0376dde8bb81de3a7792fa4a508fb2bbc3293527e31ac67bea6006552a6db897d3321ed391c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0bbba5d1dcbefec979ffb24cd3bd03519d9945aaad77434cfa18713ca533d898bb19c0af46c725af8fa6e48768f165459fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39af65805d93c533f9bf17d907acf754095795a3ce0f76f2d8fc37b052dc8ba252e1102012860b14f6cd55e0e891135dd4a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf017b538b0120bb5e1640077cbacde3f8399cff3989fdb0134c512d9541651237f2befefd7d90cc9a17bc22b1c9a80f475c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28e753e6a203db402ee958e783bebe353dd976ea70adb129415dfbd8a58f15cbc7d050ba8fcb3755b7d6a3ff3c802c6a5280;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e9ba4844d79faac11accc60aa7896007c90022d9511750d60af9526ecf254df134c6055ed7dd3c7b16424257c6a61648556;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36fb38b9cb02732454757f8737dd9eda280423f0398bdd8e5094cb167189aacbe576bbf51fac771188d11c803be88b1c2abf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5c21f0f73b1db06dbe8647ff14170ca20eaadb08d657238e39226884765e9ae2a0e7643b8c21ecfc5495f5cb366660cab93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa0f3b9ce083f27fbf101f27e520d664a8a094ecdb3adafae12425487312e3c39766c4e7dbc82f5aa9fa9a2ddf676148369e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e7534b538713fea71b2707c6353243a41343b66f8ba0548ac652c37bcfd6d7bf9931350e9513079b7c4c28d2a11842db7a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h788e144102a90a0cb03819310be7bbb110fd033f7fbb564c104f8d1a1b3ee27bd43fbe1931c2a5d47b15bb669aed85c5be1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdff6c8ac7c9781a00109c17d8920d2570cae850b788685b31f2ccaa1c5c90dfa9e59b5ba48875bb0dd29845e519e1d4a60b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h305968091aa8c24556999c3bb2e83a26457a23a6164340d1ffaebe8ab15ead05b120cc0f366d96b9c1a53b9d78b43ad281cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf80c0cdbae2bb543934ddcd16ccf62b456b45d83fd1cb09d2c0410ae72ea38e68327a3cd1acf4ae2df82d15ec309215644c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea49937305c7c2233a4689847ebd6cf276a026bc9d2d344ec5e541be373e6d6933908e02b64b26536ffc2e441a469b04b7cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h176f6ed39bc0e456aefcdb6887afdc260ab8587d4c8f84497d585f090a37527402e5f3f63715bf037cad6b3278a4642a51f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha17980721df3106bbdf4b7dc70395e08b7d09d857c92ba3e49c36783a9b34fcf678978177cfa70f736435e042be9d203122b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9dff9c4be8086340fd82c34e5d5bdda9a8c82b70779de748429dc50d7e5dfdb3153b4c28730178cf2a546932c5cb0eb061e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66e40fd59f9eabfe6645de6c3d3b650b6c64a5bcc9a4207daccd9f3eeb0194fc448860d8947d646bc6efe9e53c699720c3d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69ad69e3908304c961c7bf83781b8c4a2d73eca27a6f9adcf8459b9bdf846ced32370001ea07bc915edd87cf6f263cd30d84;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc948e699af7cd911d1b43764282ead647cd0f219fb6c41c68316e554b96a611627913265871e13f2bf185cebd6225b551a4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21196d560b0eb297d3153ca828024f4fa1e131d02abe202d7492668c67d6d5d9bc2025a1220090100222c0bdc88a5e4fd92c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h816f7878361a83dcdfbbfaee9f3ac756798e7a2bf0fbe7efa54cd50dd34927cf0372bd0d8b6d6ba718178230bb183e434beb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he31203c77784a5b15146b7bda6fbef03836dd32131e2e9c8aabbb7b4140406ac900955c09761f10675266c79c469c6b2352a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86139c02b3cd2bba8b04b4d0d6fed5147cdb971c4b3c9d6dd75d8cd7b2b33fffedf5369b14334f6e579e940cd30d9e3ddbc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a95c2a5c4275bb73f81a0fabda3eeda3c1b326694567497b9acc381f944493f12ae57e9fcd12ca5e4092284d34f258e476f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32f8b8b7f380af1742a0d7102336d3da9f8081d3377ecbce8faddcde6d58532a5ddfcbf3c7ab3dbf1647f63f39fda47f82a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf23653f5a78529bff0b71c3078a6805fc9975ca48ba788b6043e298affa2bd39417d410e786f9b801e88e54d7e92510bdad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6acf2c2f08ad2a8789dfbdfd5787ab0d1b86ed7f21e03d8e78e0b6ad29e61ba075811c0673acdc6b443310dfc993c879d02d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74d3a8e722e41db25ebc5e07d64052f066d0304659e97eedfd370e8e7edffee5ff815ad042ea7425aa163d61afd8e8da9f2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5eee6d3b408cf8fd803902eed4220c0ea5202483b94de12c4a31355f30621613f16a28ba3c4f95e1c3ab300896b83cfa9e0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f8b6661ef644ea2b2bf81b88d1e23744674d03411895dee367b248d258ad481fdb8b401906080657504f4a977d7f6522b78;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42d06f92fc53d1279eea505e90b073a4df3c77b49cc347321c9e3d036f9a1ed8cc58460d0af489bcd08ed6f5a01be41e5c27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbda8671608196ba1b85deecc4931698631f6ae75e8439f7ed74eca722ac1f38478318a692c749323fe3987a6bde23bc22ed3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22ca55c0fe43ed869e5251746e75d85b62cd2ba17b57d0ae20367d91e955708cc356387e527d980df6b86c8a80d159152e4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc910366fb7437e5da40d7688a1c721a60e7dc41f1d7c1d4dc356d9b8d9178fbc9a028f13c52c423d027de58ffda2bd01c44d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1e70ed69f8acf70d4991c9b792075ec360442b0661333b36df76fc49de2a33e97d6e206e442a806d9cc756a760b60aa632d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe7080f3d7b3fe3770fe98f4f4a10cf65a3e946de1310b5fb8c4c5ad862485aae94a53e60581715e0af1e0b5dcc799e58e47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc988c5dd7da3ce6e6fe7daa55ed27e73b5b47209ff138d86a16dae5871dc700d8660bf17c1f9832c94a587f8b95586bcc437;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2b2fa4d5b4afaa89815225173cd643b5f2c5f3db403683b8260027775699cc2007e65396f7680d84dfa0517ff685de26daf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habb766449dc7a6df65142a55c2868ea2dca3698c01b9bb4d52f1af16ce2e03a6e1ad1c866ff7b880023a2b3bcca415b5ad77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d365ac652bd28f94ce54877dbd64b88f52aaae16046d92568b55af174d6318d5fbb9d6d9ba2917a88687aea6dc49ddabbab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81752b925c5e5b0970668cc08780183302fcd04ab57a94a5da0434e50d4af239d3b859dc5db5bc9ead2ccec211c270f5f918;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d330652b7c1d40985a4b0bd66894753492b8deddf90010417cd4573746e6294560b59eddb2c10e874bc3832beb766d3da7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h743ff8fdc63c2e49d30298692ec95bbd776aac67abcf428be166769c0be49c0a7b24ca5896a4c7036e29eed2a562d01c5d47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7735bfe920b0b08903bb82b18eda3f4994ad33b5d4ecee8bc9b84dbce57fdf53677c6ab9648f755adeb18b307df2f88778bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54ebb6907def5be127a5d9d8bfbcbf0f5e5b5c0b246fc6138f809e025dc4e8e4becb13834c80615a8cedd3e95b9800551f3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43a1bede15ef407cb592ed05ca227e6c882a003418006da5f9374a94c6c451983cf510604fb80fd3a8d4686f556560ed71d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee5b97e9f2a944008b6a5cb8b69f26fe3d514c8b9f8c57cdb011c06be8fa1a9b39dc1767f7f9f8afba5a4a44d2d61d5615f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ab434341b257741b7be9e08f7c8719a8353f2c7842054e67e770b3eee95b3d4483753e96418135579bfac0063d8012649df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82c4a4eb19c4c2475b24be8b319c724da1421b39f1517a6015abcc2cfcdaaf0c475c3d34d0fa4b758e6c4a167b285cd13454;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5eb3837aed077e903614759f3c772ddacac1d4c95276d9734dc366d40257d3604c36568db0dbcf513d98fbad06283fbf8df5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b7d2b5e7556df6ee7757c8338ab79a68f32aa7fe43f0428387dc42f8118f3b6cf073160a53a65b701b8c22407d6325892bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5798dfcd32063d40d0d0fe92aa1b567bd5b8aecc6e7700549523d0098cd7599f6ae8a353a14693ae7a802f9c4efdcb45e4f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb75ca7358f8c31652f8c69e9d4dd072f52ff81d947bcda7533ec03d5a27a261ae06b64dd6e1cabd9a4a6f7ed2ea59ce8ea9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef39fb1c7995aef2d3b30364a2e2db54ecf37b8bc49ed1f0e68990ab4bacbfcc3bd7e238233febb15981a32d6d3f284ee400;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8822f1b7f98f0fdb719626b8b4e509b570842caff778e1a93c1b2fcf569ea592243ff0e0015b9454bdd2771b622446a10dd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbae7e13374874ad2aa637d6c3b3fd92dc58204b768452584bcb2e5a8336da537a2f5aecc9875516f0c8f8fa035a0632bde4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb4967aa3a7f7056611a7213908a22a2096f3c91fbd180e02690e8328ba6363f56c4abd1203f3b8ca9e82e568ec2da3d2d2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haafb49c52c0f6b54d2bac54724a293c4f9d1523d24dd2c1689a7af8425c51935b7600b91f0a90db9f1dd081f86ed928da1e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49c09a2aec0cced9fd07a30c237b4dfc6073b6b112ca572452930f0a9a07a40e5c57ea7dabf4491b80fed970c71fcc748e1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h890063e21172e16f08438fd80f34ab001c993c8441ff3e5669e92e3c8876bd1b28929f8294db5580d1299a03055440e8211;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5f5b9c170f73823e017d415c8caf41de47c99ba7aa9436d913c94cb0909eaae31eff10713c98c32f82271567f980921e61;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedad82f6b81d50f3376451319e6af8503d90d76bf043b891e058a58e86d9e7a063d129170387b1c7cd0459dea57e6c397142;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70cfaf71a18b011956b854fae3358d6115749cd6c1174adec41569fcf3233892ce6aafedb69881649616659cd67ff927e147;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h764cb1b5eabb0ca7daa4c0ae698d6c7511ff897798e8ae58aafc0ea665cdcd5372ee09e80640449c9ca1d2b5b9f5398a9218;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd54d4a248ee4d8d56650527c9b5be6e1dfb0dec56dc82ea27e4ac9dafc0f25c38805011da6540b934af4d8a221a02a1efe16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf323c739c1952f73918c7da815df124c54f0b9fa6a9334a68d38694c56142f4ae9ec858e036eb1d875f78e71da56a2b210c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5085cb0be132d31c42f59da17c559d7a47a281fffa14c141253c4a8c278e11c5ea803f82a70502a2013105862b9a0925350;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab35dc7954e1a91cbc8165a5ac49826a56771a9e5c1663f68f8316467a153b204e9977745e428e3a8e8fbce329cf30705dd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe371ab407eb76f7e6a9c37f6f5849bd3e8d8f408a9fb5297c8d10212d21aba311466287e80bccd45332080e83be19bc6d65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a32562d61648cbedf2a4972ffa1979e51ab554c8cc681732d164eea5a61bfa8b5647bf5e6067b12946a51bb95eb9d41034;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88ff5d9020a97a6b3759b255a08f31c1f7d988036dfd0d7606194a5bc9da8b2e48d7d658ba7f0953dc142211ce3beafdd555;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had633936c17990ee70281cc3e7d3e6603333c49f2223f3d91ecdf5557586db49a5f079b41c67c165d8840734079aba81db6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c6f3fb14fa5b434195e27d524ad6dfa76d8e0883a94fd95b39c8a0b017eef66116181a30c5e8747242f7f5cf3830a4ec3c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29bf8ce8fbc3d17788be818dc17c3429873d71b7d400dc579641f3918b544e2b6f4d996e202484a39e886f158e1790beb2b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93afce73de0a937a84374b587904beff089756861cb210906606061f45e1f7c6de94a2dcf886382a169e1e0a0cf0939dc9c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b8e63f0c159b316ca9091da8eee319f1b9b18fb7888fa3ec0ba85687c71b5de98486fb0255e1d0fe56a85d12ad3941d5d09;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcde165c4423adf839ca35b1dd1a7a803ff359be449d353915a2febacadb8e13c317fd655d13cd1645795d9b2f5dbb15c878b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0f9605fd03f50a2e7f0ad79d1bf0acad3c2a5605db18e0e837b350870baadccf84a16e315e96d21a43c75a52cce7b294ea4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97ff4f136e5e7420b52d62703ec31a93955acab78469ebd61e3b13541395e8cf36526295a8ca02805b3fa29d5f7c17e90d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14c688ecee848da9634382a887a8ad3bc49f9f80e1fddd600071669a8fc8ef2f57a1ee9a7a3a36ec1527901cdf077f16d231;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h183f98ade07cca84e1216bb14395ea0ae6c430f44115dd4a6ecb36866d39690fcb6f5a05d98470076749527d2d2efc24d82b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77fc4199e88470cf7fb0b0c31a87dbfdbdba54bb41e0df7db577b1fa94552a42ec2437628df73711e11636834b68fb4796f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc440636ee14e18a4f02eac97b71547097d7fcd31aa0a62ea9ec8bd6a77ebe3df47872c41fb13eded84aea60a28b6751c793c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79ad5fae7be6b31cb88bc5d169cba5e44c3073db73178870ea44a2e0aead3cbae5b7993078ea01052f82b287e9a79a69ca23;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadcf21ed474926b48e1e3f9c95b8ee54962fdc155781237cbf8be1b0c5e2569aabf1b956587386977360612a2b73f332648d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85da342b56492d216d31e277e32513f82a3793f1e9112f2427ee27303a144b0101b34a9e85e04107f78f444235f903285b9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd64b097b2090e138eeb87337d909b1e1d7423ca5649dd5c06dc22d0fb238f4cf0e622631c188bde2f7020891902743202c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h277daa4b3a1ec74ad4c4ec35c3ed35ada4eab05c0267f57b4566ec4493c325d404f8f12f519892ed85bd46330a9a6178a1be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7925f7c963d56117ea269297599f777c65428a20226766c0f40afd472df92f328d2cf4c6eb06a7cfcca442bd566147b939da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bcee15c52b89f1ba9497f89e4eda86e80c8065b1e6e111375d83cdf0db970cda5c8bf67710a7fe0ac5200bccd6552b72499;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81c587bbec4484ae99064da58e5cdc894a248a1c4a4c74b2e86c0158b31fa31c13f83a6351495e566eaa6ed71b8882dce0dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haab351692091ba2744b9536a7202a0ff0af961ddb4da46c7fd8e416a2da70067a5a4881a328591d0e2c83add4c95511b42c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82c6ce7c70ee1b6cd5346a78eb92deff8aec5a9c24de6d0703a920274c8545ea6c9fdf7e46713d92ca85deaf3343496d35c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47e48af094d68ebf7aa7d1129864d6dc0e8f19911486432c01fcd53cfb8ad179d3f4439ffd46930cfdf6ee96754ea352bf5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae26e89a6b9b27536fd7d5743862a86e86dd6715ce3b07743c3fd114200f62ba08a426d3184eb0c671a25ceb12a45df053fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4413eb2c85aaa7022a2c02afa21c5fbaf2b54fcb8f79462e6e88f5801400dbd6577a9f858e6542021fd2df5f61a4659b22f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97eb0a219cfed9f71a9b29d0103dadf01b03d1d328c133f4dbbb1f2eab7cddfea509a33ddc7a2822ce5d8e539e05eac7149e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86115cdce19550e04ea69533b6b8770e685093e085fd379229d798d36fcc8e3f7c68e06f111918a1bcebf5d090cb9f7a2bc7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46e9f83be8dfc3a6b25998f726391aa3b221dab5f22bc7435a76658f414055894fafa74b9682445b9bef63cd46e7f4132bd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd96cdf983046f81760c3c4c5f5beedda2309b671ba2032b0446362b17d63be18363a82d751c8413b0ae5c49e27dd9ca66e56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9a2c68ccb4996a4da5049cdd1dd15b522e759d4d5e21b2256b5d59c20dbf4232e6496b67f44a53a31d481dd458bd2c928a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef3818f5c2bee3ff2652cadafe4464bac41470323f86add9ac8e2c570fc3bb3dd73c3909b792572fdd1dc0de96f9a3d0fb1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8046f5e79c7a35805478621946ac5664c5562e6080833b3257d9fcfcd9a63863f6b6ca13ed4c60083e8001a3de686186556;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d2b2337fa0b077bdeca8348306383c2ede0de1e6613072dcf9fe5d7711afc35dc78ced4cd7008fda934bdf67c2e6664427;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba5a36ff931469fa5b0b2767500396d00facc1d966ea2c9599ec942cff3918667b9b09f44738493d0b408a5a101011a7beee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80d256e0d86f731947cf134d4ce15288ce55ff33367da068383c395fefa783e21902892bca3177747d2ee8beaf7c12ff5fca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8f099524248ecce8d289f367ae5929074d872c55e038a1604ad1b056382a7ac08bc2d6c4fa8d0906d97a12c5995093bd500;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4374cf9da4d3cf3c4c6c9c0f0630ea1b809673ffa2386f4e245c84bb1f87d03e37057f81021ffd0ba2fa4ab0426dedbe0458;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6270de30fdfdb708349982ad0258234138f304fd1ae43cb4e72d76e0dd9b0436fc4f5feb267bd07fba68e1cd83855e136d37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha539d8e3259670727e31e7504cd9cdd4ecdb0936fed49efb72ba00c4fdee73230c49ebb712ef812e3f80662365f8dbc556d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha17a311faeee7998d20f3bd1cb06dabe2e5aa7dfbf0c5bade6861a139ee0df7f763a6d25e79a62d4b3828635af80cd804c92;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ab231e87a5cf46c4ac0f2b76e027eeee38572707aa4973e93afe45321d332b13346905b56aaa1985bf8b13eded9f9ad64f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf97df2de011bf774bd24db9cde2bb41eb161c68085156d70a891c104bee3cf573166f5978c0d9ab83f822b4018c4ae71f9cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1876c1f6e9b5e7a65727013e2f0554e01591554c235d5f19893dc5937c653dcb5bb04bb60417c649e7673cf9ff12b3bcc825;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc335aa21a573e584172347376c7ec434cd7c569e1249efc75c3baac8b473a0746f2df8783990d33ed5164357c95ec51d923d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6249fd94833d807f24350311010b51a5ad6c33272bd15a96e50122b864d058d577df9043de938936e011e7ad33fcdec3030f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h236fe9111d49a7705da4825c10cde3fcc58c9762a179e414ee2ee5c660906ee915a56ccafb1f6f7e1033ae1e0db1f7fa16a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha35092ef7f9ffa6e8bd2b7f1dd27429b34cf6e733567d4c8602bf2ba88509509b95fca338b1258fae801459fc4a91a5a987a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95c37e8ac0cc19639b76eaf35a495436b752ef3ca1eebfd216417806986a35cd7024cbea7580a9c478494d9cd6494178a07a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6146c683acbbb18e0f30f7134df11771df818c15c1e64c3ca29aa07054aa08c10bc534808c1a1d40a646e1664796ff1fdb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9778e90e0f35ead41f4d504dcc9fc857a8072e2859cb1a74a31c52f002135994c7c736c08257ab50ad920784871b31572314;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6844e7f7408998ce408a8a8e97fbbc8c7251ea76d324ec22de1ec1b02c3455fc74eb692a1541bd4f2c8a354d0b2fd70d0b1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8af571787314e625af256594899bd388830c2f75b882778d4c43e296836efffc28f64a51997bd927c4db523e4830df9ebc5e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84a976cfa29127186a8af948a0bbde577e85740be4706901d688e8836b8bfbf58c87faf81c0b3916ba4ce4686c27d82860;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b55e461311b9edcfd20065a623ac6ac4484d571ef3a8b5f37f1a949b9ae101379fd581db8b6e90df7881a9cdb5aa2ae7f93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e8b02afff3ab73f3513036a6b052b27ec7c50d16d5cf8f84252dc202e6a05ec9b0df187187895d302bf490d5cb437ed472d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb46b004755203d10c65483c19b08beee0121ef7fff2628fa988cf7a5f4742d5c8acefb8e72cb6c367d2e0645e1e1f3f1c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbc30341075e450d71bab1658ae0fb28ff3cea651ef60109f285b77669a6b6b5a6957640fe9fd0a6820be1f3d1053f6634f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe6c7a34cb9534f5ff504efa0b51cda8a0e07f74808a3d31661a4c7d9ea46cb61aaac47e3b4eb1c93f1d7e1d64528cfe7360;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5dd1ca10f0903a108428ded2ffcff8d2217130313e8cebcf3bcb47a0a64846c1aa142351acde8cce0ca5fc7c272e808fe8ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57cc5355fe679266d34767bc565b3b0917e0ede03ce408d056668b9a7597d405611ac3e14e29cf549b95ccdd5606e6de935f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fead1ac4b44fd7217064d2a72b9a8546a2ade3596dc315c3b4b23affbc29175cfc6be4dd050c59f2a313b2b6018988c3f76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5d1cbeeb8b437a647d82e412337e9397835e6a81303ddd8c4422627ebdbbc8ce1f8e4c96eac4a34ddd61bfaf7059c20f4ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95678c837486c1404a67c90544d01c0c57f0842d107abfadb46c914ae06310bb1410ed7847c5bba077f3248c3d38a2c69427;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b1319c308c9688c23413dea077bef092363bd57edbcf632c39399721221957d8a44ee13b583caa842caebee1d165cbbb99c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8f815739afa42aa839b9ed522491a9bcbc93b70b5cd9b6d1548f13d9a30ed6952fe58a1a13274c0512fea61f94c4d675ead;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a22d6b799b2e72c8e86fb0a1c2b3e6efc8144d9486d61ec6bf7d008e9bf4d18b9626b8de9c11a8924be41bb83bca8d26416;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27adb83a635aecc0a6338e29656887e3961e55441bad2d2f44f08a4536cf0b09fcf55bcc6c9ecd7c6a780a4a1b74656cf17d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfba158d4e4c4a1e5a732e675d1dd5996b3792f683023c14588bba27f26b28f32d60e555c74c8df31f32e910d5e9120fc7b6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb7d6398c87cb49b0f10cc75ca391c558e2face498b614f4d3a6a2b3145a44163d7794634827260ca4833aaf34fac232134f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h871409f7fd25ae966309b603a2951eed8f0b030a6befac714c2f84f6a6ebcdca137df2c3ae3b1267072de1575cc688442f45;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf4ecaa4f2afa8ceb635069e4dd1923aa971a17b6fd501d35480a720643aa5f0b303218530e969e299eebc02b3d6090f4dbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1e2ccfffa581b82efb44af2b65723c91e4db4f50bf6eb8e7619eff43cc86e7a02af53f8bbe6034bafb5e8e548b472418934;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f9c56ee11486e5457f016410c8091f32c6f7d9f892ce91ff1a5faf5955d04eff821437674c8f9bbe28bf4659dbf96923fc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12f365117e511ebf0245d3314b6716359a2ab10c2dda4846f8fd61bbbbf66129d5c42905d3ee2c780bbf0d9845ded7cdc46c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3abf3a8994b872f0fd2a6c4fd8e328e7f0f842a28b5ee10ebd9d7b4b257c0314bcd1439675b4f292f106d302f3ca5d8da99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2accdb0398f9e6d3816b388bcda2e9f5c2c52c5aa2729c1daca29f938f9504dfcb109530f6167e30c816f6785ea4dd99305;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdad5db4ff53cf120f1001752b9fbaa52cc7da2b29857fe3976e76508bb80b65a8e4a6484b7240f62c450b51f09b61f3ed5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbec2a7932b06d1c33bc41115d30bd61a41ebf5583b002b6060945862ff69682400e47cc2ff7cebb295b966662e0f460e7fdf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf17958c1b93ff6455787ddab3ef9d0acf67c69c6556d93c9761e0dcdc6bf8c5844c878fbd4230e04373d5e724a861fcb3037;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf601466ec1c32ac74d68f0d5114d942e1f73d75e3faf3fcccf5716c72764b9d6aa91a6793db2d9861ab12f5440f949c8b32d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f9654e9ecf4caa19d1e9d9605797a4f1f40cbe26586147c96d38e77e82fc94b235f78a0857abf522f5d5ae4e49f175269d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a676555272fbbc95b979f82fb5f27c15a2ca47c967b6ce4af58d421a12156ff568733cb43701093d7d72689dd0c1095f88b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54096d183731de086e914dc4ccf51e8088fd6ab6a53f70061ca5de5478022e440ac18810b39042183e64b668a2ce8eb0cc08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fd9e1c87ce75976c9ac2ba32fbff1a741160c4261df2dc18a79d976574e0162f8d109271d7accc83e21728ea9412c151cdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8c4f977be31de6b51a4f4d63a2e1d2d2bd8b2fb848934a941707546e0599205dcb338207a4170d9e5a24c2a3b0cf0c84f1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haaf1d07ba6bf3bb14256d4bdd5ce6bdbd99af60907cb30b713d05129930b66fb4bce1ed08e2b61daed916bcdeb02459df3f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he419c0c56782a5a53c55084c9258a1e3e2be0313ccf7ce943e2d66fbb51d7de647b2d7a46eddcf10c9c3ef532493e48e4eb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd306ce3fc4bd340cf3d48a00eaaeb8abdd871240a742021361bdd68628f4e1868403d1cb1cb80019cd20146946b1569010d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c81eabf63b5c528f4921dec53fc4b28225ca37743e127cd964f46bfe01ee4d624be375db905715ad4790ed726209502568;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c50bd74e8258c53a4b64df4f27b48967fb59f554b84733255bcc207c04fed55be5df44c13373673fc72e6bcf4f609cc4936;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e0d16da79f3f2503f96eafd9117e0c32145665f410cd19b944dad445a6bcf0f43a93ad6e3c1c19095b36e6ad9c4fc66ae98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9102c6019bb3120aaba9c4a1913711c0abe4753d5d3d6b6b82228ee1cc82a9702920ee0c136c4b84eefa7a3f488af9de56df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed62d386fd71146674eeea35fb1d2bc574cc2615238be222ca14410e22c05b245dd765e1b37152d662daa6861c22891fa870;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8f10a029ada4d33ecdc0b0850183a20e88deb623a080c79d458ff6c06b5a05588708fec318e6a88270392292ae91590d654;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf5529fb3f96c08b78da1e307a937bc0f7c3f0e09e54db876084f16bf2dd972372a081c6a64a658866a085c7a19464562f6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he49ecdcf3afd7ea4ae685f12098f5c273ecb4c336afd2c2048634fa8f914eb26ea301c138c0ee682f9b4c84fca30505502c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcab0deef56ccacb8261ede4d41d4138aaf48b2fac28dcbdc9d14b3706b850d42c38b3d9acb18ac66722caa315f74df1b91d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9534a54cdb426ae4d14d0a501790ebdb7a8350816dcc47313e163cd3db77fbd91d610231b942ecbf32229e9ec8fdad322a13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf0942123aea4a3e2bb07734a843670dcab0a7f0cf70975e1ebdab040fdb79d5babf068d7cde508be80f875d0e6163c9417b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf5b9fc50fcd0dcd3a3b5728017d68170ef0661ec8b67d5c5e881d757e276afd17b4474b5965b62ec588e467a2a334f82c67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fc9dc2c81fe54ac7ec8b92b75614d710c0ca43d28b26eb691dda0b4f24dbde1b8cf26db7026814e982354203bfc6d3f6288;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92bc6b4f901a22ad4833d7a632bd9829876eff4efeb54d2a5fff13dc4bfa709f2e1c9de20d139cb832f852945b3994da2c1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27e65920b738341995a80ae26a0efd37081299164ba3266d755518fd09d4e3c6400b925072c1330a7b7a0f55ababc9f18291;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54cef2aab6b013421934f5b7e9bed2b1581a4cb0f7951edffe7f92ec23f3abebf612625889b9a5f17f32e1a6773e12d33761;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ae8cdf178dc4e375c8d695a6bdab936a239589a5eb476ca8bdc3e6848fb263a3281f5eb61a447dd9d5ddd8e804d52155b47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25db52d856cc182aca9b4a3f9df61b700c9de6c5814e1028a2cd45616d44f1e8e82a5bc7210a7a79c2ba852a2c6a30204bec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8eb4f1e30983a8a6704e2cec1b1d383a9889648e297dc0b3f3de41682e76a32293123e847086916d25eb4fbfe50da9f19140;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he306cc54e06e74e1fd8246209e61996b9bde67a8c03a87d346207b980df1b7654c1187933971f1fbae0c961c3110a3ccd8ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha44efca127b4700a643d7eabc3ba9c204de1d1d4e7524bf359fc97ed409f6ec57a4fba5faffecbfb6f928157abfb87975d57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb740faac2cb2fd3ba8d60ffad5b483ffa663548b9a1322acf7f05be78c78c659e879d71870f9515902e3cc7869b5b4b80a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha72ce480df1d10bae36ccd910643a339bf2a110d42098ea9d2ee74e3c20c34daa4521bf5a1b06ad595d505e90272c5576f0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9a145a9a936e623ba1b71a794f854b7ac49d22196296ad1138112fa511fe3b38c723aa9369e84382af0ef451be49ff9038d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he84339110a8f1dc695618cee82c2df0d635f96bb4a2fccda961bcc6cdd599d1bd2a30bd13ab7b01402bd79299f899062aea7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6f3fe515abc30ebc00c7c77004af2f7abf423253c5f2b6c44c08f90992519119883ab6f09cb98682297511a253fd0d31f29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9febb97f3b73dc61d1182f10fba1662fbd4a7687112ba44fa42e07042345334699e0eb3649688a08e6dd85d5f1c2ae7f4827;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f023d41a7cb4c7075f1d1fc2573a9949793f2e07f7bb632cec6a7d94b602b55e78f7a2bb693b736b0bed18ff2a6bfe52bc9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51afbd2185de26d482bedaa61c91fee7869fcfb2ea8a30ac27b88b1b91809501ea950cfcb448200d99f8379b31152dd0c048;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3e0c57bbffc781479b0ae861fbab7eef00d8da68e703b92301a49857c0e3ac8b77a0155d8df0377f777cea55e6b958b57a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h321216f44aeacf599fa44d51f166482fd3928e4476077e11e168ba0e563260ac621778f926b0f80d5399709bae82e349d32a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he12576b1d562b353c23f3a6b85b38fc94c6b2ce5f448d03d4dd99c4071fe64ac5c0c849fdaa6f0d83eb9f3602c51c0d6e66d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4917ccc9bc1fb5d8dc4e6da9f0a65fdbb75aa9a19b9ebf079530e464298d0f9eab148cd1f53d032636988a6b011a09638078;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38713e8754a4e91a2d8b00d17ce2dbf8e65efa8b73edb8d02995029ee4fe99f7dc486414b9b05a0567400ad2e1e61ddf919c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb392a8febab36cbd9caf9ec1b10cb4f4f06e619a99f5a114effc7602ded69137cfd1454a70d4daa0f3efa367e17d02eb9b35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a18b4eed0928099888bb83bdbfeb9aa9e1986493d2b18014949293e615a552877f7493d909e02e4254f45734dfe960f7146;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h880824fa563c444c562a23af5aa4a334c24e656768105a226fd34844fc6306df5371e17448a83eaf6dac69e399b281f560ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc77f8780a572cadcf0a64a6aa3df2284b020caf00a03c4b800f394d4c4cdf8c5075abbeaac0edad91fc5352db9a92c14f738;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41c86d022ed0a27c48be11a8985586d5a3647c3b2f660dc4f85f54c8e943a8b206e1377207c6e94e68809bf625953646edba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4701765bf4fdd044d309bbb04e19179d27a0aa598f045ad043862304a21ac08817346205248e2259ee554933646bd80b3eda;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4a6b6d99546504ebf73ca9022c51d615f7e4e310ee15fd6de5b30c786a5104311adc62f744a8bee96cb7cdc7e3daaf6cb70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf71d593e0eb1101f6195b1dc2ab03921c82261d7fb81ce3570c55834a07b293b315a427c16e6b740c460632a0f1e3c850e2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf449fb7bd773c412d8e4aaaa3611020907cd1d114cefbcc6a4a73a82b2df36327348c2417c1b52f45d55ace32c5288667ab8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49e86b90b4459614f60e76d56f7226bc366fb1c57fb14275df3127cb9965fe1b67fb74156cf8ac12ba5fbeffca806bd67288;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b740f3727f27a72ed992c54585ad3aca86a89c465a6ef40a096862b6e1b4db3139912dc6f3d1a5c34e707dbeaca7ead40f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36369c3f708fb8bb246d859ecea533bda7bdca7299673689cda6079c1b9cc6591a1420ea24dbab59ae1e0af338fdbc12354e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54232de1227694367abf87e3ca5356e8d3b131ddf67e970137b99d30004a6bfa372ef368e7c9976a467dd83d32ab7c751a03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c00e779ce6573f64ad0f32d11f8d01f074d0831c90012e570febea9784c761c49bd7bde01da8e564faec990d41684b6530f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d95ef8f3a214cae7aa50e61b34202ed8d836915cc672b122cec90918360472dbb186429507f20200f1ad6512db4d20980ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fcaef97c38c2be9d9904eb041705c1ca046efe5b97df900e5980941535326bd4298ebd4dea75769ab870d499badd2726bfa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4fb59601a66ea5cc8dba417878db2bad998b50bddb1dbe43b171a42d58a9c7593bf3a222685960d65b9f573633ed0301276;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he05e34e26d6e7cf3707fc79ad47502e0c21fa62679810d309fecb8735387a9fb33ada993ca3cd2e0667d4f0ffbb5cf611afc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbfdd9ac1125326f11d7e2b3a7d371ad35cc56ef45d015d852951c22dff1958a5577121eb710f52429011ce6ee4b0e25140d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf99378b1580b92f019e13c7d05b7566f0568ea6cc2fa56a3a92772b52a38ef13faf0906df1c6b07e0fc2b15a3271a2ec5fbe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb3f3fc08504fac55e528536e3b8b6e5dfbe134e4f0e13b49f937a0df5bc24708d3345fa999b05abb4b832ab50c8bfbf3fa3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab0de753297cf97acca5cb7ae8e35db362f13ce6035e4f6ce686927d270d66f7b3244ab4204539c824fdf979d81af0137e62;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb08772d1244abb98fad58abdcbb3271d4751941f2fd4ecdc748e9d41850113fdd159681490880e999b895252115dbedbf574;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcab848b9235830b5c310f365f50142d2d4681707a2f588227440bc773d315c90c20780776e87cbf8ab66268c44c38068535e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26cd8555c9e557c548a7fe32bce0560cde30ff747361bc8a6e164728c45d74248cc9b6b4e43171dfd853ca4a3fbadf26f937;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha54c593e8b3f94213225cef0c83e9ecb3bb8f49903de6c07f91a9fc4e4ab1b45be9d7c614a3df297d9d95a263b4db2b3539;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f0d9127ddf0200a4b06206372127d36d61971a392ad7cff5ff5b04e9bddd5fbe615916079f36304abcd8abb00d3648a9d77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5143eabfe728812103c51041242f5bc1ab8a9355b7e7d33928e0803458e007931ff4f6c40b597f6f62e94f0ed72c55891925;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f5152e3ef8046128e2c92311bd42e07c43736924e737f10aa54efdeb85f65a7636b0fed873d5c2e1d5e6a4139b660abeb43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70aa582cab9a269dedfef760b455a7897627d1b2ca10bbbd78d78e84388e882c741838fff107f058d957058ab96ec9519590;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7259471e5600fbecad00ac5e0c98b17b19a84e5013b204a717f0860fe15621122e3ff83808553e94f77f23ffa6f932235b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc91f8d42950e055cc0fb51750d0aa41114327c32799f239e2f87be183a30b98adea3b8b7bc519d1b71db7fe8953b60f38b2d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6461ccedfcaf858dccb95910878b7fb068d96870d5099cb7a92a26118795ecf7d661dc833e5eef4fa6259932ecbfa7ab160e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9079ff29902140c72edac877d55267b5f55aea0da5477a89b553a44d259732301a213e4747ba2c2431fb5bc5cae71da917d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cc4186a5862e50cb60a613b643315d2c6318d6d7a13dad9f175fb7cb65d522aa14b845f9512eba2f3548fe1be3eceba6974;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa967011024d1f0fa540bb3b4cc5e202cfc2fdb63a74707017e2296586ada38492527919f4b1da7769f15fd7711c7cc42d96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27f99d2276f438c7316afb181a43421e00b010a0e62c97573dcbcf11932eca31ec61d6183e69a8048226d99670317ffdc3a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc007536dbf8e938afc20bbc6ff31fee371150407b16be49aa1187dfbb3d6204f80b581c36bc610f12e5cac8ef4424e1972ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h837f39ff725bdb1cbf30aab84349c25d2c86ba64b5cefe74e27d409a36f7a6bde26bb38d635c0bc6ef93252d603640194c4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ce8b86dbf99bec44d9ad120bdee5cbea023957224d9214a787f30359c78ac467ca29c90b87511547570b9a2aef86c998720;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c412ebc47f58d2d5ffe1b24086bf1214d839abed9bc09529d3d9f144b127731996344224745327eeddc1f7d1f90fca0c5aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1e3f76d36e41eee3643300b0e085c70bbd5d397c51e0973f794cd58ecf928a56759435db14a11d66fc3a46ecc309951b4d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a44ea86ffcd566a4932b3b705d2eec85f905a3a8d1431991ad1b009cc3e3fc35500aa3cece5aeb36a3fb357dfec2ac1b20f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c64c00ad60cf9110c1e65b438221cf4a6a2e24ae32dce7e4d3f6a8c5ac5f75a2efdaf8b224de7bf3cb3508b333096bf6b05;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf2e2cded60a22597b48869d57b0a302fcdd898dbcf48be58e01e5618b9e72789a885a46dfc5d4450a286894964781ae468a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h489191c805ad0a45fb9a073d75750436c65e249ae613e2eb97aa190a29afb2770d5ab7f2311b43308f1286c5031c415b604;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeacce9fbd99992df7db7d78d0d6153cbebd804e89abce7e4f3405b2b524114270025b8f0701e92bb934f2fc790209027a45;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1ea8b2c5a22478b7c8de92baef35ace40f71d03bdd733dd692f5362a364caa64fba5d0bbee147ef925655050ad38ddc5837;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d666f4b972225ab4b7f51c5431bc94e01445ea5a42b13dee24db2f708d49b4974c1557602bc3aca6f4e0ac7c3d430157a27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7c094476a46deee6bb64305af7f77245cae194a6e3b03a375898afe1099e12a10d01ba2dde650e90093df8044d15d9e1eec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd636cfb0ad4aacbc83646e2030cb29fd246cda8a84e7bf7f23c369a1bf2a9e993ea3e99291c9b66e75bd885cae590f755737;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f8a062f3577f43b28e0695d6232438cd3b6b904d76084d5417ad0b8c159f6db9ef1295be1c3ff9a8bc4a49c82eda2eef554;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2723b38e49685afc9d6528af762a619f2166f66b4edb6af154e3fb705215b348451fa35657b57097459a040c311cd2aa95d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h753e90976ffbb8e0d1b878ec302127ba32f61fa0d79935a9fe403f49c4de23c0989e28a278cff5a7ea7463b5369466d8f33f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafd9dc322885e10b1ec32709e08689b467220c090fe4ea59e881efcf70e9aa016d182f99cef8300a9eaf43d7497948fd7b05;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1894eba2357b33c79abe93b9ab27826a5d146ec670f28713494db67a3427e131bb5e9764f3e270260ba4cfb444ace4e9412;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bee244ccdba8cf99042e905e8993e93372f585863752d73355ea6fc70257ead2149f9f614480733829804769c04ae5bcd34;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fcf63313201ed634bfac71ea91f64fb59351061e3423124417aa1bbbfec9f8e5a0d797815bb963902bb88126a25a55237e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20fa0553cec82deb4d4a603a745e3bcefa50e9de20223b79a5c3b7d7235a519f1c12627a8274297ac52877aff6b76488bc1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78df70c4fb6f0f2cd7467e64d2fc20fdb43ca952c27ea23342782044e779a43ad7dc81a21056cd4514598ed46da48af68d2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50db07207446cd5816d81363935c99b9ff8f69e78e7956f8628b6781775fe01221a63f99cf30a541e5f53d311150fa9a6eeb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he84371365ec857638982907a5ac5919452156684f6ffa4fcdccca84edbc0aa341de1346a7dd795724640ffe04f1ee80d3bee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7415cb64ef2fab1052e99055a72207dd145330e69bf527a4adf2201c3e5665d58e963413f08c2ca9d13e012badf414af5ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9277dfa910cc30166980e2f409b9417f613ec66e26d805e1228c68d84c0633049bfced4b9c9fe66482275c78a29e11421dbe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a0edf243404387df5240e78558745d14cf51580bcc0a0bf525af461f8f1ce475a3dd6a4d1747b203ca14b3ebe33f7d05ed8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4150872be92a5a9eb6db9ba785a46fe2a684583fa7a6bf4c5da01c6395f331f0054f9ff222854b7f915a1aa737434823817e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f521619552b35ab360dd2f3352b771ca42a4691e175f602900d2af5aae60853ff0ec48ce30ab4b4e7ab25c9e6571cd9a55c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc692a7f0d5e9b86e7b49d9e79c487ee0f0d4bce48e8e8069fd8d9332796a8456b81b50241825593ccbcc1287d929adb1c4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c2d044fa79930d5f2cac5cbbfb5963a692903a0accc3679fddde72ba34cf1ab44a75c0b3980294a7d6f9682ffa06c5944e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h691c80bc7591b86270b0f64c43cab0e35314ded2941610640c31750fdda9c87b2010096b0d159dce3124242d96fc7d42f743;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d45d861cc455c8d63d366e5508f350315751bb1d08b0c83f90081f1e1b474deadf8df2c20757ccadbfeef5e63f710ecb74f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88569d4a5c9f3304859153b9de082a97e9e9ec5eedcda0df1cfd68ba94bf62e4f939c72cf60e81ffe8226c9cdc1bcbd92fda;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d57491ead04c696fd0debdc38229818859262804b6867455cbd1157abf7ac1798a25c966f77cee3bd604516cbbec85ba884;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd733176f13e33af041e768659d539c42767e802b24a8fb617ff6e5868062294a1146b80dfed8eab0e511b9157437323ddfd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h423de25028d7dbaf58af0d1e4420dc8040767e0ef0682dbdd25a04f1d072245aa46e99cc6d7383e2f82754bc6544359cff42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e7d2132b10d84239b508b9c7d16f60a848946a391661adb14e96e0140d18bd8b1543f84bd8049f8133684e3b00c9e012;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44b93d8fe5846a5792562346949e43e67645e229215326355e6dbf4dc3e4fa3380fd301c8ee3aa43a7a0cdff2fcbcab2901d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfde7d0d1f5c286b6127c5ab23136d42160cd411986d17a19d87141b5ceab35c222df9601be1e33704e5692bd812aea5abf8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d5110d8c69c494175371ce67608a9cc9c2683ccb9d4954d80812b6d38c38872d7b2669d7bd860ac1cffad3e987f1e1bd528;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f39af78fae4ebfadb5e717d9b3040dbac961ee3df5d413fd15f75c935cf01dd342812621ca27f633eff59e9f10ba29b8a2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d46d3d34607539a15f17a87cf6b3d8641f2acdb4d027a855c916e41832d9afb406373185f6574325c8487036adf97e196a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1ec85a45668a28e32abd59addfa93df58a9ded48d1e20e8d07251f4743bc0f28b7cf694fb661a06f789caf34f0ab34b4065;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6b4c21ae1f3bf7ea3fbf64a0a120e52e729ea196001ce5a8b466d321e4bf1ccdba12eb3850f9c369e3c37aa2cc839bff8b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcca177fe0b6f59f57ed6548c3ece732a87935e8a396bec2d2d0f2ee9f8d765307f5f76ad480d59e987aa1d30830e91d1ecdf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heae3a175f6735fb69e5ed8d72995d468334c804f568c498124336316101e547a533d738d92fd5acfe80907ab03b90919507d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26fde0fb5e0f6fc125cf9d59709ceff79f26bafca41cb78cd7558c18fbb9548891082e63a712992982d9aa2d71b6e0f41fe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f21d8554ef0b2f70f7a71872b513f87a96215863b7557c634ebd3ef036db4ef845b05e6f3dfe119f1ffda209e76740c5805;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h313a1a8113bd1aabe8c1de8c8eacd83490c1a6ba85cf7713c93461c6690cd9e749c7fdb059b7a451095ddc97bc4e48069694;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc533c26cb54b4244f089bfee925fdb6c7f2c8a92d205c2d252edae8fbf09ab4088e83e1dbe74765fba0edce3a4bcfa87eca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha248e2cb946858834fa2b87acd91e059544fee6036e2161b56dd9aac1920490c3b14773afedaa49acf32077cc6b891d61fe7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aa7f3b1f9868514af7012b2941a34fbc66a7bec8480db1c574f9a262aac2a929ba3dfa3d22d21ddaf0a5faf6087ab451531;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b9d72d1c0edc80d7a86bda90b16b7280a613e8288cc872fc727f9ff83c3759d835795635c200b7064d7c0a628640abfdcd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h594946924606cc2e933cac9e9b61f434da4b205be822ae58b765c1b2b760b3f1d7c7811d8179395ba5fa6dea3559eb08b1bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cfd0cb1c33f195d495e6e1c3defb023faa551ec1366ac4a301c83d730da74d3def2e715461df1ec69ada215991ef9dacf89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c277e0069a62a4b31e4f7ea1d4163ae0f776eca45da71b5603a5a0fb58396dfaa683d977d48b924a41b1bcd7255ff61a800;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h670db47cd572f674451b5e23a7538f3b68086c2c1a3c5b3593a79ad4fe6c3bbf08110b6f44dfbc45fb699e3a466aff962746;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4666ee7f7da60a8334f51a9565e60198277fe7d38a3281065dc7859ae57cf9d9d017f92123aff13dfdee026ecffcd41be71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d391aefa58b32cdb13c9f9201542e3dfc334500b725c9c596529698f418200b4da7405bf2fe63409d2317a3ae7a7a023f93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd1292b5d6cd6bde51a7ccd9df230f64cd30b49ffef8956b5cb18b2098144991098a38bd4eb689e8dd6a0bdd8fbed03f5c4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b1f0cc2cab0bf01751f4180fee328a76732be9c74762b0bebfb8c7d6717e44ce62a2609aaabd5002c80db46407c9503f68a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e981733d9fc365cbbb20476a79149eb32862693635ccac4a88c000d7c91193369625de6ffb4f016aecf2f20fe8fca39e6b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b167e33d2cea0649f65d0e19b0957c51c8d66fff036a82e244c7a42afece591c903cd10a373f1447a9e00ce9128230d0593;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9bcc6ab3a7651226a2e39a3e8ca5978c928508a785d3f11dae9632a58c0f24477da4be8025095b649c64345cd75d4f5a96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbade469fd3d9fa3d488178e8e83c51598d023c989802ddf9448e6bee8d6f72a1bd00914d12c5e7f57619a123872213c8a37c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc561853e27c863c644ab40625ff41cf538c7b2412ac9de1ea76f2bc08d9ba740255761af6d4d2831c976bc885c608c25242c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81a1272089ca73de9d590c12b24fdae14f5df70dd0d98e397cc2dd8e1be9d817e245ff8bbe1a38a3c26cb764dbda1289726c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87f952307f75aa184d807e5447917191dc0e74e2e605377e0066ee87ff7ee21d20835b1dac4773943c0f871280383bbe9781;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf48e1e6d8fdf18082bc3ab05b5fdea71f21cdd66dbdace48c3bd12475181ced5a40d8180739c4a0474b8238aae73847c18b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdca33bea3a3c17a86814f1557f3cb7c6cc8e28d49aeecfd681cba1e0889f988e46cce6a2b5c1c50281a779ff90710fa152a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9fce9aa404df43528de4c45e465e446faf6b704386b7aa4d30a7a485207a9c9732274581744d998e2802a0544bb964646de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e778cc2af12e7a4079f2af357a8f5e790a53c8f47276e70b789fe23751e360e012f6c90a8777909867ea5a7e9b14c41b54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb59fde0fb98689919847d051a2c35e0413cda741ecab8cd33a0a0ee09f52968aeb3fe4a5fcd94c7338b19a18cf91350ae96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32abace3696483511089a3cdca992f59315e2830b386ed4b246c0d07c32b61d7c09adf24b10ca502aedc1b72d736f3a3b021;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d260097ae30bfb440057cfaee3a0a26bd3e7fcd2e1dc5b8c9c0a80766ca809c27da9ec3dc82a39ac02046ee9916934f5dbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cd73ecd5ede345041a9f68049d55d7a62dbff3de7a5c92df151cfbec77a0c3a6890ea4f6f09e87aa1679d90c126c6fc25c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd582b7395853608fe62fc2ca8c0a319cb6096ce919182d7d905527859f480435d6b74723488d094fc83b61ade41fc51734f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cea156db95d7ae980d7bc4353643c35f0df8ebc0b5f9f03f1ad172078cf87f07488d8297452879ac15f778a50ea6640ae97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ab0972513583d01e11bdf05d70acbeb8eb2454fb63eb3f03f89d98b5f940f124c56ac4ff9b1f8471c24e9a958460018f1bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc0dea3261b0e22db717d7889d4d9ce432b8d7cb1b7e7adb8eec60e8e0cbbe198781d50fbe44419db830b2640ece4af42875;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h912d06074eaca4bfbfdab9ee83fa745319a8273bac5fd9ae43bc524567e91711e6fb6688f751f82999fa9dc852fe5c795a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bec44bbbac91aade80e98224ca444bfef405dbb10037adcb30da5e504c3523ce41908acea516f59ef32d3be6d5214f86ea6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33c44f25256d23a4d7f837a6922918f9ae5b4379bc2f29a5bffb188bef045d06471d9c00355974a0594d55c7e67e6adc23f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf969fdab1c7323d922a28980b82b1188bf62f9005e8670f98e8ef5d5a59e54d8c9949def826ff3994658af23859852897690;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf41c9bdb65c77406fa51f08e709467935dc8bd13ae615003b3254801aee651805c02d140a4f4d0506e4ba27a618a56868099;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79f688e2716f4b7c39a4da869a2eeac83aeeb05040f3ebc821a7f539945021fed5594fee4198f3d0fb7a99485ae6cd86c7d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fcc4bfe2d0fa62c19275edc9ed72d3091cc61ae3db884a8d1386de4250d0f6d4b28940518e2a116eb5b3b1a31fbfdb6e69a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c751374c9ec07a5fc7a2acfadacd6527625ffc90a2011b7cfbb3f66c2a1b428cb6019e099318c231d24b4351e8dc3613b16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc41daf3dcfc06ccbddbe532f0ca3911015f17e5f2965ddaa992f24d67bdfb8585be09af2c4bdd4532370efaa25d01f277339;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb951c46f9abc74ac3c7f491eff30b547d8e80254f8052c4c845cb8190c9bef854395c80d9cc649028efce2996fcac6fd863;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe3f72d292e5112377bc12d5b403913a2e8144e643bcc9a92c0557058bed5ad82a3d75fabc5ddbef5baa28e6969d39b57c41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31406503358421f1433b1ad9334549a5d7af4a02d3ac3dac280203408fc147cc0dd1a4c03f2e43d3095c7b1cca6798f19d83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h224d71eaa0a1939605ab9bd9dcc03e68019d95bcf19edb6500c358f681cd1b50bba5755b4044879cd552fd9985ff5eff64e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he70cf2f02ecf082f4bd905f3f3d1c358e20adf3809c42043f5a3e0bb5a1dc68f7218e69537130bd0e13308c22e794965c5d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ad145940781889867f788b1edc2146ef814356e77b72fd89ee7e5be9077e1e1585fd20161b04d7d90d32c2a46f37c8bdf42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24449fef41111e082675a623db7cce9c2cd3ddcaa5266d9d1cbdd80618ceddb3b20443e04909e9cf27f4998fb00bdb161476;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heea7c5d0f02e28fadf574492b08da15d677bb7096af562daa60a8c092e5163f3c51394fdf56a5a3159fcb244a673200675fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44d0458e02c332afbfbeb49930842ac5fbc18ad6bb796af0c9c7dcf25f07b923d0f25c3327de92c01370a882329452a8a287;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e62cedc868614f419ed6b98577b9dccdebf1b303224a3dc44ed71cbe5e1996053464b8a8e67ceb0e65ff127e9814187dc53;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91018c4e116f710d60cab34216f43a815a8ee52c69111fd2ccd82a18f087d7f71e7d6afd093a282694028456ec3c64785350;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf417ab74fd72b0cab4b420a05ae20487c82cff6e0c8bdef7000b4779067ed013464733dceca1e292074cd59845febfe7ef9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h447bcc60c3693bc83142037e0427d656a9bbdde3068e77c64deb9892aaa30f19ff34b5abb1a326e4b59dbc5fb84a34b48f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9844e17e251b2d264040e577dccade0c82db9df130959b148447d479b2e70c7ed26019dac4e6400b7bc0a96320cc5c42a17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf722015c29a74f479255bc8243419426e8b760b252a92f55599de246afe6f7831f4ce8043ce58a1cc182023d1dbc72d648f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd500e2a83563c1b91d53db32433e554d49c47549b9015ab4fa9c5c5c65b6adf8b2939b935e7b76342a0ea66359a2e6481b11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h579de795c82fe4d6e9849a72ba823df3b526c9e0ecd96f8892cca2bed7b9526cace1f08797100ec252a1776fca6b5bc1a910;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60e258c97d16eb38bad55d535d54288129fb52e8099e51aed11f8ec8cdb89eb4c17dee38a1a80d0aa7f88e000d392119238c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bbf856be4cc377db7556658b52adb94251e0f14c5b9b102a99d358d12102ed81b159d0ff9937d58b110108d15740980905b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaa11cf60a0a762f12599aef6e269a53024ab8bd8ac985c9f3acb44fb9f5f5f5dbeb7d4f0e04029aeba53d0ba3728fd6b62b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60aa65be83c0af46610299407ad4ea6615f908185ea0fa909622fc579e6957ee83f91ee84046ef4e0d07c6203ea487cba9f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f7f735597089b8333bbe65acc10c0738b7545be423ef4f47fd61a5a323a2ad077d30903dfcb624953c8656025ed0a875eaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c3638c4186a93fd728a42b9bdadb3979129bd9a59e55774272da66604a99fea2119b99368576b58140abc0be0f6774a0ffb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h985150875e39e40d666cb28a750465493ee575f51d08a299a573504734ef1f6c1415966446ac1567b80fb978266efc7f7071;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97e61d500f29b4aef9bff5f961374058b7747e75517fdd7ffb922d9f360899b74610b8a99bf645462c23c9e3dbfa536a99fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa34d77a857b04f322e17d2313258bc4ba680d5721bb7e35526c5faaab3875b8cf51eaf59d733a75f8c26140c25aa2748716;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a8534a34dc4d75777d78fef59a9de1467075110cbd3725768bc9abbcb5874424a2ebaa05033a9a7edf095ef72fc8682df48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb3dc2f42c7bb1cfdae1706a8caa0942583950beaf698050f57985d62cdf3b51f6eadb10a5da0c1763fe52afbd2b7d932ec3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bcb93cccf88f0028e7ab5ee02cbc26ed816f0c282356725e34f46de801f46ad6a2ebcd59b624f02d6fb20ebf01ce0a6fc39;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27e74881f0225e3c13fa41ae91a8fbf91ad90c5f433c7558b56ea39c8ce4ff97ff55036500d41b5c9de54f951cc8cb82ba4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h464081ecb327b63bcba0424d4aef90fbe8510a4ffac32238e42000e46e85f6feefa650df7e8cf02f3a9d618ac18d216673ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c8c80afc36c47e7bf2bf2c57247dd8b9a52cd7cbfcf783f20980d73101efdf432e069a353d14569c3280f0944a2b7419cb3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa81cf2613f3db2f5fbebd567583992281b77d6690d98cf0d00aec7a9691e95652a2a5c7d7dc168b4e6008fec76463a6a9b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7eff823f4adc50b3711e67d912979a71b4a9f4f5d7a551fdba40b99b86983d0df396f1a0a6c339f447f1b614ea836ef3853;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8546cf40f2deea283873ef8bf3357e1be3afa56734807f31a6fe67e00d2b9052a5a15abbf54892b3e10eec20d08eb43abcb6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf03f12af5c624008d4075493168a6eca3d2e813ebe88e72c33695abb8f5ccc2219b5ef28a047e5ce46f889f2bd9e31fe5560;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbeec2eadaf71b744d5b9b61e620e7ae048b35c3244a10a7e206680577d011002cae9ca1d1b012c9edfc48efc031dcf556776;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19c7f27011e72933eaca3f94f743b87701cc4eee400c207f15ba95364046cc5f74f7b40d21db35e04b62fd626008d3bdeb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae024ac0034c4f84993705d0604146cd6dd6dca7257428f6c560442e9ebc5b9082eb2aa5fa67eebe6cd313cc49c1a586d1dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52ff3d32356632ddf59eec9af422b79fbc2ecb47b83a64c1afbeeb87bd63583319f16efc7a876f0222cfa11d61a4df941b1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf151e38c95d37c82e28e28d6812b568896b4c120a79bcd82dffe434747063d76f1b63d626db52002154bfe4276524a84ca3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a4ea74340d695936d651ee1c93d98d38275be29eda8f9da5d2cfb8ac724f295d47703461236834fde038dabb25ce74c8f57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1b4421df28556cb954c062a48b9483d2048da5bb3ac5acee2b10478047cb49812cebc56832b575e6c44dcbdecd53cb3d06c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb07a426456b56351ea4ee1e0ff4d1edf02fe33029eb14715cbc4be750e99a4c8b235a0c38ae4267434a4155409484cdbd4eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dffa8f0e41cbef7ac3d92d6f3c21065d0a7495003febe380bba756810ed7ec5282172c836fbee483942bc0c8a56006d74c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he746cfe70fa183af647ee5c24d604746ba3af611c6b8ad4cc1d96f5db81fb0215bdb8259c979a70bc41737373a28e6552887;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68e7d0593091629e20d4aec819d55cf439756ce7451c620df90bd3fa95c4eb9cc0138c5ee8bc395879fbcfb70dc8489cf400;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he830dbf808fa2f7a4f1108922198c45dc3cd2324694f5a069b8a8aab187f36fc986d98dc92bc376d944639698daa9a4980b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h588b2b2e37d577c7120860decfba0e16d16970124db94b4487044cd9cff4a97b78377cb3f54d81b7de4c7de9cd055b277bed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3173bcbd73481e4b5013941a1edd613ed025dfb8bc8383d70d12ec0943dcde31cccccd68d46d879576f894a3b4f403f4e7cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e36c60c48d43874fda8fc9510eca202a2227f085f5224fae44082c8d2abc531618f67fb71417db1720f6ec04496f995d90b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1df481c810136050913614c242ced82f60b2fe4816fc72145141aa2916b230a2498050a384a44d3cad3ac72732740d8b2555;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6be21705493af293893c894798586109626966111ab14f3b5e5901183df9e82053d58a67993542231b102505c50a1016771;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1252d8695309200619d051957655f2b1a2705e07973b78c726c6b253bfc0eb0c8449d431875dd69b37e1e7bf2f051a231000;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbab39add907a487cafd07b3e86fd988e1606219b67a61fe6c3480f078921f9c5d60e226b70e31331495de8d12bbd52774de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19eababf5d6e9cf84db8fa577672bd630240f4f18af2ca3c7d8770500c82a63c6c05961bbc695381fc95f1f50f235e8a7c4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24fa00c30b4c43da1b8b91b7640d8482b7d84f998e36d933e97f8d0092ad493057791a937d10c20131cb36afef015f4d2865;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9488b99050e9d114338822b9aadfbd684fbd0269f76beff94bf42df7aa4ab92479b25b3c1c3055e6b7a27474e867ed457df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebfe80de86cb5339ea19077f63e572ebbfd63b527ea01aab479a5acdc07fea929276cadb7521739415658a5454d19115ef12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6ed190401d2397faad289c357f3793c57ce8f67aaab82801d6272d0f86f39be99e8c878bd4ce7115f2530309b7e44eb8e14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4767d80dcbff482cb91b852cb124608ed717824f7d4914e83819453abf6626abd5acd6d93165ab49700472c2441264fda9f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f8fddd06a081176d3ba1c8b237831bc3336996706fd3ce89258f0b32de171fbf0c86b00c4ce31949e0a8d0debe405d5d77e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f066bd1645aa20941a138b6e59e3719a7d2a0bd06f2da8717a00042ea2e1393b835193aa549874a48969b2d9c3a5f60fdcf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h159b4d4f3b8c656d73f4c0dcf91ea4d244acc32166133cda2f6282f32dc4fe06f0e1bb3cb13817f42a5153afbb38b2af4299;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bcf2eb0d9e242b8a4103f5bcf935a64fd4423c769bf2d09e1eccfe34b38ae0da6610436e862d74d6f50b1876cfda1176775;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf439fc16667e39791d10f8bc744f2b3cf87fe4503697dd87c64b8f183e99ae8900de59d0f767b27e1fc2ef4a063ce82f66e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8ae0ff3a02c05538e9ca56091e947e2935d59504a4deec74b65dbc30c701fdcb7081d4d89fa7faeefef2cdf4f2f2812834b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13507596bfffff78960376876313c89366cd5d80fde78aa001e35aebf87b187c9bcfab58abd61f123d6bf1df66bdc37b4ca7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83b7d39e0ed64b51c3e6b25f17f0188f58750b2d780f0b21666bbca4f6eca2903f18ed70251ebd8d809f2ac298377cf9dc97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc36217a0985aa9cb014f09771880b5cc6879a013c09492a8f6fe7db35a6198e654bda052e4f002e0cb4835d7ba488157ecf2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0ebb3fbc57e6c4708f887ec2238254195e53cfa357dac775d2764fcf8a0d99006fa39c2f28bbe64240e0ee5531baa1b2aaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf85a77aeb8aaf6371add49aa031774505b7ab75c83f8eb9307aa6d68feec0032667032028e74d6ac72d8eac299a1cc3d537;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a6f26bfd37aa1e61e841958025b03a082ed9b4c9117a0c8a7f219bba6bf48f8221b81ae5e723dbbfdbf61160ecece5a9c76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7587374d2b95ded96e7118dc67d3b394b2f9a36f86e3f914d8a2682dd73ebcd1d15a179c4b529fa4eebc8b7c5047873eea8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3332e3d837f692779b5c56063aba690be438f2fe0a89127983fbf59a3363b6eb5d57bf2016ef43ee593d6c85cfd81332bf1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he031b7485c606f5c9913e1ffefd715253f4f73b380f8e3f052de665687227820048df6333058ac9147e3a556d6da8abaf17d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1bdd4f6f593db1b087f8f0076d541c71fba5dcad65537aee13a4c242132bdaf7db8a244aaab514f93437345393117c1de8c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeda7bd2019abe4f68943c12c0ed66fe4e34fc4b48c5fad65b4f4357b4aabb9804d923eeffdae9b19c864eb28a8ed40301be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e3ece84716aa85b020def670d3ebfe5cdd5eb054e5e29957f15b24a95de344fd591bf87638bf2e22caf91682a7ec908d065;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb28d8716bd63be09efb06e0b86c1d6749f25e963a664624c3e4abbab73c5808070a901e179144ac65247d18314ca41006068;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94b9b4789dd2bce5e1e062cd9d2bde295bcd69e6b27d041169eb4b0a779c047ae928824da9e9650aca5b578eac7a91fa12a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9f11d7d64cade3827e281bf8c6c13e1239510e2b1cfeb1bff4b425ee4915ad7e2daf6b0dfcb7c0fdc72889360fe21d8f40a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25a68b1debc7ead46205e4dc1d0c33bb8e8218b1d055751151bf4f474482e31a5627a48e2506f9adc72544ca279aef0956b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47944582909e061c4ec7f3786a7510a92276b24b8c16440f03e5d639b1a905a57b8116f4966b9cb10e04011a116f5818fae2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha337a1051eaaceb283e2b6a762f73aa0b67845297894b4f8b0fe3e501a59df5265420bb801fb2e6f6a2a6f68e8fdb78b11ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfe36542acbc7f0dd013aadf5880d77506d3eae1a9b850ba004daa8580abb54cfbf837a7ec5b54da7da6c3de295e6cc0032;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c81634d4e15ed7c319c4f9e56f689437d485c1bd0a79f7387cbb447b1030c1bd9787841b9b60346a87588cbfd0a6d03fbe2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8c6f32235a74786ed6d2b835dd12a71b0a2d52a6c932adb4b83595f785faf718756135149d0a148f4925746e96a4e3f7361;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h543bf25c17969f1a41f7ccb1c1ad81a0c66bd65dfcd7cee01a85b796c624b273a79eb10cc2326b7739ee9eb1424c6110fec7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h563414c65d4d264106df3e787d6d5c5e5c6972bea33ea67d37425827cc746b89a0a537ef3a00bb47df80719e71f474baed71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6a41e0c7c86979436f2edaf9e5604d4ad937db73a84baee09f41aaeade50854c9ee48849f499b1defec869569c1fdd94caf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h536144f7dae688b513fbc9ef32ddb9f5ad435f731c29bed761eeed39758f3ae948a0c5271b82754d4762882a232dceedf9e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1538c79564114c5b8387c4d31ad8b0062e7a49a38b5f9e5725244bf69f022c7210de8a2b45c563ba28e8e260233d8e2bf1a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2522eb3bf374fd26ab0606ef51f6e048f1cee3b5ed2059c132e95cfe67ccc0f02abc8130a7bfab666fa0c76617bdaddb319b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dc9c0566957c1a7f874379334fe43c8be9f2df5b3e1576bd1866c0ec8041156e4a4dcd13296fa003cf6e00fe110b52de939;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1ea6839d64584680b8f0d9e9ddf426ad1cb671f88ffcb52993184e0cfc522cebadc21004d07e65009e69819c884b370489b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21633c8d378f16266f4708194cb6208bd35abe1df2c336e221f6729be950020bdc550f1ee6f3f41742cbfcad6e850693afaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61e18a97e11804b1d3181d54ec7cc33c4f6333cca43cc79ec829ae7c3d61d4fd406fb2397b5b369aa8f1edb059660c0a4ee4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71f98fc4c19d294ae1740102d6b6162d9c15a0cc98e928be66ef4d17b185388ac197df1a68acd757d15724aef0e553919c1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b94eb2f7b0bf28d73042b9e57a11584cde15fa066ab4a8c590d21765d2ff325d984994d721dd474ba08cc9b0bb17af7a0cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb13160a77dc458932da489b425cf183154a8754c4add4aa08e7985862118a054ec7a0e719a46b73f8a5ddafb4cc2d1ef1e82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9c63b53c4e7ea2aeb5a2b121bb6a2b3867a91f26ed274f8de333d74bf9ac3930d6accc84d41fd8c47d983410a62720b631c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e3eeb52e4885594cf8191e2060ce0023141806ea493e27f8c724b67ceb8ab337069c07dfa3871a2b94e657fb6b482bcb801;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf25be312211187864c50898cf9b401ef1104a1860e60fa413d77e4bfd2bbaa56943c74efa9518ac6322931b86a1b48c334b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29fc44fdf5925e025ba89c34bd61def54e49c012b4e6443a183b1263fab106c641b096aef2cafa81c155cc00a1d4c4e92783;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h953def1dc2de49f8f0866f9985a22935afc4286f3e4c693b4c9b7a77467c6fb46520ac0fa795e64bac7e8d966850be1b269f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c2a0074448ea2791a83f28da34e8d1b45b2ff978983d24cbed200d6527470374a695a38e1d98c33e61f9d4c52c46498febb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9d5b25f6ee6792cd04ce48e37107edc4bd2a46f6dd6638d1c50cc74d7630e782d1caa68bd4f5c3f7c773fc1c5fe00a75b85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaca8963244fd3b0cafce97600b31f92b49c8ffaf76fae6e1cee972e3ee82711c7df30c3c78c67da99236e9049c32e7bad43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d553353a8e7a875fac66664483e3eefccfe8a0267146f4f38c5ee7737095b4d86dcb4fbde383a1cc783a48535d5f431ed28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he661783c48d5e4b8fdf3af67db47b0cd60b8fa55a38a662068a59f905260c73f5f4f8b30a5b8322348df93d199567f677941;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h767ef9a39b9d4cb6f6f05b89384237bce059ffaa159d01d8887d705210a4bb1b0561be3157c6957f841a0b7677238ea3428;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h898e7c5405e51dc6e6ada02b789f399d68d6ee80cfc1357dbf6d5d0ee8dd1cde4b478f402cf21c8dd659d2c478fe8a7f302;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a7a793fa25b4fed22338b7520ad16b3c4841c744dffe9022ecc7144dd962d75cde1892eb5831b50f25132d565a4c8532741;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d6cd9a8d80ce37a5762b84249e76107eb4c0c7fd2a6da7e332d3974e391507df761df2ce20be1b898140306025dd90061b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb57480ce9b682dd13897763ecc35a9deecddd1120ffe17d925bf83829ec1ee7c589f3d94410da57a91f52d384355b7053759;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dfbfe5dc256ed1884ffe6acc5a99573b661be4e8cd2c3560d8586e1abc04b1b079a844b3a582053e3b5b98b58c0bb0711c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h537bf1cd2afeb479a969d578ef5e0997e38c4ef9f727823e343b3b9d7ab74daac19f459994b0eaed190b4061bb3f9b1d0d20;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55bcc347b3d6596769729673e5e2962459e856d9cb710e83a9631d1714235d344ab482066c8c01bf25f581e5133fbda526c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2faae5b1251cc28fee40c657b6701e4c204b470f4c544ff784df479c4e67fe153697f3360376c6b9469dded96484cabc91d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h650a5c9fa4ebc5860be802580d18b2b7e6542dcd0c2be044a5742989dff9eca35b1e327424044856d013e34caa1945a12bd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a3578f308e2c97a899e0660bba6d1efb78df5f4040d699ef27127e83ea078df39fdf3c8f7ca1d7e7b49a89a21321493bc4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc4d2fd314a47138a6692d617d25091e7453c0e0b77df8863d03ffc82627fa5e57dd2bf6e103e785b222cff6bf97f5c7b7f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9f65545b811e384827cba5a7810d6c0cc71399ddc49ed290218dcd329451abca20a327ccff356127edc82dcd667ec09a40d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e58bc5a5303bb79220cd6e9ececed42fe0b09a166a9cabb874def1f71322f50ddfecc7b6221192b82100d4013889b32bbef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53b1a8642c77b61b5a05d95a7e5aedfe9d2df176b5d862f943cdb508f55590fe62ebd64b8a52d35b18f2af3949e1f2770ba9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d9162cfa8c6eac58373542eea5bff441ced373e2dbba1aa52c828d921d580f8504173154851f13d4e4263a7cab868be0a31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h535795af5e66b2e643337cc7a6f49a3e868d7c281d62c92775430400d06ab3d1e51cac556b7f89647c27671058388dd28d52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbad28e85af59cbde84b815f5b4b00c8298a2f74b5b8fb36a6f3350929ca6452611ceca6130e0bca46b07b75b66c83437e4a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3be5935e84c158cd03b11230f296b9fc0d75dc5f86ce2e39716eb3831d6ae42b26e7065d81fbcbce243da58c45df6490ab73;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd9d99a2f8e7256c6de39d5ed8b2736a783fb856a2bd7b1ab99ce08de4ff38e357e1f0b06df199ddb863478c891273cf1fc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac0a975c44bebc27269cf4cc0d5620d0f55d0b501d73d4dd23e4730764762793b83587651b104c30d83bd27789972d4fa528;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h324f399ec4a5081f3bda5c89928d2283482136bbe80cda18cfe6f0179306d0e323151e69b65c0ad992a08274d939d346703a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he338bdb7a63e4ecac45863022a5929cce72f3bc0f5084ef5893d86ffa98db6c4749d426e1fe6f172b6dd74739738dcc27e39;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae380ef58f1bfcd382a3ba1628c64d17fc5488a67d2bf53ebbdf8d82c0a39e2388df6af74774b1019e958058f2394a112c82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76699b3954e9f8411bf05075f1c0d55f47aaaf04b8d29286550b4e5ce7dccbbfa4900d81fb4ac7fbd1575019fbf2a868dfb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b0af3aded6b9a9c06313972741702e9aaf7d4fdc3645cc16e8d84c4921edcd871e0c43ab305e9d839c4e43b31d3b72d2cac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h460dd29d3d5721bd674c2224e6a206b3ae6c0f75479de2242dee1462a64f0b82d7c4af2351c782578252beb38cf3e2a0dd66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69a2429e0a4e09c3c853b520581e77d284153847e38a46fd861264534157f0115508f79d55882c43879cf58b155f99c71f33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf91c65ddf85a0ded9f08ef60e1e83186becbb75e1d970cbf26781e212bc5d30155bb034bb98219fd83b34f7cc9c022ee17e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75b24be348a714f8a525b96b4a31ebcd7204a3d341ce97fd94633118e9b38954cd662a4c42c1d1c52c2405e36ad68b7e7a5c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5403e7446be9ddeddc72d27e9121ef9d7ae5825b92e7453124fa11fbe37a91edda410adb63cb0e2f9858270aed6fe65f1feb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd264cf9cb4465873e6046ebeb99dda8fe976220b72198ae63ffa9fa9cd51f3651ba22082abf0870c7178b3863c655a1c8465;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf64f7706e7f2d7196ea999f46619ca1f062b768ef61110bd1007f96994d24a42b312ee90daf0d81b3df322b4cfcf566a945c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7f4dfb5182d0c8ae5b77bd49ee2958b0e26bb2320650512fe80d328d64db8738c08c77ab3cb00f5e2a613eb5503a620a7f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h456414289610cc39165fa29667d706af12695a1e1db5d47ccdd610927dff041a250b9471b870598fd79e36e9086a152ee5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe7fd2e3066694caa2de217aac26b5bf4f554949b45a7309e414afd7e01f112e3d6bfc4eec1860056574832b2cd29a528502;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58eca1ce2a29f14ce7aaf84ecc3c37ea3ac79514d18a8d0ec61caa21aa30fffa44b7137a7bc830b2ff80b1eea55a7c03ba83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd26401844a9fe1853de42e92288f16bba2742f74f393f9e8ff9598461bf3180c72c5c7b962a64686aae30d796fbc926a218;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7d62588ca2a7a8552294af7bd71ecc25816a90c87cc182284ab959c1b5980831c4e80a7db2072f395280ccdff21b1b10a3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b332c717be5e2ce4e4fe52aa69c42e6afed68d56ee8e615e5475dca45c97e952c0182678330927556300c68d5087a78b030;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2be3494c1550e8b8c7c684eeeb92fd8079674718b9aa8bd144f6e013b5de6ea38edfbff230f66b4ea65ad407728dc33e624;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fcb80429524c431cab13e8c2e7fdfeceae2f1797c5b290881949dc4478e681edc4ca08d9612d09690712b24193fe9459c1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfc6729fb808f8bff8e71ba3f1eb159a9f41faa7c9441f49bfb9d980e32d93df54df36647a3fb710529aa4c940595bc9ffdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b7020bd73eea62f71e3b26cc4691299bad2a6785526dc083f15e5bd096f8e9dbd55a46b73f69b5f2ec6c21c2fbc8df428c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haffa7f95e4dff52c8c34039fe0684e546283cd5077a5ed29e65ae03ef50fb4c685a8c5358b37cc8df1f577d55080b0e5955;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7112973eacca7882f0d6fa509178296f8a06085700fea8a37c0840ec2309529096242ef045a0e9e938adf513e826c0f01baa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98b3e6473849568e7c2c0d98e48829f608fe5d3c4b5dfcbb5664a123c66a2a507924bef0753daa2cb39dc153c079fa5c834a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7087fbb752b3db680c317d09635381e4c9d9a00ee981b4f71be7853375b9715bbc45d2d78bf72ad2770dee95815cdc1553df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18d35c523f77412b197411c93cd0fc31ab09144540cbb666397f6c258b804682af8f5d24de9d6179ff4ffd892b1543b88452;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bd7eb87020cac2cd4efa4b26b61230b1e3f0329da7031b98eb8c6a503ba0b3738d1757348164107ae4b861cb38e67d6e7d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he638b2c7a9814ee74d36ddf77509b59a4a5cd4773e96ae019230600332ab31ebe17dc233d68b312e76bf7dbfb7478af56c0e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf271ad879ad4a1c374a8ec3fcf4feea7ba51365c675cdbb898ed051e8e9a2a3fa24874af3bd5f98be090686498e20da3790c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90c1512d1b38f2d6e315a2f06f70b3418005cd6cfcd96549240557181c237f2479aecac2aaaa725456138a58a5da689df8d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he714e8c266235044a1ae4636f11c1dc2bdf804ce7aa7e2dcc0cfa797d50e943d1fde1b4e29dff9510ff7e124ec63213f3bf2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d3f1e2e33ef6e5a705360bc991238735c6d033df4d93657eaebc63f7d0890632c7648da2b4950b40925110c9db53e677172;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42c0d45f7ae7fd7e90079a851e174f36cac94b601a732bb16c01ece9d7068c426b7e542febac13b222ebc3b206d58df7d832;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h652cb69ae8e16957cdc86174bfd774a588c1e25e81396705db42368a2582f0443809fb5c79420828e2ff9af990c1b76ad539;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h574389f8a6199438f050a795feccf6682a03f9dfe53533a7aefa6c9772c0c75d99aecbe0f95195aea2da8880ac07579aac6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0455161fbb92f5dacfb0415ab75d38ee41db3f2aac34c74c5becf87f706bcf1b3e16a99fa723196799737003625c6787c10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5bafab3c3d67111f357462dc8728d357f88af67964fd4e3ab360abb1a47108961f7d7eb594c9265234d88c465b11d2f9ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d57f26cea1446b96129a63db655225db320b1460d1b787a2244c5c4e91025f8a51a7542856cd6b5f5af9bdd018707659692;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1ade99470e84ccd3cb4c487716c2da0dbc85fcc0cb0c437fb8596e4b50f5d4f225c7cecb05a30e43092fda2b28cfde96aaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42ad7a86d09e9ac27a25f1c3579708bc5aa0a30c722c55c5533bafdc58c8082a7b5a17e308a7966041951e73e1e1af38fb51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h844492af1b6dd5e756af237a613bd1ebe1896521827f85c1b3ec1b869ab18be0c428be76b21ff5f6ccc8cfc4a251066961e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1c609d29b145565cfd6d3c005d48079e25a88a71ee340d1aee10140d6f825fe9dd57c6301ddeaae310470782ddef716f865;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d4239b8e5bb7e972550e3d2ec3866076bd9ca3d7a65606da1a22c4086834b2e2c3b6de5151b4aea6511f304a27cee258144;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e5f78be472433a0fb5d01c236cb4b4cbba2becc77deccbc6161399c115fde2dd06ab86cbfe843fd2827012a533015d8f10e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hced0c6b2e237ee8e957858f7679594035fb7ad37535eb8e3ae2b1ab41960604a3842c13ba58ca7036ba4e192c629ee55eb4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83bf15c3112a453298c48c79d1d24df6b4b1268f702824182e481777dd41df4539d058a40d4dae51d55fff401af9c32c5ef5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53d59b3159b1fe7eb9c5a2056ff3e8a06b10d3f6840ac02cde86490ec9ab871caac28cc92e9f4da6ce8d95ae06c75b41864a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6c0ad38958017fb63dfc910bf0c263af4505fa7d020ef5506435278d611e803b76a7186230c92b21f571ca30471d92da5fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56aae2490d548314e8e1431fe3c9944d2ffd831886e9c9672f669a32e919d6b67369c886b10ec444127b9b6aafdfa396b5e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a2b2984be53fa4bc6f7bc173ca8ac0fe49135fae245b9ab4764f27a3816fe2133b277482265515e2b347bb4ce4685cbd8d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdf43df1642ed1afa136ee214952c42238efdfcfc76f1ef06213355ebaefa25ce25b2af8a880ca13a9bfca795cf0424410d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h323249709d7ccd40f9b2249660566ffea510173bdcd5eabd55c03bc974d1c02e794e96f2619720b3595ef7b614d314da95b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0ee5a161c7261d2e7f94c0b0245d5089035da6bec634d2a62ba4e2ec5b3aadecab744e7329dbaa90e0655daf744dc05c5c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e74e98805f5a77787b91df1981538c0effb48ab1ad335694b7df30d3033bd9bf265158b5fafba7d6f90cbf7f80bba86b1d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a4d962978388eb17449422385d24f7d0d02539817c82e31e8741c079026acaab7c6e1b9ce8f76931d0df3e088cbe2794034;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3e42b67dd709b99d610bda01dead4dbbe4f3721b4a18b540f6e20b02748b620bfbf6a54679ecbd53675ab5c7d94eaac82ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72ba4417782c1c450149e3b07ef219c2e4dde3316083942d1d6d2577388fc75908ff3bba64d102fa71597f563f9826a6dbdb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha69a812f5fbc5ba71f87d3a8931f84b30dcc8c763182a993f1373fb1e43bcbf138a7cafb800b757da01266100c8e6781662;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf374297cbbaa4aa8d269cb2cd568762340976d4f3fb67dc1eef3d92565d46c19aacf88e6e0a5ed4d39f2166c0b0be6960882;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h848bb63fc33afeb4837a97ea472aa1e78bb410afe6e3b471a67b6819225a3b5fb1294613bb1268660ac2b0c1dfc591fce2ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h952f8817b7a8fc3d1a0f7f25aca78e8c1d7704574d496f384143511f63024c2b19e0f4d877a658c65f00132c828a9eb7376a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7de1bafd52245e899c45b1a8add41f623255a748555802bff1b1f1fc715a15e86ce8d36cb3f83e8db412251f5650d9ef0ba8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9572b151e362de84ef49728a4aa3c0c7d882d4ee9ab64ec64a2e350b89c7e982338dc3a5daedcd928018cd443eca5d04da11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a6cb2ea546ec35a3863e841ebf06edcc616e858e343425700eebf2b3e8acd55b3422d669741916a169a27507be03ce0b0da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb22417bdbe98518c8052ce4e675e151437356e5eec25eceb17cca4b9382d7ba48c09d6716ef0eefb29bf864e48b2ca198f74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89a1495cca97a184d5ed7f2bebcc5cd7d7407f6becfb4c6ce20358d095cb0c968baa8d8d6d4fd9fdd7d259ef740ab49f2133;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3eaec474913520914ef10b998e4efb8c1618dfb3a9b658d52dd4abd5ae194c4f9052fd33c50255575c4e6cdad18cf73206c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7341521e3e1125356f6e70abba876573113e598d1de764d35feec82ac2119c8fdc27879900d3eaa7590d7adade86d5c9f9cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59eb133305089327831e47ee54f67ecc74a4f4abbccdd09026b54fe1aca9a4d99e67a85e9ee18c18d0330f35bfa1bf506e4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9aa9d2c067ad54d2d5442eb34830aa76384aff0f6d4491684e0a6a69c8fb87dae4989c2fd9f3ba4b9e0e72bfb2ff1d029d9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h867142eedd0629f9fec2fa1f36fde25302ba52c30243beb51178b742d1c76c1ccf605772e6d9faa99544e29ae0a360f9d44b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8df6426b701c5c087c76844805514c1499c21e921c2e0a8a12de63420926614820a702e91f798eaf88b42a3a7e41d0776b1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb99e9d60f6b2f092c0219615bfa6347e70037228ab50191b907ecc80908d2e287d036954414cebca8583e692431030caa94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd72cdcf8fe2ae7f41d138315cfc496583e4fb3472baca29fc70f78a129b643333cc63947fa9b8e5108eb422a526bb4b64026;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65a55b760502181e458ff7b3ea77fa8f8ce85092c336fa4a73ac78c375624f7230398303595883f9c82141270ab091836bfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dc3b13ca22ae01d981a94278a1f69e8ca83749a4709f1ee5f7a8ca1a00f7b3a180cb49e107d50ffb88e08934e63c6ab2d7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h188dc1c97b371e97e1281c6b0981dbc16d0cfbf712f4258f6d14a461c283f6fe0c7513668ee8bad5f3b1f2866e2da046b17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h818b92538ffab19d24d47dc3ae1058249b680f7576874f2a42583f9ef7d36187a71573fbfd13ada1702ba76d8f76543566ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bbe189cc74c8fd8cb900e684cc56cf68bbad66984aaaa09db8da3781997fd8fd487e050b822b37611c7d018b4acdfad098f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc1ae76337b75cf7865741a45f09402a173f090fe308011d55857d8d0f87d00ea43b177c7be240e62d96427a1c85717fafb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bf06e4f40a0077acaa2e5e81d3287a6a9200a6b23d5705db1c8f0a55cc2ed11570d556270c3b1511fea4d6962619f147010;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb774b9ef914c2c5596cfdc59ff3e84e243f252a8cf01ff2365103091095db775c5ec8cfbe890893c2d40bd95faba267c64b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cd4122c86fb64dfd9fd075c5813fdae573554f3deb883e42ad1a106c909fa423a6b03aef3c9f43855fb431a989fdbfff357;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d2210e3b9fb56cd021e9750a3d200610d8f6ceaf3bcb77daad366c59027b9c15d925301ea5937afaa1c573e7acaabc37daa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e123ba2dbdea819f16d164dd316ba21aa105824aabf9b02c7539df24ea74293ad0e29220c6297e32455628c17bc53bf0566;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1a1f0f71a52d07b0773273785618821ddabf3bc01c8f3266822451d462e4335a2a3de36b4fab5cd99efd3cfc817305619e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29e4479c1998a2c4da50d355d00e795763f8e0ce05863fc57ef4293890a2a357a19732d06e27942ebfa2f2e8ca02119162e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ef8c26d3751dc766cdae2541369dd516928501ac4830631e11a81ff67f11c331f80e2196fa798b1d2e29db789b8eeeffaac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd2e4ff11c3b8ce2bb76f70116e924f4314bfe5960014d11acb709ba51ef67498a5323cd6338cc19cb8a0b44dff75e29d43c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3837759a664efba70eaa0419cc2a85eff2bb4ffc1adcfb9c9a512ac201b79407d962d18d783c4943a9b90b1b3b010753397d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b3e448883d718ed883a4d95c0f3626021e08c3b4ce411b049cebaa2923a3bbb8177e914370b66df20c1b794d04bb18a28ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a078a96467afeca389964b91dcbeb65f0dee6f54ba39461f2a36669c835b959f9326c236622d2fb76a3806994ab652b2bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf081db898d0bfbe1d305dd6bcbb5310cd57ee296c0a6b55a5f8a2beff915174a0e26e8bc932ed012455399c343b595b557b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h788fa35df2f2a0e1033897e45e23afa8bd953ee537c1ad4beac41cff261304e05f74483d368c7f1df40a07f21c9b7da940bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf606f1d9ca8f2712d6cc8264b8dcd677b3864be3e5c0541186382f5a8686d74a04e859964a8ddd046f7db0d33b36679c9432;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3046377b371f9a9d2b0f6d3682f9c821fea1fef4888abbe07237cd87310ddf2592353fa761fd212b89260d35fcd8dee0dfc4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b411a2566ff2a8a98687d3a7ec69ff4c02b5c8a125f265c2337a0b4ffba917d6143bd6bc90aa96f7b8fb0b78f3fd36cbe6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e7958c6b86ca0679fbbd439a72b21ffb8623e2783904ac155f961d380fdcbc169306e08283ce39e699f712f7974619a6cfd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0f681d96ab0228c93ef44ef2cdbe815ed646796c90a8894b14047e992d5ae2db18a84208cb06d360eadd44c077c0a564fc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bbbaaa4c4ffae8ef53e6a5058557ea84c758fbf1d674256e9cd25700f9b99a4dbac81b479cb0e2c4e605f6658ffb06d8214;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c93c3e720ecfa4c070f38b2ddfb34891a995f38fa38fabef19e3bc3bd68c7d33c318045ce0426889f7359bf33bec128decb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd692504164a3d71d3781154f23f83c95b515053000ee27204ddc77b6d2927a2826ba8b220a02a4ad472ffe2aba9a099606be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e12dc4217af55947da539380de970cf1a79c61852d9b36785747fe6f2e4cfc696102291df5c640e4ca65569f7090107ae21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aa7490fde7b90a91cf626b8291bb3541aa1f477df3a8f5b2b047cc12acc2007c0c2c80026aed6e8f7766c2908831772d4fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h277280f58e8a561362dc8c2d6a9af40263e3abafd98ab8bb6e88aef2448859a96e54070c801960dc2c833f34bdf9566175ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a93a64e46cc915618876beb4660cd888e0ea2b64c77500b90c5a0e57bea7f326503acc41902f3fde36e3889ae276f99e083;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3d67143095233d41bf54cf6c0173502b79d4fdccfca28682547b6adaa4bc8724106ec0ad09247b87ee37d6b195fababdb96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cf5368491042cf803671a2cc4926bf53c6e9c1c284cc993c8f26503971f5415691d67f69e44e3c9a409058816033c75cd1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66cc333d12f2aafe9c739f35a4421d56bc542111eb7228c309d6e8ab9706a284e414b40b770565e042aa6a9772c19dba77f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h449fafca26412647e8ed0371a293236dde75014b3aeff6f2062abf7fbfc66fdd059c57130205a9938c67797b41328a325c8a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1af195ec59c6889ddc87d085a6178c0a08643d0898ade9b4bdee0daa5031b744dc3b42eeb374c88befd78ea4052e5fab64b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h112e9b490c6f0bbd23d93b85183353f9e9f7e179b2e81c5cea1291889cc278a7077977f408a9a2e1079de86fd5cbae1e45d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9671207e643552dbea91f2aa08b6ddb81312bac62cefdcb3ce87030da3e0c667a02c0f75adec48b98266b0e4afc788e1590d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90ee2997d4cd96475898a1a0e9dae07847212804abbec542f0dbb1ebec5ddc62e7d0c4fd4b417224c71a78bc157dec1d6567;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72c9a7988bdb9f4bc8244e1a17ca59fc8286cda7e15e98bb39cd5f2a6ef1f1f7aa2c23c7f30a0fc045f7110c6505e4c0c2c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc082fd1e2f3dcdbdd56ba1462050da9324bb47c5fffa6b87b0fbb7944029e403f54688e6794b44f67c37692756c4c3b002fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59d9bd04de62b9e85bfbaa91efa61e0c3838554223cf98e1c542ff43f82dc9fec2092ec42d76fdfed3389a6418a73405f93b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b21a0bbeb1a8877eee1f1dbdf1312da8626a217745f33aa0172572fcd9d88dbf5786c89d551e2cb3c45c5b4fbaa186b8f5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ec78f363f3fef0b6793b0ec2358a32970b232132c6864e4c0d0c6d42398ea8b3d9725b9bb85aacb9d8e462e5c79c39ff385;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4895d3266f6bf0a1d4b74f97c948499c3fea4c7634701ef131366548eec6c35d4e3494d8b353f73d205f5ad40f6629fe1a8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee708785321fd72ae3e020fb3128c76cb370f014e2b13072b1618dc2e6f32f3c8c1c5ff221848ac1ceb6c0c98c602b12205;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9e9e6d270d1cd84084ef3095db42aca004a997dd57a9ff30628d33713c98cc4bf12a44bbc9e03126ebde420f95415f640b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72cef861f4a6299ea58ad7225d777da1a8ddb909bb2040be5571f841c3760e99d7fe0d96ac8b083ff15b71d2b031b9407dd7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5770fb8735d1f4455400289c9d5beefc2b3d6bbcb3d29d29c6f8dd2cb2d55173b6496c83957dabe89c8784563ce44742def;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf45642ef753661ffca896ce7a5d11c87cd5ff2d4a90536d0d1e4f41ecf4d02aa89362d2e036810915f3e21d3d3b161c4c1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80deedb152273a8bedcc753938af9ef78454ac1a929615d2ab6df7afb31bd66bce96c94d4fea3b02f73d97542dcb7527f421;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc2d969606d5cb6096a04a456b582b8222b1d3b0cfc7b11e680a20f1bae2e996a1fbc07ad29ab3500429d45ccce85861bb10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f80d464e777f91a303e10be748620b7f65160299a96b0aa1e85e934071b2b1bb2231723947dfdd2ab8dcb8e24619a65903c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had3b47a41190fdae58f17e12527622903b12a9f2d1e065ece6c7ad760cda349cce584feec9b51320c410014786dc5584ef88;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7af01ea5a901c7077c270879ce10ee6e1b66c2cb7470dea1bfeda72185184836ea9af4a66fcd7ba802f3cda2b8930880ee30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1f2dc5c241e3e96c9ba6c6103beff63e81fe65de644f89aa4f3c6a316c46e3f2a08421941751419ddd611b3f4d13cb1480c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd31c5394bfa6c32a0c92d37b42eab5090daf35b082649d68d32ddc94ee5907f2a5cee3b4c5af9ea60a2c059507c6121ad9c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he85df6f06fa8418d7cc36c8deea53de47fe47e4e687e37732cd9ea51dd07c1b5aecb8e4f87c5e1165ba1e05f0b1ad00187f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1d27bfa29e536d00998179091dffec4e4be17939c734ea01daf54c1f4fa17789a1ef807bbcdd991082b058d2b51ca4ec4a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h937831d4fafb09efc64636abdc4ec5912eead9b1468cd923fb283d0c31fc99fd08d36fd673d0d16b7d06e592ae1cc0516c26;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3789f3aa5647f45310f16fa6856e4181335acf5d1cbadb1406ff8e080736d4a9e0ad4c2756a783860836d17351c62594ccc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc85b3c2852b418c416aa59f63c302b4e5a502f9917fecba04410596af428fbd4f66f6a20917f26757931768d8199681f189;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0890e8a61627db06b3ae4e84631fb9acf761414ed1c7e7c4aa9faf6052377ae0901ac41df1cc67b815e34147920db1e2af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5c4470906a76d68ba9de6608aeb794b457b64d19aa98b4476a96834528894ce6f3259152478fa47f4f608c8fb5ef3f0e197;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb284d9812a54e68bd8cfdf7a0fe4e02588048c545923c177c665f90a5172853432686e4202f17547f584450ff1e46b5ad5a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82c067d9c9eb4f5928f5a019cf28a10fb0f8d7b79c76b49793dc928d8be5506b99ec08f60debbb02aaf7ab400409d3ca56a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4aca0da912b710d0b38739eed7c9648f6e6a4c1ef3769d97c9f9d621ffef2eabc2c2902d578db31688caceb50dbd76b3719;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3bc96efdcb7c8026535fb5e94f504459fc9bc1eb46966e0a043bc091fd3100df091d6d246cd57f8f641a8dd26ef683fd3e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5d6088e532b309daee48be424cd1d7d11dc9aa2639f5c8a1c52c487f51bad452f78aa50d19dd2f0f31bddb3f1b1dcd5fefb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38cd12d009598964f6ce5b0bc4164d07aef2c0cba89f264bd374ba5ed123e8ee6a8dd379c9ed88e874c80cd6ca119d376d07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h945bc5996ea8f3351af6a461c5f0ab5c9d2aad8a2ccf19f0076b5cf6e3991e35f9207748d6721152a808a096ef392232a204;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2df05760fd79b8a2a86922dc5b67f47add323488e26c7c39b6a2a9058525c9946b20c3cfcd9226ebd02b7134b627c9e9e60c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e239b857279d8f8609bc225327e6f0550d3d6071b6ef1cc6702bcf09cdf33c44ea5d23b3247067deef16969902e08922593;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5796d8d2a45b89b09e1c09fb5fec3ddd5c29ce114cf544adb68870f16a503c339a0d43f90648c3f36c917f956579269dfc6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbdf3c7fb4a5ae360ee5a196392859de7823d19078f2ccf500f902d4634289936c1b73c837aa190564f56afd01719d177056;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd14eee375be2802f8df0e6c639231a87fbf64c85ed6c0ff3d251c8b0d0c8d3224a8e92bebaac1152d2d1384611ec86a3ad89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ef62daea7056cad44d4d517532c6c459ccd9d45705c90c1620092c58b75bce04e8039e493eb3643124d4faa1dfc91bd5e45;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fd0d7d98050c21b9d1581b794ad9b22d011939273a857422c912dcc5ccbd682cf6bd3da13f8fabc7834762f9b44d6c6218c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7931e9da9b6442ee0f3269197523a17964c4f2a08a375b18b7ce641cfe354fa9341d8786cb05593c1536ef8ffa2a300a2368;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7dbc7da2abc69f231ec250a9c0d0ba99d1e9696c0bb45e28de68bad9b8253b836f9365452d7afa48c00b178141a73cc06a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f8e33fa27c8e8f4a65835b90e206428a5b1159ad12555200e16536d5c1b565c1129f0f49f3a9161fab5812ca861022163e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45b79e762555321b633e583353c98540713aac40302a74d62252c2775de565ac4cd276e2cad70e0c960a79f7bc8dd37c5c12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd001f49743f13c588279667d5d412615f8369d86435003788b9afca894a66d0a3cf98b11f55c7462ea936bc645a34df52af3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11bc5be398cc5f79443de6d37c11461418f016f32f18a611f07467cbcf897e23ec2f78a44d40031bb49c52ab14a224915da6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hada8a4b7e447adadd18d3983b4e3acd0e1fd0b45b69ac525689d3e1b4b082c0bbdaa25872e9ae7d78fd138ba8b51c5846865;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e1de93fae8da538d230ad449fcdbf51245e010bf09d0c729bb1332b742bbc2126f7c9a6c1bedecb84e9f78bb60488be3169;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ff640c77076c6ba1b2516fdd145612e84c486d621e28055b227b2444220e7525558ac621875262243b5c13dff5198a769d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dab0561ec8d6c4d30d1ba2412d3467a3cc8fde5931153e175d04d9c9c1969b65b33de368c8f48ee7005924c44631ff16de3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aec6ceb26ba60ba1d825c3e9c272ae8882ad1c01ca9583e5d982558a81fd45525eb9155c5a7e526905bc32d79c347e01f74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3d91eceb697cb66a6d1c22cffd91ec56583239f6073ea2e8151bb70f2c5aea6c93772f11c65bf3501d8e5fc235b49e61d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca09bea23602ca09484bb40289b59d489efe7f0039aa6569aee39db973c48fa40388c4494d4dbfd70efb46868e953f18ce93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9de7062684fb8a415a9d206165422df5f5d5c9142a472b13f65cd2922eaf36e1057ea7f08b071007a7fb1e9ae92103a1eba9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0599b3ab1f5f523775f345d4ce4b23586841da630c8aa3687c2abfd4baf69ef865031b54e071455c666bd3322c1b1b3d8ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29215a676f78c454cc42eff16a6422411bf560aefb5294fbb870ec0043ece4a3835484037acbe7da639db45f7ee8e7f691c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65afca4b849de4cb88d472477140da2a2617bcd983649af70d1e6345caea7c76dfe6b4651a9075e37a591598cfd967b6a08d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfef00dfca19276e0f20c6c8e7ba89cc42581811a471f126d9612ea9aabbbac08f22eea6ffa48b77f8428a2b0bc277248e37c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5466f320502b53940ad8c6bc77169f3ecd816627da019b3969f10bdbbb491181c5675da2ac92348c02a7bf53e93e815ec02f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadcb53f083cb981ef63c1d67aa79a0edc29577f4828e1295b5362468d114f7d99d4cd58869d564a20b3d164ab6cd6e418b0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b1e7c40f74e82d0be61269ae0d6ff909c8a701ec1b609283a53a85f6dbee0ecfa951d4dc7b2c8dad82210dfdd12eccaf197;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6af7c0819739d8d90ff96995dcfdc4392465af6982b09e4905cbf87ee529f27c2a5a11016d3cca563c707083db311301c0c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd985a8bb247b2a7eedf57a827c0198aa844d8a638d43e7e65d8ef549e64a517d49ce2a1dd7a308d3f9d441ebadb88a3ff32c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee983baaca4bbb84c9b8a5d3d63ea6319dc90894e3209640baa0881893b871632d8b65c9a22851c8ce4cd9f250831cb76ea1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72ca8af62c947e6cf38530026aa1fe7d044efc9a810666f770ce56344e941a2ad576a89a3686e474ae364f8cecc02f05d814;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdacf1b1e8222e3b0ecc715c1f79a527c73ed7a73c106dc310bce9924c15e44df43616b402fe7602244a373b4cf228b4f1577;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ac734f22c59cf920a9b7b6ad75f19a7154bf9e6fbf94d3ec4af20403282b1937fc4ff79131b79ea968bfe8281aa5a53beb2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h366423758e3c78fa2efefb98051fad5597bfb7338fbe8c59d77181df003e352019277de91605ac8f4ba83e95134d1b110ab2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde1c3033cf9eedd46f5528ee3d9668130fe204fb0f978585961164eace2125c03ec994588c291c62291fbb5ee38a5d5cd35b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1a41144eaeb7949b7c4c2fb07ffb92df0bf9fdb3257fd3b26c195aa136b340012f17317c44ac618163a4f07535cbd951a7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79a67c0dfd8d06f0868f164c6964adfa9f41d0c11d91e270995a491b032ef9c871af2874919b3d00a53f92a50991be80e286;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc17c39e9996933d2a526c9d83664f146de8d1ea5aba8bb100e84d858343ab18beddb2b1cfce17b487ccf3038e1fb7ec36af5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33fca28e3abd648d3292b46eecadb2ada64f1fd1f809d7f7bafd033d1ca29cf8be19de30a52f279cccbca30926c1b6084c40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2bee15f038ea74325dc137e813b9baf14834673ddffcdf2e6d86f27cc25bb07251743878a233231c2c3651226aaeaace77e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99a27bfa714e7a58cdba38109fb879036dff3d03473390da22b95c6947df1e457aafde25a8e78aa96e62d73b008828a9c4eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff2c7d7a58f6591366edf6b27bc9c0f314befd34909631ca8c191fabdde894f8a0323ed81b806dc54edd1baa0fe1409457ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11b28afcb623af369604052a1a07e6cdbabc0285d8ddcdfbadc80c3203915b31c997a4dbb33c8079aeea9a6b6517cf7634b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a38e5ef98b06bb250a96f5da5f18af9c2b136f63959b19f940f0d5bd68e45402c6ac4f57d12e2e1b106f99dfc0416a9780d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha21c6966908d7ec71ad613ec7da2ceb801786e530ac40580834fe24d2ae726f0c6c7b3bb630f297c00531d2a8280ebcae2b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0a6c5acf49c6df183a9546d3bfb7ccb1589503945059953f6b16008a828d57c842dd68eb5daeee5d47809772cac5d9163c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5081a7b659fb6236105dc74c7a9f8b720d15b0b2de11386c0d07db50fe4bf9cd84a0f2de963bc94798ce6d36fa9280519f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27e2604b8c106c10d55e72f8dc812c8e7ee11f10b9709366b11597c3057467b36584dab4869e6dffdc278cb7296fc69d6998;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8176de86c3f62c1278bddbb6c17766966ae2838b1439b36c5bbd12d1dfc589710bdf816660325b974f88a6c698a920d1eacb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3d9b7699577213f3d583105951ccd9b2f4c2704e06744b1a97a8bc85445266fe9f379a710a2026824cc8713afdf817476d9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65f3e55fe1e8c8eab7217dbe86594c2537c3b124294455d4ca1672d17ef55b5edcddf4b48c59ada938380fe61efc559959a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3386bc967e5630bdc47a30d9261f208bf654d3774319569169da8df16237730f56c479ca0f8e8926fdde012315767f86e17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf3cdecacb380a8e37c501fa3c107bcd2fef803a6c6c20b2523f0c6c6447ac36f292b88100f1f8a25c9832a72d7f1587dd2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3091d859961074fc98e68df62995afed7388ae2cc12109698adac6c8277a00e61d5e9ea56ffdc19390444ccd03979d03703;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfacd61f34cb815629ded86b05a2be3b96f45d3207c4879a7d2773c1ecb7417db6065c0af4e402a590840e07482235241f3ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae19260aeef44699fadab17081287a9a297f424edb162ce8a4f2dbd3990b054f1ef4548e8fdfaf26f0e02e357749f658ef98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8694654b5378cce77c18bd07d4aa0c5ff481ed3df13ac214904199332b179d340e45974bfaf711418159123f6386021fcaaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe6cc111a1737a68923e9d1d820aedfc06d286a8f57d6746b6b0c2b57f897dec10a066a7dca4ce55eb591caed82531da4211;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h680470753f09ba1fbf862183196ae8b7afb3c98a0703138e4850c294544c693a66f6b2657e9243f59ad5dc7404153c01d75f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h361e8eb922b6305cc18d465cefd064ceb1beed6ad4172de8676cf74e95e1ee64643866ef7bed438d682b69b0603aaa3750e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb290a1df76a831af4a455a24632e305266832bcc0ddd2e991bcfe9979daf454b0930550a4911ec51540467936c3869f4c0fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c65a090a9436e0d3c2085464114e2cf8ad124a28ce823495d1b7dc86ab891d27acb48a6af4465869ac28019b3358f03310;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cde214d37313a56f5b58334a05531af78388f4b64b410894d8a55efc3cfb641f3faf21a9a7eb9bf54b809494cc862700a19;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd48cbc991e04463ee123b036e6fb2bbaa178d644816e727c381b461c89f8592a124a13dfae021a1dc16be96f06002decb62d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2931a6c446e6e52b76ca4aff1a5e3b983d49dd3115aa317b10f5a2a6724218a5c2a10a2deecfbadf640daf916a5f79453a36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed553ba43e33d438576f4b3d73a05e95215321e9814774ce3f773115b4f21942b34ade13f79a8576d9619214878e1a66c86e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20c2093d35c9b340d99faf79ed4c54e671b3dec7e15fcb94a611db466b8a556babb4a53f61ede32aa1b896902abc110b8fea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h114691b1d3848fac154b90bdaa256229e62d2adfac527b6b0a67f9fd80066d6d5f49488207114dd1557bf1902200b7aca8f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha75c719669e445f083eae5f682d5b904f0d908f203ebde4635dea7838ad1162c24fd46896c4f525ed1c925366830c612956d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ab1306eb81f05e20af988e4bed1d16f1d1394c8b63b3e42404d202dbf85a7f585372ff1ba2c5c29510a481024b1a19a6a8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fcfc1713de111c6566f6fe3a22fae27d9fe8dcf0dffd921064571fdaae9cc6fce167d4ac4dfb48e8f4d5d5cb69e42db0b65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb2903a6903a97db65b6eaf500ef22a97e0e8b8d876fb353eb449f94f44db7a40bcf89fa544da04ea4efdd6cb0f9aff743;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89e8ec7f45a596d799dd4cb521aec5f115980b3359de14b39f2a0d6c0d5d3fc18f901fea842be88f51458b66ebaaa242dc87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45c0a8258a9fdc94690fb398b53e8557a1ebd58ce9f2ab6c8011ebd56a25c062f1a35497fd81f456198e986f679239693b96;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h404193b4a63a0351a215d60d25a138e686b04d850f23e907f0660938fc71c1cabcf74c3361f195516f591476e4501846c73a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20d3dc7c8987e24343785ff3dbe4ab1c09f326da40cb95248d7d4dfef015463e4c9b455e07fddebe011186f308acf4739cef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5ade92c1a3b87169e9437851835e1083d03ea8a1eb70b8be391eb65a336fc8dffeddcb74085c169bf454ff5209268b1d73f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95074f99cad04334f024d70aa3bb8656ae7d05c67c942c53a59948cedcffad9d57dc4b85c9a5d00dd37d8d28646bc6978c3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc07d693f2f1c4a0548098af062205b1253d5b0d3d8f338b0e56d8bfcd50d4bce1435fb7cb97ba8a28196703be3ee5c8bff5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd85b1b5bce56b43f1dc3033eacc4d8702d4bb27d4e55c3c7b442893c2b720d05474e06f7cb5be144e03a6c432da63aee987c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6e393bc5cb62053332b3616744fc345b51101079576e33e16bab1436e448a7dc59d5637be648d1b8d614033a7a9588f609b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heefd501b68d729ecf49825c2ec5ac842dd3d055cf0a18edf64c30367570c786419a7cdd3be070c34c70fefa38a7697d829ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a20b74923dac20db272c415fd2275b650d782f959a7722e7ae28e0a48e2dcc5ec0964eae7b6878282ce8ae5380aad060c3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85dd8e3f3753da0b27749d63ffeb291baeef23700ae87c6f9d7f90582763fe56cc2dfef586715a0b51944531719c1f559b6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9d46883e309c49634efb50613664b546af28e1475a0cc4911735ea833dd51755d7d29d871445d415c5126151a61c876aa4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e965ae4a6453a5c239107e6ad48089642349b2e584d397ad0065fa60ddfba6a9796d0c9c5de2b684c77fa58be3008bee523;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h632995721ca3f0b62d3a03aea6c5173d60d5d2e110129bffc35671b635ee1d3b2a23ad598fbeaee402ddb15e461a0d592727;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33994b5bbb5659d90cbb17f9bca512e03b9889b9fd8223449d38cf34f5b8b85ae9ed3846b18cd498960deecb2f7e97ee7fa7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd176a95b36e63562dc696bf9c2597c193fa53f28c1a25ddd54c752cbefac1fa92eeeb8c8f56fbe34d8fc67f8409eb80d796;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbf46c0b6632643d0a329e11ba0b68345bffa390ae476827c0ce8579a4437a6a13b443f1ec1faaa207b8d3d294669ca2a97a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bbb4d0b363ef37c65e2106b6d84c540c0809a9c1ea22538f076882c1d614f4f4f22f23a134f79bf089a2d116c64f6fd3a77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha545f01709bf1ec58e1abca54fe77dec6d1279439225923f7485b4f814d157febabf4c0a8ccedafc52785a0304630459915;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6344c8e00d5cb11ed03b77f547c9cd475aa281b2ec9cc03cb58164ef62014de5c8a39e2fca12fa8cdd452aae74c1ffb4ecd4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d88afc31fbf8306d61c59834e1cabc198896489c58dcf8c2923db9ecd42d586a0c13b3b99063ca5cb28edf207d21cdd282;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0dd7ad2d399387eb5b920b96afdc771b3c82b57f630ffdd28b01303d728601627dd2cad159395930504ee7abeff4cf7fb7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h392e172d2635df41c22a132cd482c43a25a34dbc91bca39f18a330276483af2d896bd6007c7e35d3458f66339fafcb668235;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34f76a2b502bbdfdd6ec894800a2fa62a1ac60aaf729471f0d398c58851a54791f6166823c6de3aaa90aa796b1fafb3f823d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64cc4af1d483444082ec8cbfb5da84aea537f57e88528f545c5e30edc109f3afbc2062a03487beb69226719cf64f68ab8604;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7255067acae2a861a3b71d655591d1554ae2e7b1e381cafca03b1d8eabbc4de9d6cb693465615b0d346bc50ffb69d79489;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b920fbe9fc9279b423d48806fd12a1ee2876e2f9a4a6dbce37ba3eacf11cf3fe5348769c835066f6f6103e92eef1bef539a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63d7353b2e3e397de1194bada1a11f8ebf6788093302de5457950854cb8979b6b5395dba55d2bcc11e886dde31968480117d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb97a58ffc4449e013de528f3e3c9048d8e5749d0de267c25248196df50987cf6648e1f62199c07f75c93963f5d0734524687;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27d160dd31b6f3d84f5c752606d37dc5aff15de0c4efb1860d981c331cc9a2156bf81a2cceaae1fa98b8484889822974b3cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79c7d5f825071ec26ad2f48eabb77ba2700baed48fd6a28210524c00dbf90501d932600175976bd946249ca28352c3b2f38c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63dfd10897f159888f5d3f0b3d8232ea34f674405241ac420dc8fa3cdec66fd74273cc5acd2bd414dc3c39b721d3305fbcae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a03ba0efabce8b7e09285fe6d5bf85f92e678b9431827524a991989fd77276a44884819da966e035ea70dd08efd9794a236;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbc6dff120200b9db14e62312d5dfbbe00d14dcb387304383007e6c200ac3044247fe62814d4280f41481818bc12095afd1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e207b23c3545e70260b7fffde55f7365067a2032da71ace4e92f9f0599f7866f5c0f909056b522a5fc0f4ce9add5242508;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4e7eb546d24bc8f23938cdbdfba1ad96a1044f03bab9d6a6dee49f05f2e4418d556589dc71f6dbd76899fe898b5d2b951c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d4c19afa5b6668be608e00c739d7d384d99058120d79b40bf85cc16c2a4e8b25b6ea5babea22cc046f02900f7f510318309;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he753c05a0d76b1e36db9756bc6dd113adeff74f842697c329c75afe0104bf5d2bb9ac09afa697acaecce19c585f0d3c5a3c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a3b321863cce4ce20a8ff23227a4e123f4af1b8ed48eb9e5290b28b269886e132c8ef0999add7a7fe9c2804fad4464143f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0847ec09f2d19aff85a1458c6f5b765daa000d1a3a348dbc9f2d496154151da58765c49dbf120a3d924683c492db2f5e7d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fc98e5bc762fff7f5a025a0cb668af61449db28cb9f25a6fa9031298b4e276e780ac5f96a9bbcf153d0a75b88fa1d2af94e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c1f2bcd4650ce0f975e450ce04d55b42568b3f099edd04ad2a8b92e6108aea12b8a4f907bce0c23c6a019b1327b3ea88ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a7de67d4795c2eacc13f7ae91b68444d0e8e1e894cb5b76b3e76d465c0a58be66fdc3d7f335ebb74b5a5eb6e1e9f4f960de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h921fd6ebb4456d5f821a8310f55166e71ffcef6069afa5ba50db1c18852a1e7baf575dd68b29a29ad94818b4fb1fbc5b2dae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bf106f653c7b3c87c6b1c15172e3141761cba18f5bd31740bdd8ae177036b80205f6dced22582801f5df8236f70c6866d59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h649f2c241d8d1d3715ab374813d04d4747e4ea8e3030925f5b1218b26c2b74dd90bea70b901506e96818d0cedfb445e99f35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc311d50112184ec68dc02e7b1c16b122cab6c62f69c2385615b8a3c5192ba2e718775d92dbd345a5bbc01fc40924265f6c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e35fe852d77c9193197c3efdd00c3af041ae55bdde48b91921f54fc70fada6b3cdee7f4ff1ceef219f72082f26541218402;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa60c40e95eaeacf33b2cb933f255c1b1397eea71f37c4c7351b31e08803aac61dbbd54b9d6aed1ea954c113de1666bdbbcb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40c00869351d3cb78d91a9abdc21d3233db9ba44dd2e1c4aadc11d2cd088fe7b1fb13ea3a733e929fc548512c0feb32372a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he837d8db9ecd7a8380aed7f93f039cd5834693b6904cda387e2f8ef128cc6a261e9a6f7dab6294ae88047978cb4866b44cd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aaa5d5eb1e244a91b982fee716f5d4e6645fe698481bba2bff8aa01710b2c8850cb2f6f9666d7ec43e54671c66a9709722c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52acad7ab4feba0eddf94cbb9017ae68cb91ea0e7a5865e4c67f8d1cb491a2422fb33e59b76da314f3555b264907e918dc47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9204794b3af80b9443f325d0c6a6f36d71ba036f5a23cf4b9c7667f1e5278224c6fb623d8af0dba02af8dcc4b7465d55246;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf63db8b2b86d46128cea62f4af27ca7053b7c89a4ee76405109174dfadbb9ecd4e3836ccadd0136f2f76c2f08d263483b5c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0eea243e6347a54776a2b15aa3ce607ca7ee1f88a8499914be2083f2be98fb6b22613c37ba071a841ceb89d9f2b78b27d70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h403cb302b5f45e3b865dbce42b0caf80ab7087062622846bfc8cdfea339c0b5a786654ae315207a63eab826e600737e8a63a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45717016b0581728908c141de1fb32fe1e659c39e90a6c28294392ae6c82ab22e12836b129169fa991c7775d2e5e1866fde7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b10e539aa3905d8b383bb0fa23cd0c845dd70385cfdffb4f1232f469122dabc6c3a058cffdff8749eeb725d46b28cd360a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7ce9b327b739637ec2655b003f21110204eea2c92df46b88c5038c5f4cd45dbf2f6dc54604a7e4430cde677c4300c09fd8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13de27c08695dd9cd479e37349dcefbef94f58ff3cb1221474fd3b38f71ef04cf6f6981bf6dc7090ffc1a5d0e12166e88ad9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d0bf3f68193b806fda2f8ddd7992c79b9c36ad4bd3bc92a2d09ed3228e8d6739ac2d73136c9b6da1b722b621a2d03c4476b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7fd12adf04332bc94339e2b3282a70c0639cba8198ff6a55b682fe929c279fb2cab196fd0d1e9539f2f3e75a036e1b3360a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4032734d10781dfcba3e2801c60c14b72102a7773b3c3fe7c99950b900c8c7ad8da0bd86b501b99907d84fb388dd982668c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e5e2d98cbac3bbf3dd55f3ac2c651d943dd960dde1595ad56bcdc9b77493314e8adb822c54e7a8e0da59ccd896bcd8ab48d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8a0783e13c5c32f3d6ee71aac147b735acd74a738fd808d39fe82b03ceff73a43c8d5b4809ab7b2af736592bee0229bb531;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99f90457b8727b87f50aee7707d20f28fb6d8f63f760c5b158cb94964526b2f87833f940d1fbe6c6d19e32f08130a962e31d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42b0d53d12d7a1ec2de4d6d8e04bf739beace31ed6e8b853b69d74abe40550d5bdca6221ab954c60350012916234a0a9606a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4f7047cbc5a6d4e31ba72ecff03cd702300b5f26c17b9c4c4a22e170a31d01b31507abe3079c0ea23b23a8c0fe74e3515aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1afaad93ce1af7ad133e78e6d22e06fbf7cbaf73397a5c2940641679f8dfa866e62ef10ae8131198f5c0ac792ff268e7e56d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha97773b8dd83a81f3adc68de6f26c8ba6784e5c3d870bc3e328d961093c2107bbfb679774fecf3478aea3873efc21e864200;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c904fe4ff8143dc6a54ecec851e4cc699c0549708ecd8462c8cff707db978dbeb4eb1b93be90f91b16460627efb26674947;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a615693d018210646c28ded426b5b915e599938e20743a82d60c274e91dda36f131a78474abc03b142daef493b00c25dcd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf0477b3d46b81bebc75ebea3eb36a1b1c20509581938b382151941a5bb825fd2c1fae1f282ef37fb459d414275e789af436;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9da07ec1aecc544aea1441c2d233e7d95e6ebf75017850b23121f21643ac0ae6924c4c32e9c513b8bb0a8f52a495c8f224a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd80dd4619b2b98cfeb8db5dd39e292d1e3da4a3cfc82a8afb84c20464810ebf4838e1d447c6fba23b395c2131d82913d6a0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5cf082a882d44193be380548db9d587206f3e26410c91abbe3c7767ca06578894457861959a410a0919bbb17842c71451ac6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84e560910851b5101a4a8c226ac56460a3b7dda559b9189b39c0c46b958a5ed97cd95bbcbba03af8c27438ac2ac3d70277;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a221f3020065863d4359595f31e73c745cfe73985f967d8968d9c024e57c2a40df33f50024a0c05b07a75635d02d2d1b2c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ea77b1a21c62862fc002a1fca9abdf5d1a7a48e257ae57c14db45083a533e356aad06ff79f1c538f6adb7667d8bd7e0374f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb97574cf6bb1b1a6745cb0aad101ce794d814a3fc427e83b9a69e2d7f15bbefb2a05bbcf9055779299c59882a637a481ea81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8079acbf53d0800e1a2a556374fcfcce858d764b0aa2c56b4dc7b289035a42e33d4fb54bda465414d80b160c36cb75556f7b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h201a1383f813cbe8645ae9ae5af5dc72718351411a01f3a2be438a54325338fdc6d2533df99bf97b75e85f2466e067658895;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha587c0bdf472f2d3b75a406f83ed963656551a8c25ddf95a4d334e29d12247573521b8adaa140395ef0431e44d0de4f2350c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2dc1ec5182cab454771489df530b1449e16b950b2532d5e1e2641b5016ff76a425cf2de07a0d39e0d91f857c3e52aef2150;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93a1e0b2a2bbea20a051e12d23d518e5d80315b20036f5bf3354dce971f4dbcdc534d06d67040e898b33a51d545323de71bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41be4077b16c68799485904c6852608ef2097baed2a04ef370857ffb037749cf6fbb60f6f80fdc57d128eb66fa28e3c1082b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66c890bb03fbef0ebb98d2255b41a19e81aaa83fcd2ce11dccdf26f4c9f3054567320d58c34859e73ba6d19732b185d3a735;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e848931b8b7c0be6eb6304c9d43e1f5c44c33c8a35e7b43436519f99a001cb630da5b14ac6d13908979827ca23b9edc1a35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79ec19ceeec95a444d662efd538e6fca284d7c6c3a440d1958b9b9c0800ac89700cc83963d229969b9d6b90af669443a1c67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h145ce82d54e5a0448949c9be634dd9b0f30914e77211c1b3a417295f814df3b6c81ac231d1f18c1f13ba76dfe27fc524b86b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd06bfec75c3a1a227743fcaa033a7a635ccbd6847b96b5c33ec80c0c53131c8851f0b8cb8a56199f820657b89f1130c290;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a1c26e4423d9c20a2aa3bce473739476de01a20fdd454a75ec19406fd48dcf13e835fecc52a787b7a242e20c0839853569b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha84ed91161d021f25731aafa58cab4b929e4789247e48fa54de5017f4419480215e380e031f0806c5e73e40a1ba4ace3e92e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ba29960367489d7bebdfe55f2bf9e9d17a4d0bdfa9c70eac20e6e636ba158568ff7ecb9629efdec51d1a14babbc0de99e93;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb50c93d8eabd7c2358b5e6ba1cc2b9fd91861d17fa7b3f544045b9efddcf2009783b72ca2be4fee4aaef752866f58cd505b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f6e6724fa2ed93d9d00a57310f83618e147c82a4fe118f7f3d4cc018c3146dc31c7e0def3ca555194b01141edaf55d3e1c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h576fefbb3e09f02d7bfcaa1af042d973dfd755cedce0217038081cdf0aae248a38f919b3407c3d6739ba67daac1a63744621;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h725a1557e4587e0d4b8f92f11ed9df8e96c4cca928df7f3789b3ae8a8eb69a5e6701636b289b513e998ff839a1ae60900f13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf11d0ff424253fd10dd7e2ed6051db534e2bf6a7f1c114e98eceda54168cad2634e323f44ce40751503ab35f9704c8b1db6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d8c2e48f832ad0523cb4ad8392b5e832a9b34a3c569860c6f078ddbc64ab61ad656c94165a3b4d28bdd3b73cc917fbb98f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99b84c39ae4381de0bef6c2d9f9f618877336037763ff3b3dc37a46857e7e316764bc34a4be27a4fc123eeab720dd7861c17;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1ec513836efaa315fd7386332f8574675baa422841f2f4347a46de59a07706fe26a617cfc7c6f78c8728b8823dfa3cfa7ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31567095b049be61b3c5fcbdbd9df5134870fbd31b27e6b83ba483a1c9b25fc20e9c8d80839143f6ac3878ee670b6d1f8d0a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e2409fd40c1cf54fcdd99fa91aa27ba94a88a1260e2a7daf98544aa23218f5bf1805e3dff48020e1f7924b2cc2c56674054;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2c8068feca7ad6fe96bb407bcb0b9e323d440b90e90d79a56f516f481a55494ff71e1b579233209c9925c21e1c4807742;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5722ea6cbb61df265cb813028442a716fc7b5bf87b8a5c719e6d6a9b3cddc660eb013afc1c910bb3e7b3e3d56d47b9e0b12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he64bf6e32e41bcc5a63a79cd30e60506fc3e7579a8fd3e7224a83bd7117d084d9c6588f39196ce22729c3886fa4fb96a7237;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25c95b89fd726f0c8aa0687f0059f44c3b89c0c5317f21b94c598f8a6059698a296b67874f2133e0d05642eb309b0dd20d40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ee6fe1b89610885f60e8666a1d5659a56605f9f5dbfa80cec724f2f39e16de7f69a3d5b14193f951271099f13b5748cd0f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb70ff194ce44758e6e40dee828973d06e200dc06e8dfc69ff9e41b222d58b9722aad0e8533eb6f376bc0978d2f7ce45c2f75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1afa0119579327c9867dadde67d6a11f3505879ee78677ce8fd912139aa956e2b12ef272817bfa5d0c2954a875a44551cc6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h779486ae9231ba2e722ac2a4098bd1014bab88dc298cca1341948911447895dc0816c46fcafd5217ce80ebb9dac4cba94d94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h152a67e67957e0b8028a13ad0ef19797f31ce74c6f7edb5d22fa643f662a69416ec7cc7dbbfb27e5c571bbbdc94927a9081e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21b4e48253f5808f7f1ea8ce54819f537ddc9edffbd990d8f095d0088c8db676e7e888efc2c773ea61441182d00e80350715;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfeb9912303f245a8b94815783f644d60a9a621b579e7fc2ed7192953c78692846fe1b501e0b73bb2954db8b42dd0d7a523c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53cb892c930e6e496df2760a26cfc9145342ef2d6ef88971aa2636b2c2ee6e7096e631e5c62b4737736f73603d7654a6f9fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47250b9c96ffa2373cc371e323ebd307c9b2b046c71b1199111da57708ce2565fe64ad94c762844e245c5dd6d61d679cfda0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64872400d08ad77775c2140bafaaa716384b2e526682c0cf22f91f56f3be220026fbc4f0575bc5b00837556a1d4bbe4b12c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h718fdd815695fb6d50e38670afeaf79b64f501527c985fcf4efdc73b34358d2c21817b4cf24e9556112b2e781d854c234f9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3b8c8c2e8f9b9db2cb12f07ecdd1f14a9c8298e9a374ef446a5cd34daf176738e45406b1b08ba5e398a3c75a63577cc3724;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80165541423fe2bddae9070a4559f67760b8f7035ac77c4d8b77c8e97664aad0f9c2aa4dc946585d24b3132e6bc01fbbf87c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4e63a366a623b3d27dd7bc5fb9426a5492f502a754471f22194b998c28c4648a8c76217cdc3f997152e441b6fbab1bb5341;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd99b94967de4bb6516f1c2303dee2ebf42599115fb207738cf55e6c9c191f4a1a723aed1354048299b56728664ada02bed4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35f2d6082a007634d51f979780267c90373a3415e46bfbd039f5152b08862f868122b6c1c9dca22e29517a9ee69d60c312cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3338e15164e6342400bfa5276161dda303a9814a485f1c6b6e6f716f5287cfcb1c5b6e7a58040f31c0cfc57e0317d0cf01a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8f9d7256e0e50079573ba6a397686ae9514065f1bb07b8e32c23dac45587f9cc38960391a718c35464f93bad94b6808499f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c94e61f536f9f02d22c75707ff50b6eabf8b6d35d18ebe0e415fba0775e0a350559f40db6521cc597f4106d6219c4ca7bf2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26cfe5f8bb2f33897477f0bcf1ff1c812f73dfb0ff49f8cf58e67c34e64747ca281cf0c731a02788a3016018c291514001c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he332c774876c92c27c3988b137a3b7f96dd2a3dfe07757f5a4e9a5a30f60796f826db03d976e8ed18466bb2cf1d8183ee661;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44ab5582945a0d52000bacf8c9fe005bc6464e097cc787431ee5520f308cb9091d99161bf85419ba4ef4a556f1fe44c70bfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdca6e637dfdc2e1a4938c82434e434a1a32fed74739b790fe5bf6db87782417baee7f5da2f9ba75426a18cb0080174e21376;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68fbeafe71fcb4f323e68d594322c1d6823054b7ebf7a30f38509a670926dda3b04ce4d8342a873fe110be1ef700fb88d475;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a2ca04609acc0baffd6be921e201847e0921122e404438820299c227460875f4067f28041fd22e3d32a1d8e105915ecb1a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cafacd23fbdc8e6b703eeef426b2e5dd51e50bad45980510fbb94d96b21cfd5671320b9f5149e6401687066327a60c6e6ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cb4955aeee0370d7dfcf7199e903c14b72105f7798d4b2b3f244e561404a88883df16a9a83ce417ee03c0dafba49a12da95;
        #1
        $finish();
    end
endmodule
