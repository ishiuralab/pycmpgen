module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd6a5d84a12a62bdfdf4af7a9eb3b322b1437adf7f41e0ae2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a41e649e4291509d8d004eec4091a8e15bd2c0a7d70a76b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50c02d0bf750f48c2f8b16e479a07e00d2c5a9b3b2b9f3a2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0a81134318cc93f1cf7081244f84fd40f3c05423c63c17c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5dfe3964d55f67f7f6c53a2c063d990010ef2fbe5861c27e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf06f8f649dbdf387eaff13c5cc7f59560df31236c5c1a0712;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7636d87bfd9a02a517399f6068538155ee5ebcd59990bcf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cd8cab45c9310e00513d36b6847fd77cc919dc7211e515d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82ec0014fb2ba7e63d6898439a11b661a31bc3e1edbe0c5d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93c9d1ae39183774ddf801df3b9de4fecbc9151af06c49239;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21ff596485c73b9f02543624d6318af93dde6c2cb7dea4585;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5c9f3071f025663c9931161619caee2034ee7cfc50b76480;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c3609be0353763a8f966b0e5af273581930cd5f9da8babc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f8db5ffb61fd6da8c0456b8a900425c8ee4e0e0db5e81ae2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8aa14a0a2fff7959a77fef082cbdec6caadb6dc269b370fbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a1d4b2c8ecd9130778d3c3ffd086cc6ba570f6ac997fb3a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe1df47ccc993223849e4ba7b1c9a521dc0e6e9713aa8c528;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99b50b223d0e1ce2e82533a1ce3e4dd2a718b433eefb2af5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6886731d61f89f90bbafd12385de0b1819fed4d0d956973fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d665faa1058127e39e4238aabe535e0ea4bb9ad6f34ca74e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h510b8d7e1d4341ace3cedb74a8c77981598b5b080689a3fcf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc69991a9227c00bc438b2e8a52673b61c52f9d35ef56273b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7ef07201c078f448bb3a96d9025900d263ae5f8923b7f921;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb1571d02e83b2b58005a7a2d0d1c1c3feebc7a1f348ea521;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he483458a6747cfef84fd49cb11d1ac91cb39686e78a0e88ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d1c07c8b63a633ca470a1cd859615f8ab11b54f289b19729;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd961aa62fbff7ccb293761fca709596f4df8bc456bfa0a62d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he118dacc6e46524f9191489b46a405019b243243a8e1d426f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bb89358b248c9fc001bbcab44b380ffed66de385014495b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6125e384b97602c6b0de4ed3131b64f95a59a840622597e56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1b756c4fbdb7357adea40bb3951cf62d7e066b4e86b35efb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h372273bdce7df4b0b41a01a260e7990baa81d285273f74d7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc76d1c6e9f5e0125aa84812b81e922e02b7f0094e01e8991;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e0fac0877cb07d4b1c0e35261a4c60b8d0c77a7fc7ec939b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcca1aa522a28560c523c235d0e7c1f79539d513b04056d0d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5c50964222aac3a5b19585d7ec9ad8563c049e3fc125ea93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h332a4a286934fc290b9366edebe08a2e07cfe0d99a80dad62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71cd6b96f58b7d5f70bf0b281846d11ef74bfe53c81712a56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcde570014b666a16d3ef3eb41dfa84da945cbd939963a18b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6fd81ebb25a0d1fb9262e240454710c394537992fc64f4e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdf88cb28a810b31d1227382805eae6cf8b17c44e51397405;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96eb7cb9b325b1029c4543cb4cf7c9039dcaa5fabf9aa94e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf834d650f35cd14b96a5c4a252c8cff381097a4b3c0330c8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2c47be586641a11bb31ac2d3c8c06d52e81b710b2b634ed8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45c03ffcf0ba71f85718f03b906094741b957f5c1a7538bad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbbe19a325a66c4df26881643a17a9832aa9aad3cdcbcde37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62fde3b00a9a64c812e89a75f1514a7bcb95062b5b8c98ca0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b11cf52e8cba004091d451fac5c22ee847aab92723e42d45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd64be038a3338407d5a7f964523921361cde5aa5465ef8b07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93a298912bb4358cc69f5e94defc46631e98fb7de0bd6809f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2174c81265d0f647f29a5df059e90e48dea04ed9c4648cfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c473dc80d1ca99354258acf123bdce386d43500ead4442fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd8244021e4d26bcf0ece1722143b9f55f7dc704215c08c4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31b0d9ecbaf0f258fa164ae7e77d27e9715df7a2e2f23011e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd372e376c3625463a84aef99c3c2981d5b95df0e8b3f29bc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdf260d7bb7b2c18a23c83371e3eebdaec48ecd86cf34d572;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h846ca54d025ade0bade7a8edbc8ade7ddbd54071d72cea350;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he77afef12c6fa7ed82447c8e01929a7a8ef809ccf5adb0703;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4e889c2e9eeb64b1d59dd07ad4ab048c224d2a716a10f2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9469330aeb6ada7161eabf84afadc5517c00a31e8535a7f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0352dd79e93fa8e2604919c1ab880e6ecd1267e12f45a7ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2815f27c7e9965c5982ffdbb48c5f40323e1056713117aa76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5431918f578ea81bcde8336ff4c47d693faeb6a5eb0055a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90ba6a5924b9662e3c1aa328fcde88cf774b531a8c188a341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bca8fb412e18c9876619ffe5f720978c43d176a6113e999a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57f0290f2f88fc7198700dc171b91b2f6037c16e34af7ae0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h737dc79ca83d4c8a30d80c082a11a629a5872286c47162dd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd999202818d8b4557d6966feedacc12d3be6dcb92713fd95b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb47f76845a00e2bc2354248cc8b39fb176b2924623edead8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5405791479146adc333171ecab4fdf12a5a59c72d05ac5c8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f8fe11f3ecd8a4b8fcc75c8eba2b93f5e0864445556208;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he070347c5db299035b463861ee448f36419b9e9c6ba4b7333;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41a3f37486d74c569ec27f12b6d2158c9dd25aa608f638611;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfae8381f1c2a6178eee22dec16ee690ba04ea87c46bc0f602;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h664a1e7e312505ad359568921891ad3babf216e5e7fe808e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32aa04abae7f28d555b1b6d0e5302b92d1cd84d8ae21e0eb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7fa9087661a80cf99c5b4e3dc39158ad9a208639fe4aae8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87457519cb158565228afdf0a51da2e496827c6fa4f9f7bfe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c9511de25de34f97f4799374188894ff86ec81b8eef6810e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a924e00c32ad00df2c411743c53646666fbb103d1bedfd64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h697cfb77d793e7c065d5ab0d62784f6d44e5cbea05c374f56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7858831490c635ddf2d7fda2561cbd83ceaa35feec3322c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha22c14e44cd362da9050a82e5c9f159da90009b7b6cd398ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e0a3c3256eb19fe259034aa7517192532dc3a45421107fd7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habc20f3d3e864cc8398b764a307999f29485aa6d1df551dd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40df939be4afcf175f81fe7081daeb531f640b7c463c97318;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7fc643a07a544bc2810ac0ed7e516baa451dbad845f95d47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ef70ac646659880953612c43af0f404c54ce96614ef26205;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f0a63add5cd3023bb1266563d7519efe16c7854fb28cd66e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92cbdb2bfb4a87f4268fe10f2c5cd848937adbc4e3089d042;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e36f176bb22dd237101f78be76d87d34ce5886165e6ae4c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cd8f9579c0ef2e8d0f63e881c3c23849a88000d03d0503a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45e5344947526e12adca24e9d2176946020c489d03fe6a3c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8099e5afeccfd0da78e9b776cbba6b5a991e80c050b8beb24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93a12b12317238c555e008246ed6f3fa6102aa6ca5cefcfde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42afd15c845ab83d4241f11de9b66f0856a0090c59d8aecb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h571498c89d14d34254bb528be44780e71d90e7c6fe0eb17b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a8b377ee216ea1ef834bb07b24d40889aac4640d0f33c9a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18ccd8100102ba6f6adc76aafb2e824c7899e3d1d30d5f547;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1b7b096c5321a26d0240286d4e5faf31322d37869ad9302f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb52c192004ea2bbba1d6034dcb17258dd5c9a172599eea64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9094222ad7843c09e307952c5234937599e43359e0f2e5e90;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f94c948ea0e5dc9ec9e3334e01f530d3c8dc056513ec9980;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48a5365be56175eee7fad8893a06f3d79842870504ef40c61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he118c49bfe12885a3fdbd23064666a077ac3869fab23ac932;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6037891da614a4c4066b78aa832572194256ab064b4d6e4d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d4b5f58fe2fdf6e093afaf0a387ad358c35520fcb9969246;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab6e88a7b60d747241d14f30c98503895eccf10a72d80f2ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7be6171f2d1ecde47f73dbd5f1cb2f0a969d288e1a4b9625f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d57405120c475f0224efb4c068b3bcd1138abaf0f1068146;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ec0e89230851c249229fcf51ab25b54d0171c76ccd011f1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1862e8b48cfc2653f77b72f4d44c4c5b221abb633c3ba5cb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6d87b157697b00e36dbbd795ee66f3d1b587c164fdefaf07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac03a436e738cbfe6edc0444de88bd01507f46611d3efc887;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf0a214fd99de55d29d31b62f90e03fca3d216eb0090592e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc70138e2c4fa24071b913e9f7e13f065fe939d8655823d31;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58728baa64bf4ffde496ffdcd0da3eaf2717dd7f6a607cbd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4c68fd49c166cc4394c58b7f5c2547644739f5da01c708fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72ebf56f510fbb4152716f6af2f1af64dfef6bbdfa7a4c731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebe7ecb1d302db6b0813e006129040357597a8b3f97818641;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1ba615952fa0e8e2eea40e9891d097b805a99dd06a25f999;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbadca4a066fd1784b4a2d05afd234a6e52c2ae1b0a73e33b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f45b61d37e1e6a812ad053489a6d13f876b29d9d1a9ec9fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha73060ca6e808dd17ecada9c380deb15b7ca6d871bced847f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72ced9083008c805535022d7db352af67a1598ce66fc0bb73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31e227f328e65d88b641cb2f3a4cd31500d3f214e539520c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc63234efa0ba7d89e8fa3bb879964c607007ad3e3a86225ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddf95224657a70980855a482147d3ec6580c51495d18f51d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99d25ef361f225fff7b9278380b2456c7bddc3d2cbb6b3256;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9845264c7ef8203c165cab0809e42abcc4bf6429a2689519d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h769b179b7ae1f4b1a00e11ddb9f5302fea03d0b450895b91c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb166f19d3e3b1b1e4dd3f706c9bb72e9a19eb579b2cbb50e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h178b898f9b65d58458460a792f495b144406790acf715cb7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc14e2f16b0aadf1cfa3b3c4e10925070b277eaff6abf40619;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6950290f00d61c5f3c12f540799669ce5f3c904c1d78ffa6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5858a9438a1b5f341d408621f9c96fb58639d7ff9b6252be1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3776a610339b507d8fce25a4a893699ee090ae37d61c72ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8de54f0d7a750dcc20a69d5d1bfc901a2195b2950c7e0fba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haae9ae8b80936b5756a841cc49488d1fbc0df1fc0c77cbe4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93a8c0d7cd081b9252411bbe9abbc7bb8d1160104938f1fbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57cdec841e7af9af35638d0af22d86414385d2b633234adf2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21a6963f6a27e565eb5cb9e2c3976dc5e2c828795c79fee89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79eb95287d2a79a88266495f88ca80b00c5c33cab44ec4701;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7880e8741fbcc085bb8c1812be3654d51c593e351c2d1f03e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc009fa06cd82b1955cbcc1f7ae59a73eae519074032ff3e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdad34bf9d31630d9b4e199a82c0beb815547fca2a2fb1f60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30fbbc20d4812a764cffee7bcfdfdbbb4fb0a3fce1580f8f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14511e7df2a3172eb73458b4b529fb6abf6e626b3ceb84a2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h343d062fdab7a2e903454546c00ad8160f0f7509202a5e6ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0503b1d7c308ff5a23948654bb39fb562ebe3fc93afb1557;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h464da33e816ce995fe9ad22e993f7333f940add9f5de0dc86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6593f6b35544b517ee7a3f29874215f7c779bca135a4e95c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heed0463b73de25bfdda505532c10e8a4c9a114b9463ff3263;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7ebc366e480e7e3fbf91e30edbeacc3c0179d7b5701223a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h378b62cc0827fc65f65c3d49af06d4314756e2f9d780cef9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd0c7aa1dd699275608f482d2c81169b355e5872fc0f86a82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b7b1952db59cadc8aa43eed767cca3b0b99efb985a1ce367;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf072bca913b6be4b348016d930a34ab990d7f0db84ef090cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5df1230e01b0b13d18d2abe66d4894bb6876da2c60af36247;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc4beb1bffd7d86a4febdefd692814647d71ded7a92186f8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93c26fa514aa1fd3cd8cf5f8fb57405050749518caa5dc1c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90eca41de798007ccd1ef93a24e55e45031c35a54ef195166;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc790ac84840c515e919d6e271e5cd389a44598c59526e95a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ce420a2800fd45c6c4ba15bb633fa021933d8d524d5f0172;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9932d53426b432b38b31cd0fb260169701e487426b5d51ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h690faab02ab6447ff6454cfefe5db6bbcd5ad5870506a5b9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81c2a2d06665fa37c7a352c7266dc59e42b30ffbf8d08f21e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99a15cc9eea3d546df4032a5c1734ed23aca5e9faf0ee91e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37d9b1df2ec4f1aa4e9c9b200e78d580c6a0ef5ead5e0c73e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ae23d9a2a96503566759edabfc140fdda3cb68cb9f7fd5d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb46fbed72a5c5189294fd9fb5c17faeb4994d0cbe58491049;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd2bbad08b7ac09c95f05d14f6686782d80a801e7f5ea6908;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38c3c0050840d5b57a816e667af2f9376947d86de710074bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc54f744cf1e088ef1262c32b29f887c7ab9a075f565eed0ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13460527622246878b3060f10a4382c7b6dfde048696f93d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1f8350ae7b8eca41f76ddce83a4e1232735c30549ff2888;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h882e9634f05bc40ad6716e97c89354ca274f1863b8c4774b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bc6e6e16051d49cda7c3cad76a4f929cc516615f8ef8fe86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcc66b8413d7f56b22f4daed8936793e276c14558e1fec1f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h715b7b7090940156c32711b60fc42a00291e37e47b6d9368e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f7ebec3c813202b5c18c081562d017dd766a8c54aa0d5a81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70932023eca47611f0283bf86c441470b5b1287dfb77c687;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f2461511d311a393ac5f4e28d3cbac655f2c1d51bb9ca93b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h295af00d03c86d4a426b7537f67af8ffb93916d1cf9ab6fe2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42b61ddf8e24a41ff13746aa5a7929e65b1ec2181f9fa7ca9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31842e2e80c84f8493bfda3316564a7755cd955032606dcfa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14e8fd8a1f979c0b0049c5ba059ffe921632c04e768073cee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb53f725fef83fba90677aabd77435d1116067af76ddc972b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79216225421e2a1a366fcdd88e24a5d2225f8e7cf907f1e0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4fbc8a997ea4ca14edd69e17de5fe1a6a22c088cb1d0f7af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd61722528e1b31154c3e0b86f82d3617d5758237b72eefed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fc6f66a2ca7e5a563d67a0cc54e4308506c733fd302db69a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haed900f5a17b9a2e337aa0e408804fbde5c5a365d6167203f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5928c8fe02e65f5ebdff8918fc5687fe8cdfc4b230834c9e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h575b5340aeed0638dd3397330ed8aba9f72751335adb0db4d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b77c634de983389aa69054c9ee7eb8956fee2f341fdb5991;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a0c081439ead40d440e1a6d05dae744339f10bfaa9a23fd8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haaa9ae6bc0af38a181c005d4e991b47a702ef0465dd921433;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9a35381f44bd7eaaf94c1602ba57221963d9703730e154c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda02821745e2bf347aa1673acbbeb1e408dedb6f94465d8f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4b5584f3052e8bd34f1709718318655d8d002223bf857031;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf7c535b296e121f8a31faa9c031043f760b78c116117fcd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he065d355f74334a971051569a33db15ae2a981259fc72efdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcf0f3dcbc12e8934340d483454e7dc7dfe95c39849e03b2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40c30d2a0b18e4b281a3da493051e082f747652e70ea9db94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he968203101f2222681a71c82d979939fe202ad2836efeec38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e94ec5c4a37eec4467dc7037436b82d6b463f10090cb4710;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e4c56e27fb5f0a60271f436f60e4ebc35e23fea851e9aa7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa0b76a2bb57a05f5158cf1247374e18b37522332b5480d6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d15e4b0d18f6be45b2ad9aecb002047a504e923d485d9c75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1980781cc9076c9e30f4d1a0ea64ae19d0756cc77b90c7c68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbdd4b08b058012a0c0cfd7d062de4e9f270de982440e7219;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22d8fea14bc99355593e933bede43e3b61a8151822e32012d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb86ed71693ad27b6bfb6b7a647e935e9d5597ce09a5361089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6dd9fb28d3076fd0bc15e726aaaefe9da2f166e627ac8d98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c6ad4799e5e0e7338a20602d001ee306508a96cd4a80cb1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ffe9c914e8ad0453b51803cf7c3f6f790aea135baed6b6c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha74feea863c8666bc4b0a51a61f9ad7190cdfde4fbb32656e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he649daa442768c45f4b7f3c5a4cf19c3bfbf698096cbea97f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d3edf04b4b4cbdae1630f9c05d3e59323479ed23b9c5534a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadf8ebcd34a6ea0af4915b986abc7b01e09f1e353ca7d45e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61b048f326b2cf7c7f4b76c105100426f06fbda86c1115dde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8e2fa191af07e12fd7f0da05b9484b61e0dea023fd74adc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fa7039a5926da766ff2449632610b271cc5d809d656ea43c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3561a9368ae966261690f6cf3c0795656603d4b19ba9eb04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0c4c3285a80888bab2ffb6b73158d4b331c4f83bc36ad4c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha51cdee01f069b3e2aa9a0487f04f1d5da515daf6f80f6bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h829b2886e579391d61f23619d01c235a45e1d5eaf6fd5ea98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7af158c235aecb7e11a7c0120c49a2614a747230cba918264;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2163f978a36a0a0830666e400f81330e8407ae50fb89947fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d5af513340d328e1dcf66181e2b23d23c36da686c1a2fc9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ffa8679c3b769d7699822e0fb3d8a3a32b892e9f9f5126d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f3e22560d57a4233949df3bf3471655e51469bff10e5fdce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d3e450343a49bbf049a837e5a425f95acf5c6c36a39b673;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ffb7a32f04fc6cff7cf1c93376e06fc3c2c2eb6af9bffa86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c01b1dc90b53c49a1a52ae42dd0567bac3602575745f90fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcd2a647b2d8e082bdfb1601e457bfd6ede16426a4d9f312d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73d52436c383ae0f067a5a202276a3977a7d6bdae5be7c85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf97555e8db3f20e4dec9e7968bac3ee05b154a7b5a23fe9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd468b290084708a9a4ff005beeed1d27e8a2f615127c7bdfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a35e15240f2096c5cabdf5ac6955ca2a476c7aa07821f0a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe2a444c9e3b9fe048a2827251393f6a4cd43179b58c020d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a0672c820931dd315e90a59e97053c8826860a3f9da4f435;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ce4ee0bd16af060d6085701ed2e0483b3b282493a502c64a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e5611f730dead020cc4f5e5a078ac9173aa5b638b0aa2aab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42682332b4ac1efa72ebb32fc347fbba0f50682e341b48603;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb783617ec9dda81b41ef7b4d79c756786d96b8e17106d9a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h186de4d88065a1c39673678ef81af616a69adac04185de7e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7da0aa36147592a4a002b8a455d4e3b78b20ac9c5af90233;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce0040b02d322376c45f40b65ccc4779d34f1564c28da3be5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b1d5131e3873ac34de9d8f53801e339a3099e487bfcb02c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29f486eeb481f8b0feb9a735b1c854168f3020755ccfc9362;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7e087a0ac7ea1b40b200eccbbb9fd96a660fd79e62b15601;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0a02859d41cb25a16b27072934248e6386429381b717343a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bbd02db186d0066dac511c475b369809ee43c72fc36cc2f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h631501569ccb08e4f537d7aadde6d59e5c6873389de7ed86f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc73d61eade6738c2640e0719399e54dcd8221eae2ebf6dcf0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16889c9237445a1866e68ce2ea11933bed97294ca6a40f56e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd20fcae8e32492a833157b600a6a35120da4ee871f10c7117;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h607b8adca180de1713c998b040076446aa47a51eca3dbc2c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbdf7c588c7c277240d3a779f06877b8a0c57b50866d2b38e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h667cfb240ce7b0c06be2f7ae61ff9ff045ee9e2020ea4e1c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcec6d114d630d1d072fec124a4b40234e8225cbde148cbdf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9060fe5c0cb5b03856ddde9d639502444c2355b67a0f4af7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2f28756fbed7445d50a50111db714e984e660e9023781ff6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59a18592e143e8fc8adc76a509bd827b287b5471356e38ed1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd291289b22662e982266c2a25d15661d3543f50b53095a321;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a1fba507c5fc75221aaa86b755682db81176910ae9b51bde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72bbf6d4ad436fa2e90df9f008f224a8bdc6a6a6366d15738;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h947985d2fa4fc2d0e23f86ffc873582ad2e719d1d41f99abc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2277808cdf0cf3e1af4031e200f5c0a58ee2fcf9a5f51cc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3370d55660d50e5d842d95d384bbfb74e7fe474d03ff2633;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7f7f51c5f6786d404156193df10265da59c3d2640904fab6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe506f5c5bbdbd5e201c142c5a73ed9b9d0905c23c948083b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f20e4e041ca0a9028ef5b84113c4ec5cdd1b649ec90d33c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a26fd548aa762248bdb8b47faa699253668b22c53931b445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85d9a479b784209a6486f7e392cf4912f3c41af20276d184e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6808e4612cf3974413577c92998742c2f3c9178abb2e8c57d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2c2f336b6699ea249d78e55eaff85fb2162b124bc33dd468;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc63ede7da62b44d076a9904e6c4149790564c0a6742ed0a6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11e964f0c4d329229138f59fec659336cce7d7218704e7fd2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7758704eeeae45ebed1c4a74b1394862577e802a7717e8c37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h246e0884637679b40fb4f49c443c30ca63a232d86e315d23b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he781da36b268c634d0634bf0a59b9f6e1b6820d33e75b4c49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27ed1e0118d7ed6086bfa4b503500f7dc240a3858d79256f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h371f96099e7b18d4a940787ac4d9c8c631962e178a010d093;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f1b307110707d8d86cd78d7a4cae92394ea8e5d6d2984592;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fde6950aa939eebd129627269d427ba9a25a5fb6a44c8225;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h474a2f8ca1bf7587a2b94d17f1de4c53939c448ea215cc336;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bc0c4188b602b238c0d0d8105d4ce990b113a47168d1d059;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3b6cf34c84afdc98da79dc5d02f1d9418c5033e4744acaf5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6a5dcf28f53360d7611c70dee90d3526ecfea9d2d26f1318;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78e91d35529b721d793d6f31345a02b0e6a1205e9a295426;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha65ced8cfa3a7f058d81b288dfe56c0cebe2f52090d3cc4f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48152a9a9875c826ebcc03eec97af9a6c6773c7fd74685e2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bffc356819424fdf886ebcf95e811e763808755afe62a765;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c51d54caea8673be018d18166dd90a6497fd1671fa5dad49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf14ec2b5147253e9a9c4c2c974e0a3ae79e46174770015694;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf839964a672dbf97aacd9006cae7170a33bc027c40304c82b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h362357f841f306f5bba7ff15a1f6b5aa502ac3004d4c73ab1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b78909459598d1c4b4f8c02c64e07005cb67778906c536a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6ab5089051aea667a9a16904d9e9ce9a198d0675ad154aa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9381dbca5a31ffcb9c32014c07c9d0ff494187ceac2eea49f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf9ec7f967764a76cd98f6fe8cb3326ee556979ac78d99e00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fe37131c05d6af2712f785db17058b04e178b2b26154419a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83d919e908ece75b660112a53c8d9666a8266d79c8e0a2705;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc366c99edeed4a718643ef19d5579990eddf971098f58ee28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5443a94f359d3a0bb440da93ef16a13f8571115cbaf688f59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c5be26b80972a8c34b73fd27c77c4e9e9985bdcee27c1f44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fdc3fa15e05db9a41b91cb9ed3b669e5e9a8a91f2f3d3686;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8fa6f3997211017ef9c3aa8adbc93654fafaac8071acc66f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3635c5f39f540f138a96e06db288421c35a00ce1f7836acc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce3cc0d3952812f45c0fb264ba90b4c83bc3d113403d22956;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b516226b7aa47f4a90ea056e42bc651f0d5d3a117ffb3d00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1766cce6cc2bf0f28ba060107d95adc690a7dabe20b83f329;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddc693898251c14804491c0ff9e46e2a711272226b03615d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfaf211c951730ae5835d9b0294a00a7a02f8de1d4a8cee0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8fa5ebbb67d18fad4728e2dae6752c22aed68df07548fc6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2da2a354c173cf7bb03606d91774bce5ae2d335651e48bb82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3c2f63d4f8c343e918f0670c63c90641c18114542cb69175;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c6065c78967f30d399ff7c610bf90a5c03995ab8bfa55aa9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b068076f1c2d23feb36ed6c2fb13a04488188b95c5eb19b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha404637e0759fc22ce99aaec68c79d67b8a1a28497d78bf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1e75d2ce89d1d58d1e3dcb26e7c0bd474423f2b45b1bd63f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0e7a00e237796a5282d1e7abdbab7763fd97d072b5bf824;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfdbc331e8833fd719d26ae49c02db736022de3ac6ff04251;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haba8a3d30dbdfcad2d2372adb1ce7366a844543c7b182c1f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc400cc2e0e15970d74e1172f14ab1e547063bcf5eed6d0ca7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h425b82037bf910f4241386f1e033056ab7914e04158995f85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12933d84f584309cc6b71e034df23be233b5ad5c535419a77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98ead5f707028d8e17eeb947b75d523f8276982bd29679714;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he73127b34f2586698eceaf01b6023e03969dd002ef988b5b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb13296ddede24b5ccb3259b2a12b43afebf4faef77c864c20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47995bfa8369c0fb0d4fa9e484083a997f9a7272028b00f2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb46ca89f750a1f3037fedb7f101d5c4f73c9ba52c293312bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cb43e75756db10965a2e6fc9abe7cbaf231bf0bc2034edbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93b002d3a443818630e9715770df7c7edd2e1d0f729d6ddf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62bb17eb25b2a39bf0b74b698649d675c6a8858912c899154;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6617b2ea099e51b76700997ef00f8efb3b9ee371509d1d001;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h448cf2b1c23b943f319521c76a65c4d418a83496e5bdd0dc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1058c6c342c13329795b42be948d5e059a33d2badf4854c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1443b16a7cfa9a7c09d6fb9f7a29def1e068fbbbf1e9b48d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h722221b4a4e2a5858c32aeb4766db08c03253ff8b2f8a55b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h218ece27c73f0611e3ab386221ffdd8979c7f25e6400464c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f23b7dc88d916cef82c15d86f98f2c0f3e8f376d4fdf01d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9188e145b05415ddbc64394beb9bd3ca51bc8f540e718f65c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc85b0b6be55a57ad969126f413f73221c5d10f1aa22c55c98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33b01b1b039d85786f58dfacc833ca592e4b1d02fe81d1609;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h908f65cddfda1b40e32442632e18b64621d807a52a7bc7062;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha22c162b3409af85a16317bb89d22318259733bfcbac369f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27277e27536a4ea3dcf0d272df103ced2d68cd968b3ca4c11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dd4f5f71f1d432db7558c152926d48212452a745c239aa0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdca6551750e6047223b9323fadd7d1a31aeaf40d9dc7bbcdc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8566faa8f8faaa9fef220d355fbd4b68737cbbf7cb9fb6a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he356c9b0f530d45815bf94d66cfcee23d5c435ef5cb5f454f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc116d8cbc51025604ba5a55df1a28227e650b912f0b6abb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h763a0497cf09d43566cde38b8dd655e0b4974bf8397c8fd1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd04dc890f81fe61e2ab02a8fd31ca525391e5f8de402bc3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha78576f0e6fb45a8e182a8936a253816c5b29547559d0a055;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccabae13a763c778a0a5603ef7208f01ed06e648a2542ce5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfa807c28aeaf73e4adf5c06c8ed2e0432fe0b52a665fbebd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac902a03377077833456ccdd8dd8f5d7009644d46b7c2bfbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b71e772fb21d1f62857c01c7afcd0f0b91768220aae89020;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc234eda2a92c4b068dc4b15b6b33ee69cdbe002a40c03eafa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ae470be6ba12a3bd3338b36da55b43fdc42d2ed839fc7db1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc80f40adb555782cb3d47ff0d68c52a1b57cc359958b2c3b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf1f882e7a8be1e1a84848dda878f87a4dd4b61f16704ad3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h716f1b717c4c9e749f6362c89477d6b8fbf87d4007cea3971;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24a0f3eb0c461e37288a7fc01608dd0ac3c3c1eb164e428ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf03bcedd6d39c7ea36a2ac77eccbc897fa5a4a5011072122;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a4fdec7e9613d6bd13a2a47c038b56bcec002353b0b5e77a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c32f4076b01ff25138add8a697c394165f22f0cf7d6f49a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h449950b59aa4ef85f72d8694ea24df3f70759a5669f8f1ccf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96a0d0130e882d690e782b7113df12916d158e395d43dcc45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50e78b735ca3ed2818b8094d71248e4e477a9672f176184a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7690310184857afd135a43de1eb4865924a5c678bf1c80287;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9a01ebc3e2b05045a41d8abc775829d036f92c87f22ac731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8c15efa4ccfe517221126199b2bebbf3947f0802009afd24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habf3bfbb106d94e901d31d983735245442df6ba30e2ea1546;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c58152a5c6c3e8c0dd000e5bc71a873aa332ba7346a7312a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he02225a3af40484a509b2019eaa2920ee5c568016b3634ca5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88ea35d8bb9471687a489e120c1c0a4eb3e2bb0c3d4431285;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h603a3e5e2b5f1234c1e4d3b5c024274a52a721a5c7b32cb16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7e440e4559a1059a5da259568cca5b85ac48f781b2de829c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b635f12272b1cd4342727f286b6ad371d2ccdf1d267be9d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ecb7deed778cf0418656420f1cdecdde31856ded5b7220a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4de8c0c1df8983ea8c6403ebd397b981abadc2bf2647eeed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he668bb3e644595d57a58a35f237d8f19e2aa89e1521cfae0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1b4d3703a416509b86ecb184b839d28177a92f0b5600509a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ca61b4ba0a639fc9599a7bb8d7ba6d858b3963ac701ec8a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd5b2baa7257a24fef465957246f9dffbd87bc5746751a849;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c73e7d913d5224f828f0728a7f5ed13adec1b04c9e0e25d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10f54fb54a1d0c90ed39538c4cc00cecd7327ecb3f72b6de9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf94388e5e30de79a6cf55cd7d3448e5e6fa1c3f2b17a47fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h776dfb389c6e17fd9d91f0a7a9f737d9ce59154ea6efa6d48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h190f4335baf491b10c275529ad0d2a6131761eb764d3abc32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20f46be65f19c7cf315732d482cb3c767488557885e09401e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf387660ddadbb4aa093b9ce2331ce070894e60b1a660c9afd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdad0f26d7d2ac75756bc2a34e1cc12c2882a45451b222eda7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc073758129e5027f00b3ac15759036b530ac4eb754939da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9629fcd74a59f81630b7093fea45bf9935abc5684d01c657;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bc9a5b3d282d41f3285447d6a6038f074e35251957a8df5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdfd187b5be1cfdc93b4fa6be6ea7e7539cbdfe55ca815cb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c9c25e7377028db7216f24747681a85634cf0ebda0b18759;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0fbd36fb1e7daac3b4e3e960a2d46ef093c103d18d704f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6289b0c213f731fa90302fb3943f6f8a83db23bcd9f74ea3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95a90bf0b082995a7419fd58ce4c3ec233a99bcde69915468;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a56e90aab72abfff1919a2c731070120ce2a64e5353c82a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33fffb38bb2110ff18f6fff5914e641dba637ee7bb5e921d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f808e0d43f020ea4782ac93e723539b421ca880eb5891724;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he63cebe196098910815893c5ad1167632a4b608f94e2af0e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d616278dee7645cf73747297819a163ca080029dfebbd1af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6061116eabbdcbd4919768d79d9eaa8f9d4ae43a1563b3b6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae4d11bdfcf276585593caae345ad1c8b9565fa191c2203e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7e552706fcf71adddc5b37978be104301df69b6b76870f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h869c7f0a73c06df75a79957769f970fb869a1a9bc1d0b0fb1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60de0921b1ae44c28cc84a47d4c0b31f046e5bcc97c769b8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7add346e11afb1d878ebc09f47a79160ac4de1bd62a20fb4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4606e37df2da4a86c6ab89203d870cf47b9b030558016622e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45f5d23b0800f56027a7374284e06e044ad77cae9ec6c41f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8193c34be38b64a9177362b5934fb9cb3276c1fe31772c257;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35aabc53ec37984c7517d0d95b7dfadbd363e7ac423c8b84c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4fd3b2d5b96975b2acf1c2b5a3291ec40c0fac59a3d45fdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he18475f058ec6f5d625f7dde075c3fb398775edae91e9cd20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb562847458177e3a258b3fbb2c490088dace354548dff8ff6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he96c6880ccf3010d1d8055de6618f870155d0cc9e30e0233c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eef1e2c02c009a7caa97957a04fe116a9b9f664f5d45d070;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1195e64714da9b526686ca05ae5994c50f53b54b002b4c15d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2714e914e6ef8ad86458c2ee27611bed9b3cc0c8536962519;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae7659c03b4505bf89e92bda617e42b619f29134569568f4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a45dd4d67e274461d035f4c937fa29e176bb6ce73487693a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2db8be743a5698e3367dad9d5f2ba650235c00b8af6a868f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bed817bdcc2d1932ca010c2db12abc17915f33ee7bb7f4b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafa47d05f4900cb39f5be180c1f564ac80dcdbd1cffd2d9cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc356740708a67ce6c8aa6feeabeb248390e65041d1611ed5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b02abcfd891b042eb23b27bf09120f5a7246ce2712c41fe1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffca6f4aca9b18562661fd43fc573615269868308676f140c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96a6c06c022d7c7f13f7b033ef5fd34f72e1220cfd7c1b108;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6e10e10efc51370d4319c4a6ec47b98e20603553b0f9cdd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f0fd7d8044c56bec4ec1a6574dd84378e557872a0c4905ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0477e3b3face9c2ead1f7be4a75aa0d3d0951b1bbce83a1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99e695aff188049574479b34acbf04973b6a998fddc532718;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b7e52f8fb6fc18b795907a97edae76ca28fa4e9ea440ad99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b94cb018312dde19470b65400486b189a18b89474bd6538b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78af28feca037d2111a3a3d49e27c30a33d4fb92156bd83c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcba7e5c41d19ec98abc526c7210afd7dfb3c8c84ab7813507;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20a9add5f0f15861f203e699c117bbc964543fa6fab01998b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc56996c64612972059786be0349eb7ad607f5b49c6a31ba3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44e8b9e68931efe418272908f16a62a57c4163e19e65715f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28c8b83b9cc9bef266d2098b8a58d702c7ea33814c32a1de1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h634d6591efc46acd0911650c4478d64e23af5756efc945418;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcded0a02390575064aafec63b62cae0ffa76e78149827cda8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha56cf8635266d30405494726ce808e8c21b3f8a66bcea9d78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9682de4e586a6bb511a1d3fb56d5b8a0006f491f2b5d8515f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60ace43e8e3809548b0f7832d47e83a38289d8ea4de893e30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53dc97445d31630814edfd1bb0ee3aaafa63c4c1fd90baaa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9509e3b5d66103689c4d7e6ae196468995e2021df3cd93b5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c3d3731f4d7c6c9e06686a650018d299cfbc60f3d5da3064;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef9470e3f54099e7cd90b6ccfe0bd27bc984800125d832626;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79f30a8c4ceca6d2c84044eb04ade664d37827c8efcd3e559;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bbd91a71b827120b1994f6d86e76d84ae4cca451d8c63b69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5efdb80293e099bf83394caed3522e87163b7bd4802f05dc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16dd9502b7df716b6828fed2d063de375460e955e097c30bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7df0d5efda1e72ecd8d4d10d64b91b04117bc278b70d7b656;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h689328f625c30e5674da674aa6381736af57184599c4fb59d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd426a706d8c618243a4f044d116d66c21e16e1b462c9f85b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80946155c6edc51bdda0d95ec05d4462de8cb5eb7123b4622;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd92d0e7b824fe68e7c0bbbe20a77ef7c5b1ee2636b11b7d82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb5514744873eaddb968023666d630029b630ac17f81152bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he658d0a06ee6cd66e581f8cda4c6b134d9331e5fe690ec742;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fc20a6d44b0990b0f444dd03ebe63d8af55825b9c7274623;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3b807bbeac32bcdc08370f1dc84d978bd1fc8e74b6657f5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9d473f06e99db2d12d8301cd5526dc3ca36e5abcab9a8e3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h642f51b2e54c4fa65b14f126137453be0385f89884cf2c2b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebd998bb6b1748cb4a794b29bada64c2c8e568b4f7ddf3a57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5a79d61b3bb95e825de76e66df2c4c620b2dda1b8c945ef8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46ffb3c3ba567256989d71e91f0eb8660be3e2f7d7da626cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bc09ff7bbe6aa2047956ac3506a7fb59242393626a2867eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfc72cb0f7f3160ffc48a5c241baa60f85bab5e409e9227d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80f41f4ce52b1bdfc4a54512e15b17540833f2f498c937347;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9e334a77161a3905ab907c8f7b01c13d5b867aaa993971bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2461e4fe8271457b63f5d4d4c70e9825b3cd6a1f417ece738;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc621b7b8dcbea2904007f5ae1f9ef654ca68e73e5613f787;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbc9e35ba7a620f18298fbaffe442f0221e97dc7ee11511ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc91638b695d54a4f70099b3c32ab8accbd9f1187df04da9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3c80af5b0c10fcf4baa4b3bfb8dd1497089c027e8c5f07ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a1d723b8cc7c0934fc658176e42d696c6efc789e83895047;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15b385db7a74d4a11226c901ee6172c7e15eed6e58aa408a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he19390395026b3532814eced350710af294592483f0dcf678;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h237c1a84dd4507d20121b4b4bb8fbf1023e686dc2fdaf0ccd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3726c8309214ba1d570bba4423b57cbd42cbbc075f4bf5e91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b89714fb499c6707829d5c59c1ed15a09baf60e015a1cd24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bb4091f86ec9d6a8dd220fa945bf2a54f6247b0c5cab8452;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc305d570e62cecb442f54b0f91d4274fa20ac390f6f61384;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19468c7b27e464532c5d72beeada45a2f5f2fa0703f5aa162;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6735a55443764a2e6addac2909dd8f920944d175316d65e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc382497c4b16c8657bc8827faf8b1735a3b218b84cccc4ecc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc3bd28fd268c4185732c8bd29f9bc8b90c88a6c84d950a2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5640fecfee73ff4a6402183ab286625b9ffff6c1e1612d47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43ab53118aab700e4828d4e3366f01ab997e81239eadeef59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc40ab6c31f878329fb6c2352ae4e775e96d43d7a5a8ae469b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha14c8f22450ba8da3010266ddea68a6069c74d9b8a91e82ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cae02e4836fdc135c30eed60d2ddbaf5b2cca5ccbc39dace;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87020ba9085a7781ddffa8d73803d31abab4eddc5ed0d3b9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h992a0eefae8c52f6cf5b012d0e9c4973e608617a22247140c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3095017506de442b79f10a8972fc0ba328e6ef7be3ed385cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34bdc96605f658fc335ec4bdfdedb68216a9707921004b97e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha880272aa6b8ada6b0e63a30e718c8715d79e1e5a43888e17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dd96b6086049852f1d64bdafbe3a185bf4fdf1aa150607cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13b6a8a53bdfcdc28277bb4a47b3d4f1897e379879ab7e4d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bd870dc28bd3f460b53ccc5ab7fad52a418a898972af9fcf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc12b7d9c9933f53d3ab82b9fb778a3c66d50624edb655e36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf836e323358b1c1c52e1885d615d1ffc3230dfce2eecc78d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13abe7a3790c17cc5070dddfc12a20c042a7b4c93338d3a49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31e6d25c3396e36be1f944ba50e3ec28451cb0c9322cc07bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba5eceb77dbbd2386eeb77dda2fb1c683543dad16fa8bf3b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66ee508e707b9192ac2008a50edeb0135a1967bcf9d7eb696;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eb3835695e5c54e2a44701b0689f5f980d34da66eb635d7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdf77a6027d1d38563f9108c88b7cb8b572874bb3c787640d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ff60db2a9735752d7c24713a8fa4c8d7094e965309db57f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fcbc42afa5afbe8e72378554746ae06544cb37787b93e6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b8510c6201416c0267ed1588df4f5239bf57b43272a79a4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8a3e560f9e6ac249270f274068f84544d62357742f77450;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ed9ca96a946963e85ec5ecf5f0cf68108393096d2d2b4c32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9990ede8e2e67c013dfd48e6e7616c57f5f3f44b7e2f4fcbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f1000864e2365a7b29c6070aa258f1a422998e1f1d28ee38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc95b6d7bde7f7d24c64f324b73091d2c70befa31fbe3381da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc90720d88c7f99f8bf5602c57730e6489c828622a96eb649a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c0fe8e20973ef5752946182544baa3e767bacc7839088169;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h939a8a9e2067890d2ac8d164d328eb3c766489d6c3e7eaff3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb22056d0187ebfb537eaa5141664b21f87fed6b2f11121cce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84392cb4cfc1793b19cc4d4a4bddaf5dc5cd5f77bd0d82326;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4ce37ec80e9389e33f04783bab765d7027353910a2ecdb61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6abd0a75cc5612e09c04c2bf4e9cf1eb7540671cf6ffa2d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h982d7c9f466dce01f0c4f7294e85db128f159e3e7966933b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb558b5e295d86c1e1f7f9c3d2de0622b79f36d604dc573d6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5594e96579b5ba052854a1494f14ed078cfd8edcfdd794880;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6447af438862febb3c4a189235058abdb13437aa5bf480e92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha11b3d8cf22bb0b10e1fad51e7be4c53e499c037aa8cb1047;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9915ba5ac4ed52fc6ff3236301d4f8b16d7f04e04ec6eb9cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1b8847816d4c07db979daaa2b2138474070926bb0c046842;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h433d6fbd142741fd92e4ab99941601f31731d333e241e17af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9123496deaf769a472ab594716cd51d726fdf1c5886ec69e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h518c03b84b20c6036c6e2771ac677584f415cbbfae64748b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ff57bb27df1349a7f81d2df0bcb70721d9a20a6cc0764aa5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86ae46520d8e1c37cdb8be48a208c096200bd6c97ac59d3d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70c1d26aedd5eb5a99f767a358936092f2bc84fd7c9cff891;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3368bd54bfe9737cee3f33246cc96466878bbad8ac56ecbfc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf8912b7caa309ff3234cbb4b2e853f9ccc49158a0707887d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3be8ff5accb973d468bdeb765ef4bad8487c02f717d155519;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h484bbd546f9fdec59a9e602b9e3ab4f6c5cca718cad9b089f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb8c5fd1999a48a729a2e080ffaf0ecc2bde06661a5bcdcd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h411fec30a964d9db618e6bee2c226da7fa83b716c360b5d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a04150bf9e06e33c37ae46fdb7ec078fa6d56f505db66426;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h452f5d64022ba52dffe7f41c8937073701a8918b6d75adfd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf843aa6fa25ea303e938024c99f07cd6ff5705630247eafbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70fa3037c3154a4fbaf0be1aedad160e13c296e739054e3d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25f5ed00ce625d907a8159107436fd782ab932985f6d907f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7e32952d975d34d7bfed03241d4895ef19ba078ac11ba685;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d86c23cfc6948417b5426f05dd26cb730e12c4a5e55c6f7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3b6175430fab642285dbe1a406b9d20d8ba5db1e341c9cc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89eac6b12eeea6bfc8f04f2453804e1253fd9019101e1517e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccc9c47138f2d48aa078c2916025140200ecf73adc3dd75d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba651fc13ba896fe24e947d75bdaa526c581006c6bd7716ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80ad4b6bbfde4747c7850ad60200c3a24a261db11d47635d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbfeb5cf669ed5116962d4f03bdf309efad0e5841a9e7efc6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c420474a5353b14bdb15de85cf9b290b183581dfac6c93ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h449fc6b985b519160e542eb43c895368b58578bc336b8038f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fcce27a05cbfaecdd830b1bff287f4738e65f54e289ba441;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea119ea06b6c6d9d303760f5c4a8188c025d1eea068e13047;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5057be8a3fa00f038261f3905a1511191b68fe57d1f6d43ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf86c87ab7b0a417a3b7c93dd8b015318bb03986e75aa5b9e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56e0dd8d456b51d6fc2883c1cb6c9647ace7535901adf760a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a4ed39bfd3a8308ea3f9cef04fa4432ad64323c0aca0e4be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e79cfe569f9c67ef3560898267cf24136baaf17d51a3fe8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h364602639c8b82a692d62a696a8186cdc531da04b50338854;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6235a7287aa406d8de960ff9d1239948fa7dba21029d6449a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8aeeb043a5030c0494535ae924b489d136b153996c497491;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h738374fa2524bce043c883bd353b59e2255558595e650f2f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bfd8259ea9333d996a268a6750c24e6ff54f68929f8c37e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57834cf8890d17ab22a59aa3184f628ee42941a4186ce6753;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb668804151db14fb29d5c7f26a214d3f57cc0195ddae4f13a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bdd1c8edf8dc71044729f8be9eb2c435ac42712fba8afa1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf2a8f15f04756c2bc2daf3d1fa95ddb53c445b44108aef66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf45241382910791f4d750b05925b23df5d474bc4859a5f054;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he16c50faceab8cb664a2a781ed203aa9e2e22f70c3d1f7742;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde0d3af8b6fae80544921881226c060e7b402d4e264f5549e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7715de434a924005420ed3dc3b4263dca80cbd15694e0d1e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h179ff9a1a2218c91121ddee18ff0bcd4b2d400742490ac7f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6009b6268239e2c295431d1bb512ac2579a5eb038db2ff3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb1514a05b9bb0b0eecac900e320b4cb1b801ffdefd306789;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5ebaec31f0934df4deeb4ff3748a7ffb4a42e6a4b9778ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f629137e9431f2c1b54feec386f96ccde2c74424f83457c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4e85e5d806a963727c19d259af41f0e498040c93c0f903d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d166a74a5522e983252bcb71b3c82ca62e56f5b9f3799504;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0c5ed5ea11b889b5dd5a9923d4926194736efd976f52fa45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d3fee43a1dd1f2444842421857f191544f7ff34db9751703;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b0d561a76279e2684066f17147b2b2a0288e6f8bc0232834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h956f5672543003c60df626cd3665e3a2539602e68860f3efa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h298c4bdf71f203be46e1158a1b9db6b94c074f7162e2ff4b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdca79140e5c20f35e0a7411a2facbdf93b779398df11ae40f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98e4195eb8a391a1466cc1992f40bb2f37de5da7e2e7227c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c14e09bba3e589c8f47caa7828ec0dedecee78b7fc613867;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75797db18d867764c89a2ab5e95a5d8d3736c7184ecdbf9f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0df1abb42678cc6924e9b8c815ccdca007fa014a2b72500b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7563ca558e860f1e4f55a7300ca7ce67f0c45728d76cdd2ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h899993ae98c91fa1583b7003dddb30a8e8aefc33bc0569d11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6d71595b28112a98757deb89323207ba7d82a16b9676f984;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11bf25d8d13b70d3f828adb234782df2ffda66b5669ec18f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c8dd4a6e3b75e5bfbbce757b98f78214e6ae60f85e71b346;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d6779165dd40bcf8eb11099ed479a3999327a91063afc10c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h431cc788b7139870b9e00ffc717a54286bbdd4d6ab859db85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd91a06d071abfad162a4dd86fc60179c5c90fe14fe5c64313;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb44916d1425879151fe3c8070a0945953198cf621dcc50bf0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3216893b5a17f84dcb75ce932706b87d02bfd938073976594;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7567f289f415c42ca432c2e69271b5c4a986dd4e794382795;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h140412dea809003ee33494491b5f0808872252a14c0344c6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ef58d071ef44540c48a30514db30294f95e479ea6a55c4f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46e51fdc7fd3a86d236af039661ef94852f60b59575a9555;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb215506e7aa6efa643a1e89ba6cfc48275552e26d2be5be77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b1e00a8a4c5e7d06062b0115ca2c151872b6954cd26315c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb8b5cde6039af3df532eb688bc81db8d2ffc26494da2418e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab567fe48e48a23b909d2b703bd3fcf27011baffb6d092155;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h999e00837b37bb721661e42d5695a52c5880fce70811fc374;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea82f925564dfa65cc3af91b0fd0c1fd771eb013f2a1db759;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd170a696c2d1939e2433381b62308431b0cf8fdc78eecbee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf79b3ecbd086f9f0feac9b388a4e410958233dff7a86c0277;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h713cf453ca013d85d9067d54e7f5ae484558e801abcd9505d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25585de7eb1f39c84baf1650f72d93fb530a545613171b897;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f662c71f0b2b77e850222e437acd8bedc412d0aba19c1d20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21780d614c2a12166cd7799cd5a7f79ca754e444e1f9d20e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e2097cec876b468e12208c570e3d92325618c851ee7fed64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd677e880de6b3c12fd745332caf46a81e8779f57b54095efd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2bcc1d030941c054dceed775919633dc84d0b480b861b645;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had6118201bf25ba9ce20e2326758271812c69b1518c2183b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h546dc14704a6fd604fadc735f02c6c9c14d6234fe27c82764;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ed7d777df37605cf1a963d923d83a32f8801e53e92444aff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92478c43fd7c721a012e7263a7c8286c38b8fe2d00f8f994b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ad9f1cf3ab0f2234560955a18df546245b90b7366f72d474;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a8ae716debb9b6c071b3e78a23af12eb3dd7e703a5a3d68b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ef3867e6ce8e850fabbe7a418ad08d58c889cf5631e08ec7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h889e4ac9dba56b645df0b7bf1e7ad8eca3ba7ca1ca3f69da5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h857c0968855212766ed9dc33fdaf587dcb32cefc9b9287538;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3a3a7b08620c768332ff104ac77baefd4854d099e1edcb8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcec642ef5b99f2946d80e386a03f160e018042c92c4d2701;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf439df2b232fe7ccc488433502614c595d5b736af65cf44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4b82cadd9e447f7b9ac441916f95f838d1780d8b87c2a5c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa60277f866b0aac329b58913cb82d8bbb6f8e25669602fac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cad48da1e5d5ca3c546a72e79f9a101ce22e01e8bda387b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5a9a007f6a5c2b04fd88e49757470d1598117727a3bf18f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5fdfded9bcde8462f2eb6fc8e41d306b0ce16117bf04d315;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7e6f7a749f8d7e6e0ee6c7ff2c2af0292ffd6cf81bd571d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6725e5cc4b112195b66dc64afd262e775455c244426f01ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42764a8d7fe9352b50b59c14d2f4f76814008cd27902d57b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3225283b1a9bd7320bbb62c68699666242b21a9d5f3d7d32d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33d1d607d3364dab2b3cc358184a1e7609c877fea768ca4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he701075a573a3215a9c1aa58f273cef77a4e307e637a0c508;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5db2dde05f239b7b92daf6c30d651c638c503434f0ea65beb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89cfe2e0ace27c50c44347cb7031d2365d05b53f8a2237b0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1686b92fcf98a4d7281adc0eff1bed6c34014019c21c04f48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34716187a26db77cc6c2ebdb5ec0ab0e7702f81e06d0e440;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3524319753a883e7a3b749a241d8ae989a6974ad3d439d4b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3be9536f7fa9bebff704720d47c6571fe8dc2327631723aaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8259c8a9ee85c3abce0dc2e24dd573a581b762aed75e7352;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha097a17d4b3eb3ce944b09cdcf85e0e98bc8ae9abbf925ec7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h636b340312b641ffca7f535f6b4c6e185392c239ea9a4919a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62c29698f3222b4b6da58d11295f9aee0321e9ed1b056a93a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ed1b4054fa928d0bc423022dd5773775800ffa54073f0dd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85209710b02cdc6feaa8939b5c47bf4ec2d47b15402bc389b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a5e9d563b0d3f8181c2f50153e925483440fd2d60d8e9fae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc099446271e1140d31e6af414472d77acc19507f6892f86c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f1cbdb6d195248f65ba7ead02e9c0085ab44a955a70712c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha32b383833a468e8fa46d5cbc9e3e1695229eb4b439e4677e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h722d457f8851904171996ca57d14746126468a1568a50d522;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb80caa1e9f3cce7d18b7bf87945c03fbd32acb0953a1f4cb2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbadddfdb2860019d178d0127ba2184dfa35e307fc2fa4d672;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cf7ee3cb172f980498670c7005ea424fda3451cb445931c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31624d91940987e22a06271ddc2a205288be895b770eae7d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he611763a07050a4cf0d9e0214af5846de05360898e8f8a5c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1afb330e0c97db824fe41132bc29f7724a35a31c9d12916dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87e034cb35827ad87b15438defa9ae5456e95706e812f16fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54ae06a7bf557081c99f777ccd761efd1157d8458f4f877cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24b10593cb8cc767f1764aed7fb6c4a1ffe7f32be8c52a819;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2440c650e853989eaa4cf4fc076db7fe9a0eb6e658d29eda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90260d91f1d8a9c23a598df1a3a35b8a34a6c7fcdd471e0c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aa4569c7b991f6d758548aa892aa86649a0bff4fd63d2747;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76536435b76dda0643e50b9e06a7d47579b3c855b34a39aac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h232c8c40ada1a7f86c2a0eea20826be74fb3dab3f9794674e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e936744a1e49c51fd98a025328361d36ec0730e03135a549;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h422a46de3b061b01a5ca3bfb09d89d6ed18cd395dbbdb0904;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42e7bcb6204d0f7f7757d8500989df2c804abfbb93776a3a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52b50fcea85775567b34c404ab8e11467d066321163c72ef4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb317dede97777eea68020c62a7ae60c1f6a06be6410632731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb2f0e50179e3adf893eae646e59a9240f067addb928869b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b14e9ddc8986eeae848e9d1a37bf24ca5239d4de9b87444;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78c2f0a463863cf5bcdb6ed0a564a1473605c413bcbc64e29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h935e10b42d8aa6eef3831318db80b58ccb9fb0dd22a653b05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b64007a98e53b9e7eb4d0b207587672e6af422931090a8ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ada4b9c3ad9e71d075e887d740d5525c51b6b5c1076dd97f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h156e405fa217647a3472983bea07d4a80a166ab19a8d680e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd503e2a93c739199888800479b2a1928ad4d5ae8cca5eaa81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fb14f01b2ccc829445c593141be726e532be4eb18fcce5d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82b11315e8ca60cef5d6c7c2b67bb34b957f6266e4b96ce87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf404cad8060939df91b685e94be2cc4c312c60ed6d662ae91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb76481b8a6c62448cf79fb4bd70f58ecafc91a373ea0ae716;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h140f7f9f706ca8a146b4e2017c8e216cb8c7043752aa4b56f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12b14925911b57ab31ef366fbb469283cdd6399088707bcc0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e7a6604b3f284c6e5f0663d5408a9083c3f2f84180b91706;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b4643503eb7f296d46ec9d71d7113df3bd6a524d58302fe3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcf1ca0556c0ba342c314d6d4c7c4873ee9548922e009d9f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc34aa77cc580b2d479bbb0ea4be072020bafd531b5898c6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1a005e5b3c900ca845702e1b8257989a9558240b15bbd6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he17467ad901726b4297897e2ccf03556f4871f1bd6185bd92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5971052eef589c23a0ac048eccd05130844211a2e8eec91d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h743b5b7b1a5b4d89959112d29751cbc53e096ef9b180ecea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1aeb25b75816f8cfc17f6cf56dd720b85c74bf494ddcc667;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0d76f805450ea763f63779482fc67393aad291fc5ab85c4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61bb7031d9fb8630acc8eafed7aea2d02d9f2507c90e6e70a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66a3a5107b206b628591aad5a67e5c4ba9ec893843241f27e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bc0f118f75a8bbb0897cd49cd1e27a951afe2d326130195f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b9ea6d0fc50895b2a2f8e47cc059f96333fa66c976449341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b02aff7d2a867c8d68eb3a683e3e93763fa3fe82cf234cde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h457ce959838ee131d77fb64525863de5d8b6cb08abf410dca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74a72e129753d576079443792988b859ccb4c36b7f34f6241;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h229fdac3d235cd59fa296ca9e110461350fdfc499c5301c93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93937fb21ec8994925c4779fdb8ad0f81d45c817036193f47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc432a3bb82ac55f5bd97b10310c59b04e54d9c518758a0ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h612abb1222d38886f974bb181e34a01ff5bb21f13dfdc1447;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b2fcdc25da48c766d0bed063d0ee98bf7c697725efbf2cf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd952218c3efdbca19bf1145e078ffc4b1eb18192fa98f7832;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a0c13c09c587f2873c9d04fd1438ec6e1b7eb5808b0145a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f0aa2faa7dcfc65a8d58d93cdb08aee5a115e48fbc1b5853;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ef578d424a05c3e3d504228e9681b87087105a9d611bd555;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h691cfcacb9e301cd6f82d4b6cbc225b15ffde048adc214a7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4590fe50902d39c976878bb6f6b428fff845c46ab8f953c15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb707bed8a6031fd0d19f55c979163105742465e2223ae195f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdb2972f351652fac94b9c5276571e77c1e9552ebaa118037;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba395250146a1938a0335ec80163fe42b6c506958468fd0e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e3c10f6bb9f2e40138e3db9594156801e2d17c57e815a7bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a16a932977656751da14796a060a0888d1751a5f64f2678c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h801923a3cf92a4713fd6d25bd478f709389d3e897c85f2998;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he00eec14f1c1d6340650b122f2d3443bfb06929984c421eba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdea5b2952a89380e82bf9c32f0a4c337b334c463a762bf3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae4f8348b7f7f34ed055c8a438cca3b504bd4e19975ce5d47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha804104cada1f0639f619f149f9b5623fb5674a9f9cd6866d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10301fd28ab457e219e44c440a17712d6439a8962751c3f27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83f7572104a0447362d173eeb8525a62c0d4cdcad5a5f8461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2268772e58c93bf23c2f83a1a9f68dc6a834a8c08350893d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95b83db97a8b166fb648f3e18a579d0a5f8023dd3bc8121a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11a82baf8b24eb0856aeb35a8e7d1dc7f1b125af3f3cf0923;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1749203fdb9a6a4e1239ff84a4c9af36137791b64ee1b4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h731390af4c82c4b8ef7b3c293009a3cda1cde2c88dee4975;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90355bd6ab4f24f86c58a98deb705bd1f3bee40376d4488df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fec2a6eee93d65d11a6203c1a2dbf494a0ed755844224a8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc226e3089b5214c26bc2f04de2f34674d0e8e8f535db377e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21346807a490e31ab203ecc0b50cddcc5fd85e764ac6acf9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h717a1d35a9a139d3ad5c810b5ba2b10df6508a742e7fb553f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc825a4f0a5c2792f100b377144d369bc577afbed770dab0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h650189fc4cbe2f30242136465a4ee2459eab131e07670e993;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38ca2d57e4091e8b337556eab0acc01fce4e13d2f036ed35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc317a2d7952d4d76b3158ba3d6d8bee327bf9b50f6781f9ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff85da4a37c5a0bc7c4dfb928b038b9d3e4c32815d163d7a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h236a9f0cdc64a8dcee13c91199dfcb2c64b0484f0f0439c49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb52891bbfe1c22cb2a24f1df2b9134057aaa18ce2df12d0fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14387ba3525212bf65ee5473cd8f54701b7b7f3a8e2bcba7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d0c6a94fb1a6374d8c06164ededfa1e20f32667340f05835;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he51325a500a1844ead1261a66c9edc74ea7445df4ec67fc53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9aa24b3fcc440a784e478e0706244ff38a50706dc0be4c7b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h109588007fe3165f3ff228a3a893ede936b90bcf159b3bfcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4831eeff1c3dc07df5aac2d18a621f08ac395ca486611cf3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bf4122acbe2cd8ba27fea945b637956d592948385b07d5cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha45141afa3014c0937b1a3a85d552a3282017cbe60351fa68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0df18f24adea55fe8ec399ac665601395132fd22ae03f2f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5e3072f831bc8b84573e69bedf24fadceb0cc7cf99964efd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26cc525d31676cf901865b10e3d9bb79c22636dd3721d5379;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h971a0fa1db081b6fedc0ca74b4be97c2fc5a8d299447e8aaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e8c97caf2cbdf9c645d0cffef6ca0a744130fbdb986089b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37ecf4a7070615b6c771e01ca0283e24e4769fa80a57a376e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79b8d6d5defeac1ad6e10ea6c0ecf5ae6894767e473317e3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3025dc2c1480a8f11770e4a07e5ee6201433129a1839436;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2b0d5d5c7e1ddc379bf073fd6914736ea102ddc0b61e11ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71dce9cbbf10ab10324abfcef59591790419584f53105f8ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7656cde6d80adb5f9991aed8452edbe740ea2a011fbbe714b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78f495e025e252605f61ebb5d8e7f2bb4a3540c51bf3f8b9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20fc7d034ebc02aff26e074830151f39a947d963283368975;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h476abc5a7bf4c191cadc1d89c59f84a989b6046c9529e4aaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h821ac907eb43325ee572de2c1128356d4697237e9bcfb5b8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h877742c2c244da514780734491674ce74b7144dd5047de07c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11dc30f428aa3c7cfab1de2820b96e86b2b4da7430ed957f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5e250e6b90f582c1e31ecc3caefe0e8de9906acf1f8b77a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5681db4c5a80cf4f2ad5725a245eef817cf95de60eb377df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae3a15cc869a3abaf8ad15fc9d67b64ab74ecd71317b816de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebc53b2b5fed28e7e8e8facfcb53f68d49a5185f9580d8a11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0747be7588b86509aa0523df5a971f01c31af0272a799c3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he985344cc082347402b8561d452157744e4c4242439d157a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc06ef792cf4dc42fbba8aeaf233b3b1b9a1b6938b6f0e5ad7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f9acc1740c1e89479d0b5b15ae7f4eba354b5916a4460449;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf15d22e690fc8f9ae5775b9a9bcf83d1e7675c8bc2696cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36b8e4db98957c6f5ab7e41701a47f74c3686ef7d6e75e6f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d0b5eb4525ae76d6747e36fb84b87c60973f65345ee8e03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h696ed3c4f6e153724a00ad5bdc5568a130f64d32494b48d6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c04d83bf1c0e0dcd1300946f3872be48dfa34d839bd3c2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d2b0259a1d2327cea9fbb8dc7b11009949a857fbccbeda7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6960eb3a826d86be7ec492294027f91be14844d45dc3c6eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9493a4d5d182aed27bb0f1ea0fff9d5918fca28a5cabc112c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dfd20dd5a46f665a991cc44504a2ab058fa94456ae459fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eac92a6d938679e66b8980c431e97e56a83e38f98764948a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0a1b93de64e6c8bc64a984d960ae42783dafb777382dec71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h612a324ab5b56d029a81937673d0721e3b27c81fff168f00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1006c2731bccd2260814202d8cede7a988ec9ffa707d8949;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f2a121d8c29aef700e756a89cc4cb66c4247cec9645c0a37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7afb6e49d035e083e1a5cd39bed696028166a6d9c65a75e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4078772ce805abaa6ce9202bf5f277e2841b74e1b2b433481;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3b444a7f8c79626888f0f20a504aeba671aca0572f17ebfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c97e216e77f9bf79f9094f66e6c7356dbf9a5aafbd490dd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h948a55c717b9bd2e7d6ca03f5a5af732c657f61de66dcfc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h479fb6864b78ce87cbe0bbcf48abd0a326854c0c362967c47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fdc07af315bfd5da52913858e96dfa474ab05c9dffc9df6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72d8acf31d3121490eb5db9ec6a35b99644ab298124cf3604;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1020c8b35157c162609656b9aad1d36e338805f22f27ca2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8526b979157ed13a1c9742ca60bcb5b5e97d75ffe14f8dc85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b5d6d54e390104d48ca82432e3686e6581b920bce11b7fec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a364b0f12ddd1fd3ed0b81455f2283103494898cf231f3e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb835b600421f207801d310e81967c380d7b10ab189b47ddb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b47993d95a070c440c780243cdc6e8fc7bfa03952f7e2d08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h218cd4a296cf508495fabeae6344872fda92aa95ac28f2925;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5026d05fdb553a241460a7708ea18932de349e5924de4f31b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16d0bc534a9de0f3e27255e3400cfb3369f54b181dfe65643;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1107646a27e0d76d0b6c8b430f7bfa847e4239644988abde3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65971b0e975a2461cd789509a3688052a459abaed278580d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d1bfc88055e8506073d93d3b924057ab0356c0d8e85bb1f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30c3c31e5b66937bb67d176ae2056e5961d50fd72496dda28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h575fe6c3cbea77883608a0ca2b3c9a8cceaad9979dc3e8dba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dca39af59fb8b39ba5a3966e0789cf826590f54a0b427f42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5649f074f55bb71c7e0f0b6ee926f66f33d62bfbb06ee99c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fa617436cf185711f62857509d3ee5ecd28e59f4520b4da6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32a1638bf4f1d417bc1dfdfe295bd416576536285506468cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fdbc98ed790022bf82bfcd7931125d0b74259b6a30002c0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b265718423433dde45c685c925d30cf4bd42c77471050c7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d160e4c611de0d391f346211b2bb48106f70668ad8f9ae70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4af009ac3b4401d34a274d780f042697278a64f61110ff226;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafee16a4ad0312ef7a7f6779ded0bf1eefff893199d0b60b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h851d76826673361b98ff8a0a5c0f7bb8f171c00dc017fc43a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c29f5925d79a091144467be058b4b26954a055b02e694fd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaf980d68283bfa43c98b86fcaaae930431b392d0f2b1059f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h613e477fa1d1fd65dc3eb3d8845aa679f354dffc8e40833b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d54c158de6757aec7a16a851b8fd68208b35c09e5316a3a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66203ccbaa8cf254d6958439b40b089a6e624113b3bb1935d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d358dda58b09e6b144608b3a88336dacb727289fbab64ed9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd52c6f1b448e5dc47a99334a30f6a8a0b40d113658dcece41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76453dcddc346944b768777bf836c1dc35175b07d910a519f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb23614d2715d65eaae1eabdd7f3b0352005c70c498990f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe5ac2d27bbbc4d37591720a376bb513979684a645fafe97c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23f63739f34a2ceae8c3f68ccc0da819cd5f382106f7e6cb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h419f232c01ca6bf1cfc286b30a6ed6f872be6f1a143987ce0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h458a571c406c31376d4494470217cdd3079b6a357ca95b26e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53728b509d8f331b94beb7462f19cc5f053f4ac3702495793;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h802ef827c023c07ef90ba06457087c389b7d5dcdd921c09e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1f7abd4ad5ef49425bf83153c74cd0076942cc661fac2775;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c4d585dbf867e617c6762e8bccd14059e19a1fa8a30ff812;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefef95b8567f3976cccd188478e8d7323819994f2d16a3113;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3384b47bbf1fbc016b0b0adfe11f03108e5bef3f685d66d97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa8020de4ffa47a5bedb3d27ef0e8812831304c117d294220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d87f3064baf5375a45552a28642dd6fec4cacd715556649a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfefcfb07b5a853914233df7bf571c3b72f4e538678b5b1f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d17aef17b1f6869cf29a5c3de518efc754093b9f7f514013;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0a1904c0abfddc534f189550310460eaaee061f727c41e60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7c926bc9f59730280b6d6f5d801ad9b8679045a83765abbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24a06d2083776d512b766ac5bbde4a661758dc4c9a6d6c348;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61d4e3118eeac3a78c9daa9172de6683e792b13e5bca5fc5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96f6923e7fd783a9d6ddef4380f3e7af842df0f0095ec7aae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2106fd04d3d492525a75f7cb9f3ec262d2967892ba2f7512;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha90915b05eca62a46aba2bc1283444530e7db444ff0b9e02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc75a452891762c64f2bc4628a5028560b6303d3d42a30b919;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf42a81c017f7dafe23b959a379631d81f9a78dd4cf2c72831;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31c32ad7385a39e055c9e92a954a70ee68f21b25e2a0196b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8ffbead4694caf9c78191748cfa47f4e61737f9bbe5a55e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49ca8ca4a87a54429f0efc645df3bf2c5854f5b8c8852e60d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96929ad1efead3c02356567b0d654c5f221de89c94520b396;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eedfc9fff7d8433a8197fc876d63cdd01f65c2ce75f038e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65e195e28438120a46c9fa56076f86d55bf9012de65bce8b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haff1ab8526b4105868f3cad090c3f525d9697726133a3cc09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he49d91dd06c50d72555b48e77b2205cf70a5bae33bc25b9ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7f7ef823b14f84249dfdcc974b90374e5fa6cbc5b4bf1d08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51374d839500f3936bf4b4ccf6651f61625be4b8571fd9f2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89a0116098071d8775ac9ca1eb953b4bdf509d742a4e04746;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf33ae7ec73a1f4a8647bb602332fc44db846887410f712c23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf2d52212ab0f98a26812fdc464ff5fc46df6906c7f627ef1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e96f2e4249f2293d0cd203b06bb6d30adf65db59e34791a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3573d138349374a94927fc85308b7d38276cc9383082b523;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf59d4541ee40c618c71b4d988ef1555fc768ee9cf50099f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36e8995ed459dd893fe2f237e40f78f7bf955aedcb1879510;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90a22adc6ce3e68cc0a856a440699127de7f94006301a0764;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70e8b7eca5515f7fda576ebf3fb74e7b193602ee46e698988;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h584e465664cb98dfce68b40da4c6cfef44f9a8943b3b71375;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h329161fa39900ed8a6069b851fbfc5b0fe25fba2cda5f5428;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33c8fdaabbfe073be93293d377c9187acb4c9d0f275408faa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c8156cc3385d51c7a8bff2631826dc2545bbdbff639131f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4ecc9f03782350d64d62d0ef043ff9110abb45236ca58ed1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc79b59cca0569a85572bb3cc174f5730c6741e0d2e88483da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15bc30f93c3ce2bf07513c530bc71d44622b576bab28be137;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc5cbc0e3f218169b5472945f11c6ca7b40ca8c7314e066f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed66e1e2be7632c3122f891d58548084fc8a871cc58846f17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91fdf9164dd5c6687e99c757c3370233a0536f485349b9661;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h676b00b9d8be700b10308f71c01afbd7727cce261d64e671f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98dee72b7e4b46f20d0d14b675d7a807846e10d24630aa307;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a53a8850e8a2a41ee9fb15c3f8cbfbb1d7ea2308fadf3323;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h450cc5d954221cccdca9bd7f17f6e9e3fdab32c851e1247ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4597826f8fdff04b9c65144475dcdb17a408ca259fc08ae4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h391d7924cf5cf482e358be880751649ae29fd099c4b14ff5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0a1d2157676b70251c0623ada6765e3082e388b73159f082;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha236c83fb193e6db64e8164dc55601f9fb722c607d33eabeb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1bab198fe8d55ee400d1a42d0062d2ae2013000cb699f8b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdcfdc089909ce81be8543341fa8bdb2828e5d3235c3657ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h627d4329d16c7cbd1d28d2d9d43b06ac2cb175da074aafe49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dabe8617a659195ee557d2a959d764eff83bd79867e562d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb243c4fe043bf06c04f5c66c5e764023e7493dd6a85b786f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdaafb7eaea9ea1cb3bd8438aba62a858e644f090dfa4d71bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc77620387b061cfb440d63601d4e93eda8903afac1a6ffad6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7180f57b3cd9b3e97c1ba966e5e1ee5b2c68d206801aa863;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69937bdc895a551d2f60b5edbdf8a64cb07703c901abd5537;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd17011c50c2db3ea1da57a821d698ba64d6dd878429f752f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a84a7f988c6b4b4b61c5ffdc60aa1d7917c8d302e3355d16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heba88c8f083caa16a1215a9509133eecb15d6eac1beacc6de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6cce2a98cb16bcbd6d2cb4a976ef398f5950e1de0970a1b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70a30b9fcfa6436a4bd7e9cb313b71336aa7d9ea677a10b32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8efdfad79b1207eaee431be0026c43aaaf5a0a3549175e952;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b97cd2531b1ea6b54f7a75ded7fecef9e676534055e69d6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe857c6357fe36dcd4e19cad10f76586b55939b756fddb5a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c103db5c8062fa5ae300055d6a1ac670f9b0b86758f00b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33bfa60d44a8dfff813061a0eeb81091f97c8faef2838d518;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ef5317dccd9108c37cfb8d530f9c0e6fd06f15f8063cca8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c48d28609c7821d7d29e1e52be03f592a1825c0512d28b63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha67c0bf4bb3819f68981cfd38813325ecdef5cdd215d49fbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5bd7fb71ebcbbfd1ad6ac835b1d91c7f4f3c87c064a67396;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1e3e1b21fef3416edce408432a460632798951bfb0a078e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hece53b2879d387c6ee7b458579266211c540eb1ed22a2a065;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87cee3afb3c019a84d7ab63b1f1b4c6f6a41eec5c9d0cb2e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h436812f0d0c5affdc3cd5ffad17fb38cc3784dd79bd5e6881;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9bb95599a326cbab5dc2a583439ec3258fde52c1379409c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95b47b2f9dafaab8e083e434d77225880a7fcbbc72484e10f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h412fe182e869e0b2a596b4c7b4563c6b429c61d0e06e82c4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1cc6ecf001114d0bfb198a714bf08ab8ac7305284b02589b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17eb01c72cccae05f048cbabe6f416e89650e8f04c45b4b57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcec0893d65d1f02865c3dacd0155c8121f2261f22aa40ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f480092af3194ddbf6d0d209cfc0f060180ed20094601acc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb11f4fe61543431f321477c67b0e81315544e03d9af1b40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f6670d3b223264e12d03aa2800bc7e7b748c92572ecd5c1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6093f119c249b2b00732587a2e03a218e70f1f9919e1a8352;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb7ddcf0bf9497a84f86716ca9cc655ea53c9703261336bc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h510ad41b26e30d4edfdb16ae6c6022fcb4ac56dd3ca518222;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14da0dd6e27febace5e7ceb2c66203805654e728775dd8b7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7585c8374abcb94c52c6dd6504eec3f9507cb3007594cc536;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b876ca4075e827269d3792d444c9e6cb0d327492212ebb7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1341bf62764f156827600ccb31f8524d278ff4bb01c2af8bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f48fcd8e61ed55dcf93bf97a600a1345f5bb7b6269f03e12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f96856dae3e6efccf40266fea149df24455883a1a6e3d582;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a7960e6ae4573dc0e8638280a924038817e84376629a3a54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59bb98ac7f090da3cf24ce5a46e2e3e3433caee8cf03baf73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab8dfae58e6c69667bb4b13f45ce5b84b93686a2463131516;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d8fb2b3a6926759d604456e89c348a5c0f04272c70f41e5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17d436f559a967ff230a12b2324ef9dc8959a5ef3b2d64ec9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd82fc34adac022fb4b3c10d636a5fa46b94df5f07ac49219c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf911e63518d8fd8ebfbc89b8a5f14026c8e579284905e21dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d1723716b8b47a22711fda797d571b3bf69ea5a4e40e1755;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5be5691b3edf61a696dfc320152eee3f5d2ef1b5acc0ebba7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h276e2707bc77132ce7e9af8cbd8391cacb9ef74d11a6c2a5e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3206b66f7aaf663385371c65286f068222610494c394a50cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90e9978e51a3b726c1c0e3971faa1f3e740e0bdcc74dd1aae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b70733d9356ee4e2dd226aad6e95905147f98be0b7cc1dd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf35c7f2cae44326cf3130cd8a6bfad228962481a075d49f42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b4ae981c59c342a539ee01b8454c7f038f36dae8fe5af401;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf79101dfcfb326b2003fc20571ff3d4cc3e8f0adb4e868814;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb7fafbb8aba7c36f0d99cce0dfd25bcb4a44764eb1f238a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6836f4bff8a242d860ef3dd2c4671f32ae4bc0a626a07830f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h879c7c37ccb64ba830a408183cef79f1d1ba716c7c7c9d492;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha493819755079ea39463a95482788f58164638f84bcba38b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf99d3028261786689c3c61b7f4fa0073bbe258988ddcc13a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he85f3eecdd98a6c043e72475f2bf94b9d82ab5b71ec750f81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1819c478752f972a24ab00953d616e4bcb9e65ebcbbfa0c69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h422a9704a3e0f4201dd640d0e57a4d245b238a2ea29f67402;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ed6b52b3a5f23d32e2862a21a34cc0e2116e2245554f73c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd78da0519998b64b0c1b56172f706ba83d75954dfadbf2c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf1a59b44bb36e7da7f4d59496a717095ca45e18dbcc2803f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e2ce7684910693f7cd673586d3cb722de83fa910cf12cf15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2146018fa0d9020b06aea52c4bd07388a7d9b83327b17515b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7776d0b626a2c14ca4a959ad981652533f7d23220efc9335;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30e2150373373cecde0cdf59527fd731c13b8e098348d4d9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18e0b39f38750bbbefe358d9d5b63e039eb0ca6f6f7bbbc3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc5d5c5ef0f2ed53ca208776b9448d89af51c5a407938933e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e502cfd0424cc28caf4767ffad7936c1b4e68edeb79f6222;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6808115125cbd3c16404ade882a6048ee3cf1a32ea20a2547;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb2ed3a21499a1c2afeafd70c88b536c56c79cd239c5bcce8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h722024f4da0b400dda156d963289cffa2535b90bb7b47fbe4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb081e5efa9def2e70898b3cf50a53630f0f438a63368a4d3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c269a038adeded6d8728e7a2eaf75a4aba552085fb9dfd91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68546d3e01de7ca18265121d15622466217f2fce7f19b7444;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0f55b6bec2205e7c59884104241921efac2e4025e3f12391;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3c8445036d732e4100e389eaad03d5abcd479c94e0060601;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eaa71ee631a7bd9ceb92dcdc9b34e22295733d001000875d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf92f663338c0fabefd01db63029475fb3fda41a6786f185f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5d02e644cc8a02b9054c1c4e089f53a846161ac244ed9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h318a08433c11bb3044cec8db51f0a47dc90d7544cc8136261;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbfae75fd7a258aa1933863fc0a547de4b6e725604231eef1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h768429067b63a3a3de394dcf80c9e3108c40a8ddbea82cd18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h996683d3604f644f08d87cff78a49fdaad357d68ade672520;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha103da13121b7ca5ba41f6b1abff77d03544cb4ddea1c7ce1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1e8d0f164878f927146d50dcf19da9e3fe7e9f9c27e77dde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5af2d2ee057e4c139d2be4f6be2769cb51aaee4fccd7770a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h497d024622a55a4f1c59d0d60dbf1ee893c09381766778514;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a6f789995abe0418920b35c1582e0a51d2b701402b66cf19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0174fbbc6e8080992fe460eb90c1cb2ed4b82d86e549aed1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cfee44cccc4c4402a98a3415019cbdb570f8a9099d468233;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd281adb1d663fc8190227f7fa73774bfbe99e2152ae6c684;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cf7a7b4fddd5db7138a10908652e59f4ba8e8b77c89d31b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a4753e472cb69dd11eb9b1305c3acfabacb293e18336cc8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf59711064785493a9584f184de9a86974e8a06ae7bc10cecb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96f3d24037688fb86c8022b264f88c3ab4292e7c19357bc80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h733d3323b349d22ea20981aa02defa54b393af8f848965656;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9ffdda951fc30e34b50710d540520c54e69d7ff7657aaf4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73b9132136c92501e2cae0c06e73815314b4719e625f783e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a1208a45e6e7223aac0bf7065d24e4cd20ac3114c1650295;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he829920c34088d0caa31dea7f46a42ea4503087cae00fce97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2266e3b009baf1f1da5af5a37c6a102482dc73a907ee8cc3;
        #1
        $finish();
    end
endmodule
