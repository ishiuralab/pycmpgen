module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    compressor2_1_32_32 compressor2_1_32_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
        src16 <= 32'h0;
        src17 <= 32'h0;
        src18 <= 32'h0;
        src19 <= 32'h0;
        src20 <= 32'h0;
        src21 <= 32'h0;
        src22 <= 32'h0;
        src23 <= 32'h0;
        src24 <= 32'h0;
        src25 <= 32'h0;
        src26 <= 32'h0;
        src27 <= 32'h0;
        src28 <= 32'h0;
        src29 <= 32'h0;
        src30 <= 32'h0;
        src31 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_32_32(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    input [31:0]src16,
    input [31:0]src17,
    input [31:0]src18,
    input [31:0]src19,
    input [31:0]src20,
    input [31:0]src21,
    input [31:0]src22,
    input [31:0]src23,
    input [31:0]src24,
    input [31:0]src25,
    input [31:0]src26,
    input [31:0]src27,
    input [31:0]src28,
    input [31:0]src29,
    input [31:0]src30,
    input [31:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [0:0] comp_out33;
    wire [0:0] comp_out34;
    wire [0:0] comp_out35;
    wire [1:0] comp_out36;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36)
    );
    rowadder2_1_37 rowadder2_1inst(
        .src0({comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out36[1], 1'h0, 1'h0, 1'h0, comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst0({dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [0:0] dst33,
      output wire [0:0] dst34,
      output wire [0:0] dst35,
      output wire [1:0] dst36);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [31:0] stage0_16;
   wire [31:0] stage0_17;
   wire [31:0] stage0_18;
   wire [31:0] stage0_19;
   wire [31:0] stage0_20;
   wire [31:0] stage0_21;
   wire [31:0] stage0_22;
   wire [31:0] stage0_23;
   wire [31:0] stage0_24;
   wire [31:0] stage0_25;
   wire [31:0] stage0_26;
   wire [31:0] stage0_27;
   wire [31:0] stage0_28;
   wire [31:0] stage0_29;
   wire [31:0] stage0_30;
   wire [31:0] stage0_31;
   wire [10:0] stage1_0;
   wire [14:0] stage1_1;
   wire [11:0] stage1_2;
   wire [12:0] stage1_3;
   wire [18:0] stage1_4;
   wire [11:0] stage1_5;
   wire [12:0] stage1_6;
   wire [20:0] stage1_7;
   wire [11:0] stage1_8;
   wire [17:0] stage1_9;
   wire [11:0] stage1_10;
   wire [15:0] stage1_11;
   wire [12:0] stage1_12;
   wire [14:0] stage1_13;
   wire [12:0] stage1_14;
   wire [17:0] stage1_15;
   wire [12:0] stage1_16;
   wire [18:0] stage1_17;
   wire [16:0] stage1_18;
   wire [11:0] stage1_19;
   wire [12:0] stage1_20;
   wire [14:0] stage1_21;
   wire [11:0] stage1_22;
   wire [13:0] stage1_23;
   wire [22:0] stage1_24;
   wire [14:0] stage1_25;
   wire [11:0] stage1_26;
   wire [15:0] stage1_27;
   wire [16:0] stage1_28;
   wire [13:0] stage1_29;
   wire [22:0] stage1_30;
   wire [9:0] stage1_31;
   wire [7:0] stage1_32;
   wire [4:0] stage1_33;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [3:0] stage2_2;
   wire [4:0] stage2_3;
   wire [10:0] stage2_4;
   wire [5:0] stage2_5;
   wire [3:0] stage2_6;
   wire [5:0] stage2_7;
   wire [7:0] stage2_8;
   wire [12:0] stage2_9;
   wire [3:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [9:0] stage2_14;
   wire [5:0] stage2_15;
   wire [7:0] stage2_16;
   wire [5:0] stage2_17;
   wire [5:0] stage2_18;
   wire [10:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [5:0] stage2_22;
   wire [3:0] stage2_23;
   wire [8:0] stage2_24;
   wire [7:0] stage2_25;
   wire [5:0] stage2_26;
   wire [8:0] stage2_27;
   wire [7:0] stage2_28;
   wire [5:0] stage2_29;
   wire [5:0] stage2_30;
   wire [6:0] stage2_31;
   wire [6:0] stage2_32;
   wire [2:0] stage2_33;
   wire [1:0] stage2_34;
   wire [0:0] stage2_35;
   wire [1:0] stage3_0;
   wire [0:0] stage3_1;
   wire [1:0] stage3_2;
   wire [3:0] stage3_3;
   wire [6:0] stage3_4;
   wire [1:0] stage3_5;
   wire [5:0] stage3_6;
   wire [0:0] stage3_7;
   wire [6:0] stage3_8;
   wire [4:0] stage3_9;
   wire [2:0] stage3_10;
   wire [1:0] stage3_11;
   wire [6:0] stage3_12;
   wire [5:0] stage3_13;
   wire [1:0] stage3_14;
   wire [5:0] stage3_15;
   wire [2:0] stage3_16;
   wire [5:0] stage3_17;
   wire [1:0] stage3_18;
   wire [2:0] stage3_19;
   wire [5:0] stage3_20;
   wire [3:0] stage3_21;
   wire [2:0] stage3_22;
   wire [3:0] stage3_23;
   wire [5:0] stage3_24;
   wire [2:0] stage3_25;
   wire [1:0] stage3_26;
   wire [4:0] stage3_27;
   wire [5:0] stage3_28;
   wire [6:0] stage3_29;
   wire [0:0] stage3_30;
   wire [1:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [2:0] stage3_34;
   wire [0:0] stage3_35;
   wire [0:0] stage3_36;
   wire [1:0] stage4_0;
   wire [0:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [0:0] stage4_35;
   wire [1:0] stage4_36;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;

   gpc1406_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[4]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[5]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[6]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9]},
      {stage1_5[0],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc615_5 gpc7 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[7],stage1_3[7],stage1_2[7]}
   );
   gpc615_5 gpc8 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage0_3[11]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[2],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[3],stage1_4[9],stage1_3[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[4],stage1_4[10],stage1_3[10]}
   );
   gpc615_5 gpc11 (
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[5],stage1_4[11],stage1_3[11]}
   );
   gpc615_5 gpc12 (
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage0_4[15]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[5],stage1_5[6],stage1_4[12],stage1_3[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[4],stage1_6[6],stage1_5[7],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[5],stage1_6[7],stage1_5[8],stage1_4[14]}
   );
   gpc606_5 gpc15 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[2],stage1_7[6],stage1_6[8],stage1_5[9]}
   );
   gpc135_4 gpc16 (
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16]},
      {stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage0_8[0]},
      {stage1_9[1],stage1_8[3],stage1_7[7],stage1_6[9]}
   );
   gpc135_4 gpc17 (
      {stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21]},
      {stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage0_8[1]},
      {stage1_9[2],stage1_8[4],stage1_7[8],stage1_6[10]}
   );
   gpc135_4 gpc18 (
      {stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage0_8[2]},
      {stage1_9[3],stage1_8[5],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc19 (
      {stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30], stage0_6[31]},
      {stage0_7[15]},
      {stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8]},
      {stage1_10[0],stage1_9[4],stage1_8[6],stage1_7[10],stage1_6[12]}
   );
   gpc1343_5 gpc20 (
      {stage0_7[16], stage0_7[17], stage0_7[18]},
      {stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[7],stage1_7[11]}
   );
   gpc615_5 gpc21 (
      {stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage0_8[13]},
      {stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[8],stage1_7[12]}
   );
   gpc606_5 gpc22 (
      {stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[0],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[9]}
   );
   gpc606_5 gpc23 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[1],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[10]}
   );
   gpc606_5 gpc24 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[2],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[11]}
   );
   gpc606_5 gpc25 (
      {stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[3],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc606_5 gpc26 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[4],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc606_5 gpc27 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[5],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc606_5 gpc28 (
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[6],stage1_11[8],stage1_10[9]}
   );
   gpc606_5 gpc29 (
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[7],stage1_11[9],stage1_10[10]}
   );
   gpc615_5 gpc30 (
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[5],stage1_12[8],stage1_11[10]}
   );
   gpc615_5 gpc31 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[6],stage1_12[9],stage1_11[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[2],stage1_14[4],stage1_13[7],stage1_12[10]}
   );
   gpc606_5 gpc33 (
      {stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[3],stage1_14[5],stage1_13[8],stage1_12[11]}
   );
   gpc606_5 gpc34 (
      {stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[4],stage1_14[6],stage1_13[9],stage1_12[12]}
   );
   gpc606_5 gpc35 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[5],stage1_14[7],stage1_13[10]}
   );
   gpc606_5 gpc36 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[6],stage1_14[8],stage1_13[11]}
   );
   gpc606_5 gpc37 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[5],stage1_15[7],stage1_14[9],stage1_13[12]}
   );
   gpc615_5 gpc38 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22]},
      {stage0_15[18]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[6],stage1_15[8],stage1_14[10]}
   );
   gpc615_5 gpc39 (
      {stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage0_15[19]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[7],stage1_15[9],stage1_14[11]}
   );
   gpc615_5 gpc40 (
      {stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31], 1'b0},
      {stage0_15[20]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[5],stage1_16[8],stage1_15[10],stage1_14[12]}
   );
   gpc615_5 gpc41 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[6],stage1_16[9],stage1_15[11]}
   );
   gpc606_5 gpc42 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[1],stage1_18[4],stage1_17[7],stage1_16[10]}
   );
   gpc606_5 gpc43 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[2],stage1_18[5],stage1_17[8],stage1_16[11]}
   );
   gpc615_5 gpc44 (
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10]},
      {stage0_18[12]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[2],stage1_19[3],stage1_18[6],stage1_17[9]}
   );
   gpc615_5 gpc45 (
      {stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_18[13]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[3],stage1_19[4],stage1_18[7],stage1_17[10]}
   );
   gpc615_5 gpc46 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage0_18[14]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[4],stage1_19[5],stage1_18[8],stage1_17[11]}
   );
   gpc615_5 gpc47 (
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25]},
      {stage0_18[15]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[5],stage1_19[6],stage1_18[9],stage1_17[12]}
   );
   gpc606_5 gpc48 (
      {stage0_18[16], stage0_18[17], stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[4],stage1_20[6],stage1_19[7],stage1_18[10]}
   );
   gpc615_5 gpc49 (
      {stage0_18[22], stage0_18[23], stage0_18[24], stage0_18[25], stage0_18[26]},
      {stage0_19[24]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[5],stage1_20[7],stage1_19[8],stage1_18[11]}
   );
   gpc615_5 gpc50 (
      {stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[6],stage1_20[8],stage1_19[9]}
   );
   gpc615_5 gpc51 (
      {stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage0_21[6]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[1],stage1_22[3],stage1_21[7],stage1_20[9]}
   );
   gpc615_5 gpc52 (
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22]},
      {stage0_21[7]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[2],stage1_22[4],stage1_21[8],stage1_20[10]}
   );
   gpc615_5 gpc53 (
      {stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_21[8]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[3],stage1_22[5],stage1_21[9],stage1_20[11]}
   );
   gpc615_5 gpc54 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], 1'b0},
      {stage0_21[9]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[4],stage1_22[6],stage1_21[10],stage1_20[12]}
   );
   gpc606_5 gpc55 (
      {stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[4],stage1_23[5],stage1_22[7],stage1_21[11]}
   );
   gpc606_5 gpc56 (
      {stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[5],stage1_23[6],stage1_22[8],stage1_21[12]}
   );
   gpc615_5 gpc57 (
      {stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_22[24]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[6],stage1_23[7],stage1_22[9],stage1_21[13]}
   );
   gpc615_5 gpc58 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage0_22[25]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[7],stage1_23[8],stage1_22[10],stage1_21[14]}
   );
   gpc606_5 gpc59 (
      {stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[4],stage1_24[8],stage1_23[9],stage1_22[11]}
   );
   gpc615_5 gpc60 (
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28]},
      {stage0_24[6]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[5],stage1_24[9],stage1_23[10]}
   );
   gpc615_5 gpc61 (
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_25[6]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[6],stage1_24[10]}
   );
   gpc615_5 gpc62 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16]},
      {stage0_25[7]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[7],stage1_24[11]}
   );
   gpc615_5 gpc63 (
      {stage0_24[17], stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21]},
      {stage0_25[8]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[8],stage1_24[12]}
   );
   gpc606_5 gpc64 (
      {stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13], stage0_25[14]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[3],stage1_27[4],stage1_26[5],stage1_25[9]}
   );
   gpc615_5 gpc65 (
      {stage0_25[15], stage0_25[16], stage0_25[17], stage0_25[18], stage0_25[19]},
      {stage0_26[18]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[4],stage1_27[5],stage1_26[6],stage1_25[10]}
   );
   gpc615_5 gpc66 (
      {stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23], stage0_25[24]},
      {stage0_26[19]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[5],stage1_27[6],stage1_26[7],stage1_25[11]}
   );
   gpc615_5 gpc67 (
      {stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_26[20]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[6],stage1_27[7],stage1_26[8],stage1_25[12]}
   );
   gpc615_5 gpc68 (
      {stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24], stage0_26[25]},
      {stage0_27[24]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[4],stage1_28[7],stage1_27[8],stage1_26[9]}
   );
   gpc615_5 gpc69 (
      {stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29], stage0_26[30]},
      {stage0_27[25]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[5],stage1_28[8],stage1_27[9],stage1_26[10]}
   );
   gpc615_5 gpc70 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16]},
      {stage0_29[0]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[0],stage1_30[2],stage1_29[6],stage1_28[9]}
   );
   gpc615_5 gpc71 (
      {stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage0_29[1]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[1],stage1_30[3],stage1_29[7],stage1_28[10]}
   );
   gpc615_5 gpc72 (
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26]},
      {stage0_29[2]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[2],stage1_30[4],stage1_29[8],stage1_28[11]}
   );
   gpc606_5 gpc73 (
      {stage0_29[3], stage0_29[4], stage0_29[5], stage0_29[6], stage0_29[7], stage0_29[8]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[3],stage1_30[5],stage1_29[9]}
   );
   gpc606_5 gpc74 (
      {stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13], stage0_29[14]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[4],stage1_30[6],stage1_29[10]}
   );
   gpc606_5 gpc75 (
      {stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19], stage0_29[20]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[5],stage1_30[7],stage1_29[11]}
   );
   gpc606_5 gpc76 (
      {stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[6],stage1_30[8],stage1_29[12]}
   );
   gpc615_5 gpc77 (
      {stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_30[18]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[7],stage1_31[7],stage1_30[9],stage1_29[13]}
   );
   gpc1_1 gpc78 (
      {stage0_0[27]},
      {stage1_0[6]}
   );
   gpc1_1 gpc79 (
      {stage0_0[28]},
      {stage1_0[7]}
   );
   gpc1_1 gpc80 (
      {stage0_0[29]},
      {stage1_0[8]}
   );
   gpc1_1 gpc81 (
      {stage0_0[30]},
      {stage1_0[9]}
   );
   gpc1_1 gpc82 (
      {stage0_0[31]},
      {stage1_0[10]}
   );
   gpc1_1 gpc83 (
      {stage0_1[24]},
      {stage1_1[7]}
   );
   gpc1_1 gpc84 (
      {stage0_1[25]},
      {stage1_1[8]}
   );
   gpc1_1 gpc85 (
      {stage0_1[26]},
      {stage1_1[9]}
   );
   gpc1_1 gpc86 (
      {stage0_1[27]},
      {stage1_1[10]}
   );
   gpc1_1 gpc87 (
      {stage0_1[28]},
      {stage1_1[11]}
   );
   gpc1_1 gpc88 (
      {stage0_1[29]},
      {stage1_1[12]}
   );
   gpc1_1 gpc89 (
      {stage0_1[30]},
      {stage1_1[13]}
   );
   gpc1_1 gpc90 (
      {stage0_1[31]},
      {stage1_1[14]}
   );
   gpc1_1 gpc91 (
      {stage0_2[29]},
      {stage1_2[9]}
   );
   gpc1_1 gpc92 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc93 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc94 (
      {stage0_4[28]},
      {stage1_4[15]}
   );
   gpc1_1 gpc95 (
      {stage0_4[29]},
      {stage1_4[16]}
   );
   gpc1_1 gpc96 (
      {stage0_4[30]},
      {stage1_4[17]}
   );
   gpc1_1 gpc97 (
      {stage0_4[31]},
      {stage1_4[18]}
   );
   gpc1_1 gpc98 (
      {stage0_5[30]},
      {stage1_5[10]}
   );
   gpc1_1 gpc99 (
      {stage0_5[31]},
      {stage1_5[11]}
   );
   gpc1_1 gpc100 (
      {stage0_7[24]},
      {stage1_7[13]}
   );
   gpc1_1 gpc101 (
      {stage0_7[25]},
      {stage1_7[14]}
   );
   gpc1_1 gpc102 (
      {stage0_7[26]},
      {stage1_7[15]}
   );
   gpc1_1 gpc103 (
      {stage0_7[27]},
      {stage1_7[16]}
   );
   gpc1_1 gpc104 (
      {stage0_7[28]},
      {stage1_7[17]}
   );
   gpc1_1 gpc105 (
      {stage0_7[29]},
      {stage1_7[18]}
   );
   gpc1_1 gpc106 (
      {stage0_7[30]},
      {stage1_7[19]}
   );
   gpc1_1 gpc107 (
      {stage0_7[31]},
      {stage1_7[20]}
   );
   gpc1_1 gpc108 (
      {stage0_9[27]},
      {stage1_9[13]}
   );
   gpc1_1 gpc109 (
      {stage0_9[28]},
      {stage1_9[14]}
   );
   gpc1_1 gpc110 (
      {stage0_9[29]},
      {stage1_9[15]}
   );
   gpc1_1 gpc111 (
      {stage0_9[30]},
      {stage1_9[16]}
   );
   gpc1_1 gpc112 (
      {stage0_9[31]},
      {stage1_9[17]}
   );
   gpc1_1 gpc113 (
      {stage0_10[31]},
      {stage1_10[11]}
   );
   gpc1_1 gpc114 (
      {stage0_11[28]},
      {stage1_11[12]}
   );
   gpc1_1 gpc115 (
      {stage0_11[29]},
      {stage1_11[13]}
   );
   gpc1_1 gpc116 (
      {stage0_11[30]},
      {stage1_11[14]}
   );
   gpc1_1 gpc117 (
      {stage0_11[31]},
      {stage1_11[15]}
   );
   gpc1_1 gpc118 (
      {stage0_13[30]},
      {stage1_13[13]}
   );
   gpc1_1 gpc119 (
      {stage0_13[31]},
      {stage1_13[14]}
   );
   gpc1_1 gpc120 (
      {stage0_15[26]},
      {stage1_15[12]}
   );
   gpc1_1 gpc121 (
      {stage0_15[27]},
      {stage1_15[13]}
   );
   gpc1_1 gpc122 (
      {stage0_15[28]},
      {stage1_15[14]}
   );
   gpc1_1 gpc123 (
      {stage0_15[29]},
      {stage1_15[15]}
   );
   gpc1_1 gpc124 (
      {stage0_15[30]},
      {stage1_15[16]}
   );
   gpc1_1 gpc125 (
      {stage0_15[31]},
      {stage1_15[17]}
   );
   gpc1_1 gpc126 (
      {stage0_16[31]},
      {stage1_16[12]}
   );
   gpc1_1 gpc127 (
      {stage0_17[26]},
      {stage1_17[13]}
   );
   gpc1_1 gpc128 (
      {stage0_17[27]},
      {stage1_17[14]}
   );
   gpc1_1 gpc129 (
      {stage0_17[28]},
      {stage1_17[15]}
   );
   gpc1_1 gpc130 (
      {stage0_17[29]},
      {stage1_17[16]}
   );
   gpc1_1 gpc131 (
      {stage0_17[30]},
      {stage1_17[17]}
   );
   gpc1_1 gpc132 (
      {stage0_17[31]},
      {stage1_17[18]}
   );
   gpc1_1 gpc133 (
      {stage0_18[27]},
      {stage1_18[12]}
   );
   gpc1_1 gpc134 (
      {stage0_18[28]},
      {stage1_18[13]}
   );
   gpc1_1 gpc135 (
      {stage0_18[29]},
      {stage1_18[14]}
   );
   gpc1_1 gpc136 (
      {stage0_18[30]},
      {stage1_18[15]}
   );
   gpc1_1 gpc137 (
      {stage0_18[31]},
      {stage1_18[16]}
   );
   gpc1_1 gpc138 (
      {stage0_19[30]},
      {stage1_19[10]}
   );
   gpc1_1 gpc139 (
      {stage0_19[31]},
      {stage1_19[11]}
   );
   gpc1_1 gpc140 (
      {stage0_23[29]},
      {stage1_23[11]}
   );
   gpc1_1 gpc141 (
      {stage0_23[30]},
      {stage1_23[12]}
   );
   gpc1_1 gpc142 (
      {stage0_23[31]},
      {stage1_23[13]}
   );
   gpc1_1 gpc143 (
      {stage0_24[22]},
      {stage1_24[13]}
   );
   gpc1_1 gpc144 (
      {stage0_24[23]},
      {stage1_24[14]}
   );
   gpc1_1 gpc145 (
      {stage0_24[24]},
      {stage1_24[15]}
   );
   gpc1_1 gpc146 (
      {stage0_24[25]},
      {stage1_24[16]}
   );
   gpc1_1 gpc147 (
      {stage0_24[26]},
      {stage1_24[17]}
   );
   gpc1_1 gpc148 (
      {stage0_24[27]},
      {stage1_24[18]}
   );
   gpc1_1 gpc149 (
      {stage0_24[28]},
      {stage1_24[19]}
   );
   gpc1_1 gpc150 (
      {stage0_24[29]},
      {stage1_24[20]}
   );
   gpc1_1 gpc151 (
      {stage0_24[30]},
      {stage1_24[21]}
   );
   gpc1_1 gpc152 (
      {stage0_24[31]},
      {stage1_24[22]}
   );
   gpc1_1 gpc153 (
      {stage0_25[30]},
      {stage1_25[13]}
   );
   gpc1_1 gpc154 (
      {stage0_25[31]},
      {stage1_25[14]}
   );
   gpc1_1 gpc155 (
      {stage0_26[31]},
      {stage1_26[11]}
   );
   gpc1_1 gpc156 (
      {stage0_27[26]},
      {stage1_27[10]}
   );
   gpc1_1 gpc157 (
      {stage0_27[27]},
      {stage1_27[11]}
   );
   gpc1_1 gpc158 (
      {stage0_27[28]},
      {stage1_27[12]}
   );
   gpc1_1 gpc159 (
      {stage0_27[29]},
      {stage1_27[13]}
   );
   gpc1_1 gpc160 (
      {stage0_27[30]},
      {stage1_27[14]}
   );
   gpc1_1 gpc161 (
      {stage0_27[31]},
      {stage1_27[15]}
   );
   gpc1_1 gpc162 (
      {stage0_28[27]},
      {stage1_28[12]}
   );
   gpc1_1 gpc163 (
      {stage0_28[28]},
      {stage1_28[13]}
   );
   gpc1_1 gpc164 (
      {stage0_28[29]},
      {stage1_28[14]}
   );
   gpc1_1 gpc165 (
      {stage0_28[30]},
      {stage1_28[15]}
   );
   gpc1_1 gpc166 (
      {stage0_28[31]},
      {stage1_28[16]}
   );
   gpc1_1 gpc167 (
      {stage0_30[19]},
      {stage1_30[10]}
   );
   gpc1_1 gpc168 (
      {stage0_30[20]},
      {stage1_30[11]}
   );
   gpc1_1 gpc169 (
      {stage0_30[21]},
      {stage1_30[12]}
   );
   gpc1_1 gpc170 (
      {stage0_30[22]},
      {stage1_30[13]}
   );
   gpc1_1 gpc171 (
      {stage0_30[23]},
      {stage1_30[14]}
   );
   gpc1_1 gpc172 (
      {stage0_30[24]},
      {stage1_30[15]}
   );
   gpc1_1 gpc173 (
      {stage0_30[25]},
      {stage1_30[16]}
   );
   gpc1_1 gpc174 (
      {stage0_30[26]},
      {stage1_30[17]}
   );
   gpc1_1 gpc175 (
      {stage0_30[27]},
      {stage1_30[18]}
   );
   gpc1_1 gpc176 (
      {stage0_30[28]},
      {stage1_30[19]}
   );
   gpc1_1 gpc177 (
      {stage0_30[29]},
      {stage1_30[20]}
   );
   gpc1_1 gpc178 (
      {stage0_30[30]},
      {stage1_30[21]}
   );
   gpc1_1 gpc179 (
      {stage0_30[31]},
      {stage1_30[22]}
   );
   gpc1_1 gpc180 (
      {stage0_31[30]},
      {stage1_31[8]}
   );
   gpc1_1 gpc181 (
      {stage0_31[31]},
      {stage1_31[9]}
   );
   gpc606_5 gpc182 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc183 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], 1'b0},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc184 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc185 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1163_5 gpc186 (
      {stage1_4[0], stage1_4[1], stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc187 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc188 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc189 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[3],stage2_7[3],stage2_6[3],stage2_5[5]}
   );
   gpc7_3 gpc190 (
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[4],stage2_7[4]}
   );
   gpc7_3 gpc191 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20]},
      {stage2_9[2],stage2_8[5],stage2_7[5]}
   );
   gpc606_5 gpc192 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[3],stage2_8[6]}
   );
   gpc606_5 gpc193 (
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[4],stage2_8[7]}
   );
   gpc606_5 gpc194 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[2],stage2_9[5]}
   );
   gpc606_5 gpc195 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[3],stage2_9[6]}
   );
   gpc615_5 gpc196 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], 1'b0},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[4]}
   );
   gpc2135_5 gpc197 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage1_14[0]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc198 (
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc199 (
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[5]}
   );
   gpc615_5 gpc200 (
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[3],stage2_15[4]}
   );
   gpc615_5 gpc201 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[4],stage2_15[5]}
   );
   gpc615_5 gpc202 (
      {stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[12]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[3],stage2_16[5]}
   );
   gpc615_5 gpc203 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage1_17[13]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[3],stage2_18[3],stage2_17[4],stage2_16[6]}
   );
   gpc615_5 gpc204 (
      {stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_18[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[4],stage2_18[4],stage2_17[5]}
   );
   gpc615_5 gpc205 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], 1'b0},
      {stage1_19[6]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[5],stage2_18[5]}
   );
   gpc606_5 gpc206 (
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[2]}
   );
   gpc2135_5 gpc207 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4]},
      {stage1_23[6], stage1_23[7], stage1_23[8]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1]},
      {stage2_26[0],stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2]}
   );
   gpc615_5 gpc208 (
      {stage1_22[5], stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9]},
      {stage1_23[9]},
      {stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage2_26[1],stage2_25[2],stage2_24[2],stage2_23[2],stage2_22[3]}
   );
   gpc615_5 gpc209 (
      {stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13], 1'b0},
      {stage1_24[7]},
      {stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[3],stage2_23[3]}
   );
   gpc606_5 gpc210 (
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[4]}
   );
   gpc606_5 gpc211 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[5]}
   );
   gpc606_5 gpc212 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[3],stage2_26[5],stage2_25[6]}
   );
   gpc606_5 gpc213 (
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[1],stage2_28[3],stage2_27[4]}
   );
   gpc606_5 gpc214 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[1],stage2_29[2],stage2_28[4]}
   );
   gpc615_5 gpc215 (
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10]},
      {stage1_29[6]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[2],stage2_30[2],stage2_29[3],stage2_28[5]}
   );
   gpc615_5 gpc216 (
      {stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15]},
      {stage1_29[7]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[3],stage2_30[3],stage2_29[4],stage2_28[6]}
   );
   gpc606_5 gpc217 (
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[3],stage2_31[4],stage2_30[4],stage2_29[5]}
   );
   gpc606_5 gpc218 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], 1'b0},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[4],stage2_31[5],stage2_30[5]}
   );
   gpc615_5 gpc219 (
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], 1'b0},
      {stage1_32[6]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], 1'b0},
      {stage2_35[0],stage2_34[1],stage2_33[2],stage2_32[5],stage2_31[6]}
   );
   gpc1_1 gpc220 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc221 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc222 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc223 (
      {stage1_3[12]},
      {stage2_3[4]}
   );
   gpc1_1 gpc224 (
      {stage1_4[15]},
      {stage2_4[7]}
   );
   gpc1_1 gpc225 (
      {stage1_4[16]},
      {stage2_4[8]}
   );
   gpc1_1 gpc226 (
      {stage1_4[17]},
      {stage2_4[9]}
   );
   gpc1_1 gpc227 (
      {stage1_4[18]},
      {stage2_4[10]}
   );
   gpc1_1 gpc228 (
      {stage1_9[12]},
      {stage2_9[7]}
   );
   gpc1_1 gpc229 (
      {stage1_9[13]},
      {stage2_9[8]}
   );
   gpc1_1 gpc230 (
      {stage1_9[14]},
      {stage2_9[9]}
   );
   gpc1_1 gpc231 (
      {stage1_9[15]},
      {stage2_9[10]}
   );
   gpc1_1 gpc232 (
      {stage1_9[16]},
      {stage2_9[11]}
   );
   gpc1_1 gpc233 (
      {stage1_9[17]},
      {stage2_9[12]}
   );
   gpc1_1 gpc234 (
      {stage1_12[12]},
      {stage2_12[7]}
   );
   gpc1_1 gpc235 (
      {stage1_14[7]},
      {stage2_14[4]}
   );
   gpc1_1 gpc236 (
      {stage1_14[8]},
      {stage2_14[5]}
   );
   gpc1_1 gpc237 (
      {stage1_14[9]},
      {stage2_14[6]}
   );
   gpc1_1 gpc238 (
      {stage1_14[10]},
      {stage2_14[7]}
   );
   gpc1_1 gpc239 (
      {stage1_14[11]},
      {stage2_14[8]}
   );
   gpc1_1 gpc240 (
      {stage1_14[12]},
      {stage2_14[9]}
   );
   gpc1_1 gpc241 (
      {stage1_16[12]},
      {stage2_16[7]}
   );
   gpc1_1 gpc242 (
      {stage1_19[7]},
      {stage2_19[6]}
   );
   gpc1_1 gpc243 (
      {stage1_19[8]},
      {stage2_19[7]}
   );
   gpc1_1 gpc244 (
      {stage1_19[9]},
      {stage2_19[8]}
   );
   gpc1_1 gpc245 (
      {stage1_19[10]},
      {stage2_19[9]}
   );
   gpc1_1 gpc246 (
      {stage1_19[11]},
      {stage2_19[10]}
   );
   gpc1_1 gpc247 (
      {stage1_20[6]},
      {stage2_20[4]}
   );
   gpc1_1 gpc248 (
      {stage1_20[7]},
      {stage2_20[5]}
   );
   gpc1_1 gpc249 (
      {stage1_20[8]},
      {stage2_20[6]}
   );
   gpc1_1 gpc250 (
      {stage1_20[9]},
      {stage2_20[7]}
   );
   gpc1_1 gpc251 (
      {stage1_20[10]},
      {stage2_20[8]}
   );
   gpc1_1 gpc252 (
      {stage1_20[11]},
      {stage2_20[9]}
   );
   gpc1_1 gpc253 (
      {stage1_20[12]},
      {stage2_20[10]}
   );
   gpc1_1 gpc254 (
      {stage1_21[6]},
      {stage2_21[3]}
   );
   gpc1_1 gpc255 (
      {stage1_21[7]},
      {stage2_21[4]}
   );
   gpc1_1 gpc256 (
      {stage1_21[8]},
      {stage2_21[5]}
   );
   gpc1_1 gpc257 (
      {stage1_21[9]},
      {stage2_21[6]}
   );
   gpc1_1 gpc258 (
      {stage1_21[10]},
      {stage2_21[7]}
   );
   gpc1_1 gpc259 (
      {stage1_21[11]},
      {stage2_21[8]}
   );
   gpc1_1 gpc260 (
      {stage1_21[12]},
      {stage2_21[9]}
   );
   gpc1_1 gpc261 (
      {stage1_21[13]},
      {stage2_21[10]}
   );
   gpc1_1 gpc262 (
      {stage1_21[14]},
      {stage2_21[11]}
   );
   gpc1_1 gpc263 (
      {stage1_22[10]},
      {stage2_22[4]}
   );
   gpc1_1 gpc264 (
      {stage1_22[11]},
      {stage2_22[5]}
   );
   gpc1_1 gpc265 (
      {stage1_24[20]},
      {stage2_24[6]}
   );
   gpc1_1 gpc266 (
      {stage1_24[21]},
      {stage2_24[7]}
   );
   gpc1_1 gpc267 (
      {stage1_24[22]},
      {stage2_24[8]}
   );
   gpc1_1 gpc268 (
      {stage1_25[14]},
      {stage2_25[7]}
   );
   gpc1_1 gpc269 (
      {stage1_27[12]},
      {stage2_27[5]}
   );
   gpc1_1 gpc270 (
      {stage1_27[13]},
      {stage2_27[6]}
   );
   gpc1_1 gpc271 (
      {stage1_27[14]},
      {stage2_27[7]}
   );
   gpc1_1 gpc272 (
      {stage1_27[15]},
      {stage2_27[8]}
   );
   gpc1_1 gpc273 (
      {stage1_28[16]},
      {stage2_28[7]}
   );
   gpc1_1 gpc274 (
      {stage1_32[7]},
      {stage2_32[6]}
   );
   gpc207_4 gpc275 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc276 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], 1'b0},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc277 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc23_3 gpc278 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[1],stage3_8[1]}
   );
   gpc2135_5 gpc279 (
      {stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[2]}
   );
   gpc1415_5 gpc280 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage2_10[3]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[2]},
      {stage3_13[1],stage3_12[1],stage3_11[1],stage3_10[2],stage3_9[3]}
   );
   gpc1163_5 gpc281 (
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_15[0]},
      {stage2_16[0]},
      {stage3_17[0],stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2]}
   );
   gpc615_5 gpc282 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], 1'b0},
      {stage2_15[1]},
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage3_18[0],stage3_17[1],stage3_16[1],stage3_15[1],stage3_14[1]}
   );
   gpc1163_5 gpc283 (
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage2_19[0]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[1],stage3_17[2]}
   );
   gpc615_5 gpc284 (
      {stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[1]}
   );
   gpc615_5 gpc285 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10]},
      {stage2_20[2]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[1],stage3_21[2],stage3_20[2],stage3_19[2]}
   );
   gpc606_5 gpc286 (
      {stage2_20[3], stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[2],stage3_21[3],stage3_20[3]}
   );
   gpc615_5 gpc287 (
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], 1'b0},
      {stage2_24[0]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1],stage3_23[3]}
   );
   gpc615_5 gpc288 (
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage2_25[6]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[2]}
   );
   gpc7_3 gpc289 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage3_29[0],stage3_28[1],stage3_27[2]}
   );
   gpc615_5 gpc290 (
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4]},
      {stage2_29[0]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[0],stage3_29[1],stage3_28[2]}
   );
   gpc117_4 gpc291 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5], stage2_31[6]},
      {stage2_32[0]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[1]}
   );
   gpc2135_5 gpc292 (
      {stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage2_33[1], stage2_33[2], 1'b0},
      {stage2_34[0]},
      {stage2_35[0], 1'b0},
      {stage3_36[0],stage3_35[0],stage3_34[1],stage3_33[1],stage3_32[2]}
   );
   gpc1_1 gpc293 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc294 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc295 (
      {stage2_3[3]},
      {stage3_3[2]}
   );
   gpc1_1 gpc296 (
      {stage2_3[4]},
      {stage3_3[3]}
   );
   gpc1_1 gpc297 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc298 (
      {stage2_4[7]},
      {stage3_4[3]}
   );
   gpc1_1 gpc299 (
      {stage2_4[8]},
      {stage3_4[4]}
   );
   gpc1_1 gpc300 (
      {stage2_4[9]},
      {stage3_4[5]}
   );
   gpc1_1 gpc301 (
      {stage2_4[10]},
      {stage3_4[6]}
   );
   gpc1_1 gpc302 (
      {stage2_6[0]},
      {stage3_6[2]}
   );
   gpc1_1 gpc303 (
      {stage2_6[1]},
      {stage3_6[3]}
   );
   gpc1_1 gpc304 (
      {stage2_6[2]},
      {stage3_6[4]}
   );
   gpc1_1 gpc305 (
      {stage2_6[3]},
      {stage3_6[5]}
   );
   gpc1_1 gpc306 (
      {stage2_8[3]},
      {stage3_8[2]}
   );
   gpc1_1 gpc307 (
      {stage2_8[4]},
      {stage3_8[3]}
   );
   gpc1_1 gpc308 (
      {stage2_8[5]},
      {stage3_8[4]}
   );
   gpc1_1 gpc309 (
      {stage2_8[6]},
      {stage3_8[5]}
   );
   gpc1_1 gpc310 (
      {stage2_8[7]},
      {stage3_8[6]}
   );
   gpc1_1 gpc311 (
      {stage2_9[12]},
      {stage3_9[4]}
   );
   gpc1_1 gpc312 (
      {stage2_12[3]},
      {stage3_12[2]}
   );
   gpc1_1 gpc313 (
      {stage2_12[4]},
      {stage3_12[3]}
   );
   gpc1_1 gpc314 (
      {stage2_12[5]},
      {stage3_12[4]}
   );
   gpc1_1 gpc315 (
      {stage2_12[6]},
      {stage3_12[5]}
   );
   gpc1_1 gpc316 (
      {stage2_12[7]},
      {stage3_12[6]}
   );
   gpc1_1 gpc317 (
      {stage2_13[3]},
      {stage3_13[3]}
   );
   gpc1_1 gpc318 (
      {stage2_13[4]},
      {stage3_13[4]}
   );
   gpc1_1 gpc319 (
      {stage2_13[5]},
      {stage3_13[5]}
   );
   gpc1_1 gpc320 (
      {stage2_15[2]},
      {stage3_15[2]}
   );
   gpc1_1 gpc321 (
      {stage2_15[3]},
      {stage3_15[3]}
   );
   gpc1_1 gpc322 (
      {stage2_15[4]},
      {stage3_15[4]}
   );
   gpc1_1 gpc323 (
      {stage2_15[5]},
      {stage3_15[5]}
   );
   gpc1_1 gpc324 (
      {stage2_16[7]},
      {stage3_16[2]}
   );
   gpc1_1 gpc325 (
      {stage2_17[3]},
      {stage3_17[3]}
   );
   gpc1_1 gpc326 (
      {stage2_17[4]},
      {stage3_17[4]}
   );
   gpc1_1 gpc327 (
      {stage2_17[5]},
      {stage3_17[5]}
   );
   gpc1_1 gpc328 (
      {stage2_20[9]},
      {stage3_20[4]}
   );
   gpc1_1 gpc329 (
      {stage2_20[10]},
      {stage3_20[5]}
   );
   gpc1_1 gpc330 (
      {stage2_24[6]},
      {stage3_24[3]}
   );
   gpc1_1 gpc331 (
      {stage2_24[7]},
      {stage3_24[4]}
   );
   gpc1_1 gpc332 (
      {stage2_24[8]},
      {stage3_24[5]}
   );
   gpc1_1 gpc333 (
      {stage2_25[7]},
      {stage3_25[2]}
   );
   gpc1_1 gpc334 (
      {stage2_27[7]},
      {stage3_27[3]}
   );
   gpc1_1 gpc335 (
      {stage2_27[8]},
      {stage3_27[4]}
   );
   gpc1_1 gpc336 (
      {stage2_28[5]},
      {stage3_28[3]}
   );
   gpc1_1 gpc337 (
      {stage2_28[6]},
      {stage3_28[4]}
   );
   gpc1_1 gpc338 (
      {stage2_28[7]},
      {stage3_28[5]}
   );
   gpc1_1 gpc339 (
      {stage2_29[1]},
      {stage3_29[2]}
   );
   gpc1_1 gpc340 (
      {stage2_29[2]},
      {stage3_29[3]}
   );
   gpc1_1 gpc341 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc342 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc343 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc344 (
      {stage2_32[6]},
      {stage3_32[3]}
   );
   gpc1_1 gpc345 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1163_5 gpc346 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc347 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1]}
   );
   gpc135_4 gpc348 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0], stage3_10[1], stage3_10[2]},
      {stage3_11[0]},
      {stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc207_4 gpc349 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc606_5 gpc350 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[1]}
   );
   gpc1163_5 gpc351 (
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[1]}
   );
   gpc1163_5 gpc352 (
      {stage3_19[1], stage3_19[2], 1'b0},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage3_21[0]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc1423_5 gpc353 (
      {stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[1], stage3_22[2]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3]},
      {stage3_24[0]},
      {stage4_25[0],stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1]}
   );
   gpc135_4 gpc354 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage4_27[0],stage4_26[0],stage4_25[1],stage4_24[1]}
   );
   gpc615_5 gpc355 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4]},
      {stage3_28[0]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc2116_5 gpc356 (
      {stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5], 1'b0},
      {stage3_29[6]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[1],stage4_28[1]}
   );
   gpc1325_5 gpc357 (
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], 1'b0},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[1]}
   );
   gpc1_1 gpc358 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc359 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc360 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc361 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc362 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc363 (
      {stage3_3[3]},
      {stage4_3[1]}
   );
   gpc1_1 gpc364 (
      {stage3_4[6]},
      {stage4_4[1]}
   );
   gpc1_1 gpc365 (
      {stage3_5[1]},
      {stage4_5[1]}
   );
   gpc1_1 gpc366 (
      {stage3_8[6]},
      {stage4_8[1]}
   );
   gpc1_1 gpc367 (
      {stage3_11[1]},
      {stage4_11[1]}
   );
   gpc1_1 gpc368 (
      {stage3_18[1]},
      {stage4_18[1]}
   );
   gpc1_1 gpc369 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
   gpc1_1 gpc370 (
      {stage3_36[0]},
      {stage4_36[1]}
   );
endmodule
module rowadder2_1_37(input [36:0] src0, input [36:0] src1, output [37:0] dst0);
    wire [36:0] gene;
    wire [36:0] prop;
    wire [39:0] out;
    wire [39:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[36:36]}),
        .S({3'h0, prop[36:36]})
    );
    assign dst0 = {carryout[36], out[36:0]};
endmodule


module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor2_1_32_32 compressor2_1_32_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h521534f7019ba947408991153a61ef2002dca621a3cd46109316c95fc81fdc8175d780eb3e2dca76c0ebd726e52f5e15a29412ed12e8bc0c233beb38a5c9cd587ac12e6ce6deb9a9dbe89f71eda2633a11ad9e69ee1b9c9949aef761bd641f6c8b6fe65b2b0f0f3277424fc2f5daf03546f26a7bf998e768f6a10baa94c2a855;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43c3c050fc49c83ca6db39af0e6a3d94e56a2327d9da2b8da0e31300ab71d283f468c4083094edd9e26308ad21f3db914ccee7241c2e8045577b60ca4edcccbd3bbde28e265ed69a0351c9d3d6e62cfae4696d9b20d36a91d9121b628571d6360e74584bac43719fcb37839a2b3b61ac8b98ba09c257ee9c59d9b43f9469e8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbe82e879dcf6919889a31c39b4954d07db66b8ca11afeefa82754c970052d59e28a8b32d01477eaaeb7b4a75e6311b694c4a2710717ae76ed96d21bcb677752aeaf0cd760bd131f00891fb120efc28ab053703985a9d81bc0bed7ddf5ae07e61c065ce1b4e946a4dd82c85a6da1d986bf250b1c8116b4e027d560c710310021;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80e598ea8d14326724ee253af83b595a94c16b1dce525f232dc95f0a8773dff54c61ca0f5460e33ed6d3c6d7349b2b6d735dfc66866b6ec20f7a91a6d4bcf90d3d84f3be923e876b565de224cbd50807dc67f2f4eeaf780857943ca8ecfc8e41867025d16813df0e6ee3b7e2224363bb7eac92c58082227585dea04376448964;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcef49129db3def436667b416917d72f50ea9884a96ce6d9b52b531f865c378f0e3d6d4c617ed07a23338d13e8432272a6054b70050abb4b20275f6b73be512068385b503111ccbbaaca35d584c18d2f16a59899cd0e8c4483311cf9c98fe25b48df1e12cfab4635edc2fde1f4059d163f45895a81a0fb3bd9c961d16f84ed294;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeb5ee490b45dba30f4ec91ba53f7998b5a07d07823a3b25a52eea2f94a7ea5691e5c4e7755c42d5ba546d119ff691ab42ef0d907b3d79dd1b12b619251842aadb5d27c2935de752e8102bbfea94b7d2cde40c7d1117c362f5176c5d89eb440d2e59b5ad907117866f68c462990691f750e40cbfd5c1c97b12674f332a759f67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fb30501a30b4c3aef5b897fd8f294dc22793c4a84a1594cb224a67238185675fe7dfc441ccf67f0600a9abf816bb484c0e40208ce9cca5beec508679aae70a3e5eb378d25573df0dfe97ab31513a98304ff51c7e2f5626fc9554794dd3d0a5fbe6785218586329de5705a6898b7a7e36b7ea8b6b9f5c8ab6454a9e5c0868b07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ec8bdc5ece3fceebfb7d8b690c747970d743e3b8b521253dff8c23fdc82d84f0e4706ef36ce08fdf75a23225db2733be014ce2b88bac89f2b77e2a3c6be63244c7f92b84fd36c2d4e88607f91b5c8da33c54a259b18fcfcbfd48726eca6642b5190c0dc1fcdbefab71cb4c94d33d3550b4cad0183a13e85dfffb3a6bf3ea1db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h413a331b1bb3820fb24fd893404ee9c1b5a9de3ebaa5f69e26f93834bf832249da2f24045bf4831e539636c9a422f94e33752d7dbdd8095b1fcad8da21c8af0d23d164f13fcdceb8e465c8153d0f6ea5eca6b23aba04d4da6a18216d65d6cc9f4161061e1a2729a56a4f4e2b929916a4514938879eb6c8984216deef53b0c1e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fabc2d85fbc4edbfcc510bfbddbb7fe4376d1cad72d749de198c1be2df253f4813bba5ba5bc2b27dd63e7ccd142325fabd0bc2290ef61cf1ae2b525a1ded45463278fef0c579909b18b6238c845a413d4d011e9bee107a74c4750beafa30e04bb885879857fb5801006302eb272e4af0d122506116bdce85cd8a3d860a11d76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5698dc6752aad4ff5ac2cfe9fb43e4b819c49d4abcd60ecb500c2f3e61b71f99820957375138fa60fcf71a4ef023c38ca2ce6310c3074172d1bbe1eff86e4843f78fb838de8225ae094eb364c1edfd5cafee6dee1217dd811e3daf9af92ab63f45783c60d3d9b6f377e2f0b9969ec6da2908ab4cbe41bdf6665eef804017ebdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac02c22946fd13aa05c63f52030743f2a4656a9f503802b9b0ac4565f8405ad9d7d1494f0390e93ed455d764f4fcd58bb5b92d6a118224b9e1a6484b9c6f484d50cd332c175314f1311c88013b9a917c7dd06a933c60d7592b6e0101e4e062f3a9779e8224c34427864395c1cde8b18d839da0ce80f39dce79535a0816ace4b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h369d5ecae1d5bd00fc454006d7f9314cda8b4031390478d69b8933fb5d3fd2e213fafc9d3ebe4e82ac0cd5937bb98f67623441a69887b521e4faca4b2c5c41c79bc1db5711d4f1761d759402abd82be3a723a529795abef53aff7688b07c082e17437bc3696bda5eedd78f69c3301801d24b10f1f379ed1df48a127495ea361f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a0261c5e98b14a64aa76b02a276ceb61dfd89f87dede031cdefe9fa071ac931f2f87f99de0b0c1fa33909b85e97d633a88107a622720040a8c7e4ecf6f5c73da24d7556665e2449f44b79870aff9616b3f2e378d5f4ad1ebe8d6836b19cbe16b011aad02feb55ad5a8fc54567744c6f5ab7138186818df0aa7ff74214776fd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91837ddaa666ea0ba5305afeb5145f04345910c04e0926ce5ef7e887ce938abde38d8aceb06ccad0f4af1080ae837472c1451dfd0eedd89ec0078e539f302da70e0e69b49c45431838feb06496fb339881723031d5fcb5b71a11d1c632e536d7ffd2ed977cafe092f0e0a8837244b65be68e61240c273e4054fa77b7cef9f861;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc360fc2dc408ede4167923d83ef51188614864291f960affaeef0f2113f4c868a11c2effc71418eb6118b033854d2b704a3caf254d807be98b502e72c5bd6d86c8e3a4bc61eb09dd7a78447270a7d58c3a6e1c7afd04358b575c93d63ecff29eddbd9b4d3627b387ab91301263c3d95a77a0b2e856cd3727921a8d6225a608da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5759bd7ea114da58f9e62ab838ea6d36c529b4b8b7f42a81331d355ca8777d337e6f319ecd449b9a2a9c14d844df0639429b6caaa27e90221ae129ed73b7895909f82057bfa8c7368e562f0fba09660eba5b38375c3caa328639a26a41736862b104c8d48c5613921a46bf2fcfbf2e3231050c827bd63c1099697efe0aab27e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf7d3bcbf55a76594a4b79b6f37f4ad92292737d9456e0781243eec59fd9e036d602574a8b35babcb51d10a2f0a91260f60de977002084a821f5b7b7df771668ac3103970392663ff29d9a478f2f2ac036f8a3b958a61873d1e71a4a9b2ec8d169c069d4e03524f835d35af3ba9879cb691150743d26d7c978af331ede6b3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35876c790d35c34e1acf4db8a1d1b4a2833f06254338678f0cbe5393d1f47f31b20f341e1ccac7554c35e4dbb45f4d03e4af634ce8b2cdc3ca9bd24713fb79eb5cf84479bd372b92da6c410e3fa2861b5e74ffb98fc18ff7c67ae9219b262e2712a8c6a06a4cfeddf05cd60bec1a3fd7a96ac7b44e4ae6cd8aad508ed404025b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2edc290fb2a71b74d153cd6806f58877cbbc658ce17ecf5d34ce81daf6954ea1ed594f1db5e12070d22093cffd76519c9ed72fcf66a4c0fba90e2ddd17d74a47b5b4d3bce4580e842debbb0f130fb3fd539c24e89372bed655b758ff05aaf3f8bdd7a05574e4b2216f427aa49735433473eb01ac37109e8e4568a168bf8e3b89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f4e4563e86d30146aba06d1c833fec44b92df9d48cb0c2c760f37da1103a47813ce065646ebe354353debc39d87eb078082b090955e1bab58edf9870e005cb997d36f56fb4bc61bad7822affc97653b0a3021959ab7f5f51677bf773a7ff12d7437b4b9785d3a851001887ec30cc5754db6e64652a1d32410e13db9ad992290;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd61dfc9952b86bbfd158712a809d62ae9f0f5f70862af6fbb5b87f47df73cbf37a930516286b7d14ec5d5d780f9140f5c656afcf1fc2bc7720bd615a6e2c12a1e4ae68aa98e392fcfaf9e5fb43488e12dc1fab3c3089a1c58d350d44667e429cf2b2ff7bb3a2297e1cf6b841c9b1305aed9181d7187b3249a8e4cd297c9e6bdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8849e10dad41f78c36f336b178b15ec340e694cc2b12fb3f86102d195e13b0b18226332f6ad8e605fb26a0bb9e192ea973b8aa9d0c5af88b35c44a2d583a01ffd21ced60123e501be6622159c6473494241e2494b47855bb42324ec77b06f6442147ed5191016ce3a02b685a79390698a0d1843d568db021020cbaca50fae07d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b20ebc54cf86fe251bfbe9a351f2952ec9c7cba70e6ed91c6a22ad40975936bb0dd4480e2e6b2af1c452e6059420924767b57f9deb1a00cf83ac333de6a92b0428fdb9c7aebcebeb1b5b97c17e151ef3d3f65877f83441fdd9da8f09d929ea8a51a6223fb84ff47e34046e13352970beddc85468fc2e9e22e6c1336d4f905f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb000af4a33f687700d42cf83b725d833b374dea2962a48a993190622a235d7547acac031e50ea276da6314070b754fc5dee203926d05e2d1360263e3de78b45d25297bf2b37d4163430b51d8410e15460c5190c306ff5a1edce90d6eb8c5ed37dc523e067f2a94456c3b0b8bfde54650a3ae638cad655defe37f0a8f80429d13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde55d4f949b506ea0ed1a4241c17fcc10e47ffeaf62b2ce76ed7fc0b6e3b2e86eee146c9f7c54b6bb037e48901d2cab8ef43ee4fbf60787040b1a61eec38fc5e854ea74e46f6cfaf3c6bca724f61f52fe2d4ca3e8e4bc2d82cb927445fcf5c877c1dd218a3bd757811c28ef051aeadfc35fc64b263e4e949f6a7c9701286b72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ff7f4791dd871d91d26cb8e95e5bec7c32164f324f76cb533bd1a27380824010c352a1042f1ddc353dec7bd08470c2fff30151189ac7c4517f796cf136a4353350b8118408cb1efacf4926afe61f26796e57015ec931324fe77618e46bf000c1379d001067d99abe45bab92e4fd42785b3b34a5efc74fc1d552bfdcf5e814d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74d60cfdba92b91ff7cd85a991feefc840d5f6986c2a5e5057bc4c9d4f8e6665a1e10c97391b4fe203b7fe3aad581d8db69c3e5ca240aa5c88d68c777a3b4da09c038458dc17eda3ee2d67895d7ca5ffd7662a6a601d89c4dd2e0dd9f9cd286efc346cd2468c0b57c3d6b729004362e04abf4bf1431c85523f55f3e5f2af1839;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd0ac38e6e0de19139cb1484ba2b49130e6b41cc40eba2c511178a30f4b342e0e9350e53d8069df5d93ad3481f6e442ba0bc7319c8653cc4c95e42d367a7c292df48b5b9c373ddd0988bfa40b41765c30f43f98babd6e617fe2c606621865588c16caef978068a03ea432a2b55d874d396ce0837b665db4aa94da0e3b109e47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b16a4327f7aa62c15fc59417b1fc91ec689137ef11e2aa93193e1dee6661877b8ecd1fe0751fec4343169500d6b81c654c626ad954ca56e072383353f69b69ed9ef0f81071e4a2ca7b9833d956f828b76d5d026e3dd39c713e94104af728c2f763a703e455150e8e648836b13175203ba6a812e683c4d8ecd06c539639fa0cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdb19c376d57018edd957bc221b84aff3bf61590f8b2ead1fde23f7c752830c4760951b37e9b017910594f17fcb9c3bf5fb4b92052d9cd0c2853a52d99aa18041abb62c64fbb340f8ce7eed5af7b59b577aed8e77b3775952af33fb8d727e74cc5dba72d8fd388aa8ff13e719bee1799d308ea75f8c483accbe9a88da249fb2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf89dbac59a19c8460b722e9c77366ae99d1921b08ff25376f2096f237632dee1d53337131c399577a528535cc40d9d0706d186f766ae187144defa65341bc06e3c2cf7e74f669ddedd88dad8f0595f0e1c26665c63a185d93af4daf4d606c70c8ae3dcbad78d34bdba3b5d125f989654d0c0ac2a96b3e90695891215afa40c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1efa07b0aa54006d8a2463d9da9253445fe516d769f875940e9d90aad21ab8ba2fcb8b025cbf8322ff0cbaa4b727be4632acb43c5866acce9dd864acfbeb76d5d79657d63f1e70f7cc38d103c95d52c29ebbbf01332245240c9dde136c53fa4cd828ca2a235b0818dac8cdcec0ad98f83559a1724675338e0d7534ef4c4a1faa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53399ebbceb05aaee476563adfa7084d9d1d8ee86688d1de687e75de138c055e5fe62fd943b48c8c0b0a4e142743f422ca3d1011f3ed031cde3954dd27c4a197788c9caea4cb5e38eacdf7d94e6fe9037f7b7ebc6a21bd47da2bc4e14464cb0f224e6585d23a8812e39f4da5f014dde670bec845b40bda7718b0b22365438d84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72631accb60ba9a2c7b8863fab497d40018be51e2653363c025d99181dd30b6ea083e472f50cddf93ac8eac84a4cc506259185110baf6a41a3947018c55eb8f36a0a1981c2dabcc50151027c027e48ec4ca9ea267b5a729bca035102a17e3719e83d2ba4714672627c25fe77787529e4d806933f7e4d7497f5e696f097a3f45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f31a7db50dcaa2a8c57837815e259ef8ee9c6d1e1d9b61c39c8461f4032144a8606d111fa2847d38c02d301bdf871adf5ec66df67f3ac016611c3e3aaec22f73c43ccb828e66eec9886c3656ca2779646e5a62228f87049fd896db4b2842c1bb1383b39b7ffe1bc6ed4fadb4ee419db55415ab99ab10ff7fd1f357cc896b3a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73a63c39b324a6921503425f7746c73cba16c569e969f2ff3af19630840f858923f55e14c19a8aeb8bfe5487cdcc2e6470e71630a7bf5ed53e0dc7dd89f966e0dba42e55a4d7d8adec471ddf64a96d70691b943017ac4a1f019d30356852545447b551d6635e904bdf031ee5ae92e72790baecdd9d0554682a26cb053d8e4fb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h656ffc616ac29e1057464b4a496f93b9b62ca237d06435ba82934abd7097d3cb13fdc960054adb089947ac45601edd3cbbb590cc0b524f4a06fdc95dbaa2edc0b2fb8ba29665ee32e88f8bca229122cafe135fadd73b286fcfc7e057237e6a9e11bc7e717256e72608c71856eb7431bca14e35d484d9e7b6d45cd0221c59848f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd086185954b8862c534a15e73ce59c698222dc7a68036bb8fa83576d0517adae6d51fbd917fc5ca86b0fa5b865acbf347197100b5958ba167ba08c0e774b7687d5f39ac97b8cabbd7ace36bcc4699619dcc7138de8bcfeed330a3a50f391d4ba6169d7a5d097495d339051f1ec02055680da47a54934f9055d80aa967f2197a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20ec22d9c4848da8a5cbb8cab89396c3ebdda9db51943ade89477fbca38856a3cedcf8b3ca11437edbe2ae6f001033596714fd68039cf2e1ae652eee3630f41cdf793b7b4fd60d3ec621e1a4cd6c41bfb33e06644abd28846176e0e5bef624436cf0a821edb2661832bc85961b38a7641420ee8cfd2f40fd4356a8fe7721bd26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf98d3415821c2be8953272526572f3177f30d5433b0ba9c9824f81debaa9bff287a4b7c322382d7e80ffd0c0e439245b1b20e86f57793e0ed0cdf6632caeb7c4b40eed66fe1ab3817b30b8aba5cc26cdb971207a54c8681ef2ee62d14ddb4897410f3765683676bea0dc19191802dd30e0104121e368d9c49aa9ee52b845645d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d084655eea07ee3872b67135cde5f333e43c9cfe199e89564ade57e53c1f95055e7f29fc6f786a663dabbc62ab953c5f17242b5066f60b03430f1651251352c99277dca589ab02adae826d384d98d472cab6c99d271db9d28b14ccda52b01d02275622eedf654c5cb151ac8831a7790d798109583e78c863a808b78f7ecd5ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h507945b368cc4af7e11e53d81ba916aed834b04452db4dd888065d5cbd46e2fc3d0ada7c9629ddeb54148a9ec07bc63ba8f6316d36993f977c8343413ab1bf264340d9848e5eac13ba3fd5bf9b7ac2bd59bee9a19bfe6fa349df5ee656ecbcc3926b2e8086777d6c5ca9660b4d8b5eb770860f45dff59137ed12d733c444e3d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34455f3f604816ce482da8a93522642f69bc8c7aa3a3b9da4cad12d0847843203c92c69b8e5f6b1f9eff72cf011bc20aab265548f04d9fcb94bbd6e06d45324b787c3fce39b18807a5374ae2616cbe1772dafd4b4af73710787225e6f2474cfb8eddf6f9e7b30c6274225a9b10ac9bd62bd0b10452f2e8942f3fb98f6d1b82a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc155d643c1aff818fa47b1c5a231c5cdcc8d06273ece507db8b2c5ccf91efcf0384bae761dd08c4b8d5b12d709f8de4f28818f2834f06b09cf5aa7ca574d027a9efa8df3287bad42bea00cff875588be5ce7580d18d898db907208ea0206e4bc4815faa2b509be0c50279e36fc5fed0cb3bab5c54ec45cb3f7f002195a0e17cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21f9bbe7b226681488cbcd103b444cc44d7b1d3458a3c6994f0cca012020ec7f7c2752a34af5a27c1bd2639ca3cf8a702fab9dee2371374535dc36e7bd7ef0cfcd23f10c1507adb219c76869e66c1acb059aceafef0cebe7566b5cc4199d424f2a72f52a3ff36d607fc7e4b841e16cfe5d604fd52b5258de9d5ddd50c403b37b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb1226b1840292074d89213b6806be94f77090a72a7696f35e11f1c89f9f0fb6518d8335345e690bd9a099cc0145bfdddff07ccc683879b6399ae86e1a4c2a15f6486af723d11d907b074cf31471f2632c0c3882dac5a06683fc90c52ac40e171a5b1bc33bd1c234955bb61b42fb042c7c4912016611489d66d3910c8c62ace9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8255e258fad5555268bc9ff92d57dd1a53aab05147eccae5718d29d222d1979419c7d56d027aed427a46ff8a107322b18188b3d044ca8c09f1473855ca92fe0ef0b93d68271239d8c9b54d6789405472960c4170b41039a1f2b135af2db5e5666c255aeebde2e2d85cf1b6566b9bb9907142bc517050473ac95dbd060be9fb52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0ac2ee463a1d85e1cf9a30ddd1026294189f4afc7d509bfbaf8b83b9b1b92a94e20eb2c254d5be9e701283adf5110e550d8a7e208ad77037596fb4a5ec7119a266b39bc308f1718d7f52c8ea85a1e5858dfce40cfd83937092eb16fa5eede76d6eecee630c12f32d25e01b866dfb027951e04dc4c0879316f3ba05f08a0fba6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd19b195cdb6270a9c6fe7ce79714e9ab21587094eac7e0df51e9115d7434ec21a28ad8d938fcdc74d30dcd568c9d852b5a430cb6b0754c809f40d24e84d5927ec3c22b04df6a6d89f3e184e56b52ea79e8e180cd90a27c167944d6269b2bffb598739c240d15ac622e220a96c25ec38fe520fd707e79a83ec28170c41c2e5d75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a7ac16ca1620e418d41b2c7e782d577a6b99ebd3c5183d456f865b9400d8b3f9ede380f74d1423369bff3e3552f63bd99c6093be86086c9263acb644f47c55a843e18745cf02feb604c4139877e3d785734856a0e251d29f1dfbb6a5140f51da263b49c055d1b2dd2e9898deed9a0413dad20e20f5de0794414d766a05d4c96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h353e94221b076d7f411fff7aa2d4aabe8950bc4885d3919d6f15972dc6301c87dcc9b15fa240eca9ce165daa44b41cd1210137851fb569eeddf1e027b3a1de99e90c2ca8068a43122a9cebb334341d5f3334cb8ac14415580a246c40a65bc956a14e9edd6f86607d5ffe0bbd85e8256805e58c0c5d5d2fa0d5e35b78d1c5c4dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d9668c59f37400ca6f6567ef3c8892bec7bc0a851cc942beca4c79988e855cc703ef502e40db9cd70c0316ce0f24b06cd606ce2ebb8c911502bf76d2361c933c4b65d9d497eb9e7946cff69282493a645e80a498a072bd2a6d0aed06270e3f915dd9387454ac81ecf6c97eef6aeb5640c473bb2125e7308cd5309d63bcd6f0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6977ec9fedb76580d4c7199385cb81a22eaa51a5fb73f39b134f76c43c09de87987d564fc7be019be5573b5ee326bbf0513068e9391e1a402549ab77e3e8a552e49946351f889f5f404311cb6a064f4ee4f35fd536deef7bc930a34dd96cb12257176745a21521d018bb8f5b633954a128a41bfa95d7d3a0d349cd2d3912d05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37cef7d88974d92bcbea4dc3a6a5317514fc60c0c4cc504ceb69c8938dbbeb4a5b27f1be440a2f749e2d3ecd8ad6492bbf7311f22411c626c3e376906825b8cd4d37c369cdeb886b51074d5e567b7854f9ead5acfbb8794db49c263653f774b17e294792f0150529beae16f307fd72940c127e2ecd49083bc8f46b8e435aa944;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b243dfb1ff2bd30730dc2be172035b5064fc913305c7d21206ed33480ca99e57e85ddd7081c757acc1b9110f5c3883dd7db6cc18f4bb7d7a74c9c384093c7b532852184dc72735614fa9bd768d29a2511b7fcf4b862ccd4e13ef37aa2bb0527c12d62314951067d6d2337d8353ea4a2e46b936bf20369ba1f52dac49582768;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2ffc05333230f77955ba90f3ed8f68b19da2bd514454ad29ca4adea0ce59b79431b69e47c98c291187aa64df656a79e9f1a281a948dd82991ab5813194ca9c010acee41734f9847dfcbfbe8f5ed035f2bbb36425fdb3d3b99450af89239d7d2ac86f4906c1612e1836b77918050ac04765b6986be0922e5c9a80461fdd4c40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2241e11c577057b9c78acf3fae75e3996c1505eb1799ae6357e7f5a62285024ac5d54b10994747cf48f8628bf18a183ee1fe7c5d021da261932dfea11dacc1ff479a8c4c5ddbb05a3c7f7e6045541eee428f5996e2b7524fb7fd230cba170c3d0a2617c5eb17c77d550fe16a73f779cc245792ac61a04f05f4582f92a77d0662;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e1a33e5dc285bf3c72b7acd8fa8ba34713b724df1c299adbed0bf5ce01e54edd0fbc7035b3e161474de108e63821268ef4e891177561475ad926309933d3ba38f14d41f3b953cb111e9c81399bdfd60bc5461c7cff4b378911b021780cf8fb7e63d19585d44ee6f2091c975162e2e39b81aa81dcdc5ac7de60cdc68611b2cbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb81b5f6de16934e9740d8a122d2b6ce6d876ca4ed7056e74df5924930d293c56b68c29a0986fa0efdde5be529ba81fd7c4b57485f88a25f36f82839f766744a3966fd07cc66072104dd8d7a798d907966cdd8c90908a1fdd069da9db9ce1fba4828f2fe29cd400e0594196cf0946ac33e0a7d7fc42ac78280e05a4c2080db98a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95d37570bd9bffbdfcf7845ac7f8e49caee325e7c31f287ec28375c9bcd4e5e692b67b3d06a631ecfa979b105a3966291b8f3f35c7672b23539fda7493d7cf4294360c33afad39e36439e34063766bc93815ef4d2680901c8899eae9d24f83a0b38eb15205a3dd1d5daac37f2be66f6f32fdf1614addd1551de5477989721379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h560442664e3e12f12f23af8906286d69cbe287d1d27e12c60596d7ddcd6f99353d169aa7ce1c5c4fe9c34bb6cb7e9f622a4d4301f48115ddfb55f96ee094a1571d0089c46da04c7045a720f98758ddb49082505cd9d2e845fae724d10184aaf507da3754655e93510dd8b9bd3621128cf6d31c93ddef283011746b760b7a3c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87fd90dff6a51ffb897a2b7818e8ad36e243c7c7a8595e29fa0f510173310541b125ca60a12d5fbe7488f8ce22db0afd3dbedac4d15062f15ada2b6a5049e704521a1e0efcab6d3284944f7b744b213f87697d26e8c522a0b2d1235490b231eaa1a1be2df558b550a28e563ce98e052c8a872b215e96fc20383d551ee3f4d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7d716c48a8cf80e5d5e5d1d0d258ea985a6eea6a5f8114779ee29cea1c715356dcbcf5961af546921892518e9767ed3157606482556c6f6df678261a6a03e4ef148ea2e45595119a0dfc7eeb3c65c1850dfaa010187a14911fb35c473dee7c0181294dc3fe7ee110acd2389bb56e3d3a6372ac7f91ac9e827301707b9f6bea7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he40061233eb12b03fd9c48e7b19232ea8d065de1043105ad8c1a24df9ecda65e5109785ed116103f468c38d7a96912695a76879462c9d95cc8c9cb5bfcadb6e87955e47f0a144696c2c2b148937c160e5964284d1a2c411095831f50a3ae243272367f87911a3769d6c92ffb67343bd36eb9f7994ffebfd9de656665b3a619df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6da82b8c1ea1a3c9e47a4510c48c0f332f654c2c35059e6685f84d961079c3f70e9defa00a8a544a8fbac8694d23c563111bb16f6696e2dd5f714155efa3e3f84e3df413914e5a207c75270f7c286eeb6464edf1e4fe62d782bad5db0d50641855bef8cfcaa75c39bd61c7fbdf819964756c7bfd8828b7cab8a53b9eb0e1abc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha66a9a338e23bf0751466d4be0a42bd3ec9c8ceaab702b3b4fdb50f89a32dca8326f5ac68c5c87a18c07a96f25ea2b6c9786373df0a6838d87a6b7be85547c58b4f40b2d239329d299e50387572049d11d081388409bd190282a39525e14313596ec5556343a67e34f45a36f089be9644e3bf83fd553f9148af060752b1a963e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h823463fb5d26175e227c99d4c1bfcb38dd89ae7741a1dee5cd25e890432a3f0cf1233159b10676db04d897eb5feba783257fe7569ca434e6d7424ea6d8eb4672a924c077f32e856019b5b3d83bafe837da08950b3dafdbb878fb51cba0bfa948065636374a7415ef3065ffc1fd5d956c85112f95cf2fe710b4bf3399f14a2eb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97d010a36f103f71cf8e7707110d6d037f58aa9ff2dd4a94b5143203a9387a18411eb29f6a8232a4d8b8771ee743d0a0ffb3c9e5a55a15c0dc9655773d74da1d14ff63dce5a37536d986cf7e1b3a88d90f23ed50675f239e8306d9d73f95e6245c74698e24eb0a73caec4c8a51e4ff32a2cbad169c0e2791de5883becac0d3a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3607cd4c9c160b9a6b5ab5d816fb947d4b538dcdcd6e38231f62fd47da92a730e3b160a23e35a9402b14c44d35311e84a0492f102f49a285f929224a52681e875092fbd533b5da7c8e61c62bc846695fad715afc8ca0f4eb2ca1f2ff22131d931771ebd474ded2b4c8314d0e9ef9560325bcd1f886211862a62fcc432a648f18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h665f387f828ff8c4b7f60f41c056d34353fd677c15dc7fb1f32664add745eb26e994b15303ba669e3d36d6443974068a58184c3b592af50c6508c60c7bf25e1cfbe90bc8d045ef6af3ae0d242d96cce88e95bb728bba4461cc04598e7fadaf11942dc77e4a8164ef9f8108170bf4e7cb3a7112bb355bfdb6fbf74fa3dc694fda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heffac50a154a2a76ba43d7fc2fe3bc52cf7323ae98749ab9a61eb5536b6943a393478b31f0f47c6a70fbf0c23487f5fe682476ef8c6435f076260310f3e5ea786144898ce301a5a213cdf05951286b4da60d0c3d9a3424cba8e82c6b7730773ecf3ee7c6ddddb61969a76f12aef8475e2a134517fa040da5eb57a7af31a2e7a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he55a23d3e3f49c69dc5db53591e98af8ede5df2520d495f5ca2fa820aa7305af1acc7ac43d1be12b34a7746578fa4008d2b4ae36a6affcae2309d93e916b3455dd6f54930f3885887c0eb5df07d6acd2df9c7b61de5070e2ab986cf93f82a1d31df9a44522cb47e5cda83ee04984c264387348315da5501ec9844437a3a17e56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c22f5dad53110590aca8974325613e6b7349c22e1d62fc4f575182cab3e94c913f00c505a8226f5d5e4fe293fd5d4a245ee12a2fea60a1bd7e3b3b2fe97487b78f8b80c3df953c268ecf6b9f800876d5046b37e65fd1a0741987f9bd27f8114b991d7b528d05e5913ecd4b34a9d7e02fd5d0a2ef6799b5f9c26f090092ef7ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee2196c7658ffdf9bbdea264febfc159fe8aecbef6344a857c76ecf381fa0b7826aec371b07288f273ab83a3ab7d6e749a11c14eb6cf33374de11e3c70c9717faf85af948036b712e4fdae7370039e1ca01fc2075bdcf4f14e8091426181b54114c770785b53283c0ad81b0d3bda44658f0c5eb5623357cffba555b1262edeb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4ee84e1472cc546d5b553a1948466e7091b18e5906d5b6383d202e7f821df4b3dbd71ae6c0044742b30ca24723a1dacc23ab108c0886049196a26ccfabe3417e9456623fd40203e2363f7f9d1dabb44ad5c1e43bcb6095b478a89e3d61f1db67b16d1ae06f28be7ee24aab91a037a086fde0a19946f2710f0c574acff328866;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54e06f7f7989ff264ede3b058cd14a28fe2ead4c6971ff7be9644732517ff8d2b458c3849be3888178d741d08b391db314b315ca6ef32b5a1bcdd091ee07dcbd5ea5729a183a3e9d931fc07a2f8350ee8c81a1a3241cd396b4d56e2351639490d6d4b4e47260c9e21df5e442fef3033e3b3b410e51ecc2741f926f4305ae0547;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ed0d8f6c2ff51c71df1d5c21da96bda7db343050af420e1b498b7b26395ab7bd50298d96f053575af10a0a5e6b9ea2bf7ba9fda7b697812232bd0c774427516c6e2c03a6e8371064ae844b7b77db59518cd7cb7dcf04f2b6106e45d3bfbf0c5ce870971f7dce4d00310fe44aecabc91534d969e17e61c106b0d2930b3044685;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6df9e1d4068ab6edaf7dcbad2128df51c49c933b37a3b931811a3c86ebb9d9f3f7047737543798b16a8c409f3224d8db0a24924d2dc98ac5d605cf0b2ec0534bf9c0a091fe1af8057739048b61eaba40ce11a842ef47f2c76649e172744b52f60f87c11df9d64be81a3fda07b50ea2f76a3c5ebec7c5d7806862b9cfeaab12f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8422fd04d09d8184b4c4edfc7c8975f58ba2d43d9a7043f5dd75cd3c0f6958f5672fe0a2edca86636cbe336fb76ec349a9621b87d1ba6ae4f46304b163a110ed45f2aee7bdfd59f4c743e024a91161bf5e28afbd621be1730f7cffa3a81ff31573538c840508ab0a6dd663c14b42a628b1f026f125d5098372ac22a5a6233dbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2d54ec7577282764b1a09f5bc8f9141b0940dc298cdd55d77067d0b6396f8e0fff8854eafd8ff9b4093198c81dfc202bd2214086eeb25e56bf3be8d60c570cb13d3763bd49ed12e8a07065d956c9fa7dd57a34f0fde94e3333cceb5feae1b1ab0c72fc907dad49aca34fe50200278090f1f731b5ccc9457351ba0fae899008f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32a049947877e224ab53b24a0089480feddec837381818349c20e96e2090461cf7eb53f44e1bda7338da847e31ed91f5e2bc4384e523d98a784fad9d5b1be7d8b13112bca3001083e13da0f56d26da885afd26d9a37e10da25703f3f34fa7f6ef560401fa512fa215f10385ee9c4bf93bb0fa94e71e9c27f97b6bd28e7be32c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2762e021c2b1688092525ecd7086841bd25163474b7ec15d12d3a24568040927b876e1cf303f633ee93987001981c545ae432813c7651e56cc7a405d03c12c667428e4f8057b25eb9090104b7466b799d5d0e0332b0fb14bab8c1cddf220b756cdf69e96ef092d68c5148fbaf1376f1505978d71744d83892727abebac4afe9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h901f70024148890b8f7b3f68d8948e84fad11bab6e5cb84654beb53d28c3888d07924968f4a2b085fcff2580b802cb28933ee60a36c4c353d9399451662aa7af635d709abac9836c2bea4d97dda20c0dc7bd6c4ad881ea1183b6dd5a520fc84dc03aaefce3834ab4f592757127df247f133c11b1c0ea630de4037901f3d2cb3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1cd10ef54d32ddba5f4c148138c674825becc7a93eeb0d596337c36c3174c5c3c640270ddc7bf9b3df46fc05ca8a32ca161c3053430b296d5fc83337e8682086ff576918ba867be30087fd1c43d4b5a37b355108ae73db63ecf6480eec84540ad7d9f0c97de172970b372ee21549234d82cff17105ea3462f36870d6c194a86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h318c011fb52f5d33bdbeee1c3224a5673787d5a9d2a83086ac0c865272ac607957a6ad3f3553b4ede15a1ad3bac33ef5010f2d06778757da9135c4a2ef6a83b5469ea813ce9cc8b5f2875efaa63bc07cbf7178e714b3e637cfd0f724e5e7c3c042131724a1cca232f7dfc4b7d5c64d68fc69f91544784b54e6b241249ea6b646;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34f6fec4282a37099af6f3085cfca940de8ac561adfd612adb333223161fd523076d3404c8819b2bfff4c11bf0892b8df5edb3157138b53fbfdb2e03e6bf0ca763ecf6169b757b848115bd7c22b924a0a85749de9cfaa401d26e1485f0c31e360f669e44c9a0aa51d4fc511d0ab0547ad4271669bd9df327c6462fd05acb6cab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h963957c93f7588d7186924f6c02143173f17a91f758acbc97dfe0d44afd56a7716b619a2745e11648f82913b92cf1f52998457031470cc91d603d7ab4901205b7e4c7a5f4909f68394731a0c71c2015e3527b763c2ee00e1bff7efa6d9151c284f75e717e73ea512d448562cd403ab6914a4a38178a50c5d1187dbb5d963cb8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66be8c9d4ed9ba5cef250acb1e119dc46ec7398c7db6d7529570eaa0bd542649b42457aa48e3d68bc100df96804c7c75a0e414749c71b3888c316cdb93012134ef517b5c43b580fd870bc1a52560c696d401d888d9e2fa03a727863e5ff5b5412ddaab854f2f5f0a4e94447923370eb063a1b5d0aea131bcdc379b96bbefe75d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d12c1612bc83200b27bf8cbe12f17f2e7ad340b2904851797e3dd7b2b4b7938dde4bb3f58f5dc3df533ae7dc4c20c65244ba93feed729d23f9cd835fead5147a19ba90839b11c05757520772274804fb77cc35b1341dcc3e008a7bbf3bd5dc9a722c29081e76269d161e1b198fed73d73ca1265db0d16457f4a28d67dde4db4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94319e7d75e598e7e8197e1335514760161c4ba7676a900b64dcd3fa89abe799e937aad6d039be8a8fa9f4a54f297faeb9bb0c0207a6eeb0de7fbe1d96a5bd8b33285d6a446d20fe19195653ad5bc21c19f41a39b596cb6d9c7f51c84b739f4cbc3f02dd591b5616840c1db372e8e669e113bc354d897eaff1b7009e00466369;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1575dad2b19d486d499aafedcc123730fc5ec53378e5f079ae982aa519093a21b461bba898b81cdf386ea1903861ac5394f156d4eac75cc5f1a601f54eba62605389b5e4a4b80b3473ec1383f8726ffd91031d9a1dc810f9c1b40a095d7e0818998784f7b67042e2f29dfeb7f794939fc36530735373746590aefc2f620de827;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dc9917e886e9d9b41e9a19f42668760f5a027c5bb57c49c07fbd1a57450949ee41fd25331e70afad3bdb3ffe8bf3d8976cbf8540c032abad9a752bdb325435858e089c17ebc38b7d5b8d0649d9d86ec9bb732d288763202750a8695d27fac15f2ec1d6c04b130a056954fc1649f47b6be0da45e43f806c8789aa81f5afe54a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dd6dba7546c974471dfcdd7477db82c925b29752bba0f14c9c03cb7154e91a21e20eb96a9eb11b0f62e7bff365f1864629231dc9235c27d8e70c10ebbd7c470eba2519011ddd025f750789c449b7cee4d684972a762c254f0251249af77a85b0dd52c5bdf8a2d64c83ea2c73c14a874c3a0575f08fd5c1a653a2090b8f01ce4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13cb201088b0af21ac24d0c89bcdf95c4b619f58a6de77eda7375acd9b2535fb7d015a36d7893fa34b5cc460208532610b4b11381a724e8dddfbbb7473f101aab0d0062a08be036ff86316274487b4dbf3137979df6e1c7389e749c7f6d460e7831ed6e690e8a23564098ea2ad61b08edc7996a54007bd9838f8538bfd25ce7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55650d8efc977dbe3567c1171ff02930549f2ddc026d1b275e456f442c2fb1854f4e2013530af59db5cbdfc10b6081bb1f13857b85c0b76f132646922f4fb51794d727316206b8e6176488baecfce410c7309fef1d1bcc1e04a8b484ed4612a3a743fab2835c70cc0ceece847f1276529bc239bef4faac9b49c8e4b63d6d9ccf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70966969621ccb70618c66bed022da4a38530e98393ab672c175bcaa719038b7a6dceb611f288833b118a52e8c362de792563db24029a1e4b0bf626e742da9d032a1adafb8acb8d47f60b295632621bc8a3ab4448f93c9cd34679b44d9e20fe6be02ebec6771c2b57d81b16851eac59275dc112d24dab31ee1da6ae086ae3023;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e468c85585d0118f4ab39fe1398ec63d4f4c8458307eb4416ed83e38311e38b74ffff34b1205fbb40157ada3741192f32e76eec352571236463aa25ebdf7b6f4d5d4da373b1aa5eb830714614938b14b4f5627248a31f8646231007cdb35390f9ef94048b2ae3e25d9859e9701bccf39eb3393099a9f2eca2da6a44bb014bf3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c9f7ad9e1e2e46922e7b5a2cf0f1b1ce444ceb912437f2f503f022fefbccc452ed14032f7ea6548d8f34b3ba42aa4ce640773535b7469fe6e20135dd2803b4eec3e99f8f802b6007fb2374a533f2ceb76b3102c2e0988fdb3db65398c248e4f2e9d74290a41e2d82c1e2411f4d852b1c7840fa21e4e304681538e950aaad79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f51bc255d53937338ccc2e5105ecaac8f51952472ea8347a32673928eae06e019067c774814af8a9f977d3121f87b3290fbb2af36ce164e89772b67b8f9831f682f98bcf37671ac8ba097db1360e3b4cb13fc335a7bfe230041977ab0c9583655b4f568e21652fd845b5011087d4340794adbdb51bf012b54f5ecb6cb89441e;
        #1
        $finish();
    end
endmodule
