module compressor2_1_162_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, input in_data128, input in_data129, input in_data130, input in_data131, input in_data132, input in_data133, input in_data134, input in_data135, input in_data136, input in_data137, input in_data138, input in_data139, input in_data140, input in_data141, input in_data142, input in_data143, input in_data144, input in_data145, input in_data146, input in_data147, input in_data148, input in_data149, input in_data150, input in_data151, input in_data152, input in_data153, input in_data154, input in_data155, input in_data156, input in_data157, input in_data158, input in_data159, input in_data160, input in_data161, output [19:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    reg [11:0] src128;
    reg [11:0] src129;
    reg [11:0] src130;
    reg [11:0] src131;
    reg [11:0] src132;
    reg [11:0] src133;
    reg [11:0] src134;
    reg [11:0] src135;
    reg [11:0] src136;
    reg [11:0] src137;
    reg [11:0] src138;
    reg [11:0] src139;
    reg [11:0] src140;
    reg [11:0] src141;
    reg [11:0] src142;
    reg [11:0] src143;
    reg [11:0] src144;
    reg [11:0] src145;
    reg [11:0] src146;
    reg [11:0] src147;
    reg [11:0] src148;
    reg [11:0] src149;
    reg [11:0] src150;
    reg [11:0] src151;
    reg [11:0] src152;
    reg [11:0] src153;
    reg [11:0] src154;
    reg [11:0] src155;
    reg [11:0] src156;
    reg [11:0] src157;
    reg [11:0] src158;
    reg [11:0] src159;
    reg [11:0] src160;
    reg [11:0] src161;
    compressor2_1_162_12 compressor2_1_162_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .src128(src128), .src129(src129), .src130(src130), .src131(src131), .src132(src132), .src133(src133), .src134(src134), .src135(src135), .src136(src136), .src137(src137), .src138(src138), .src139(src139), .src140(src140), .src141(src141), .src142(src142), .src143(src143), .src144(src144), .src145(src145), .src146(src146), .src147(src147), .src148(src148), .src149(src149), .src150(src150), .src151(src151), .src152(src152), .src153(src153), .src154(src154), .src155(src155), .src156(src156), .src157(src157), .src158(src158), .src159(src159), .src160(src160), .src161(src161), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
        src128 <= 0;
        src129 <= 0;
        src130 <= 0;
        src131 <= 0;
        src132 <= 0;
        src133 <= 0;
        src134 <= 0;
        src135 <= 0;
        src136 <= 0;
        src137 <= 0;
        src138 <= 0;
        src139 <= 0;
        src140 <= 0;
        src141 <= 0;
        src142 <= 0;
        src143 <= 0;
        src144 <= 0;
        src145 <= 0;
        src146 <= 0;
        src147 <= 0;
        src148 <= 0;
        src149 <= 0;
        src150 <= 0;
        src151 <= 0;
        src152 <= 0;
        src153 <= 0;
        src154 <= 0;
        src155 <= 0;
        src156 <= 0;
        src157 <= 0;
        src158 <= 0;
        src159 <= 0;
        src160 <= 0;
        src161 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
        src32 <= {src32[10:0], in_data32};
        src33 <= {src33[10:0], in_data33};
        src34 <= {src34[10:0], in_data34};
        src35 <= {src35[10:0], in_data35};
        src36 <= {src36[10:0], in_data36};
        src37 <= {src37[10:0], in_data37};
        src38 <= {src38[10:0], in_data38};
        src39 <= {src39[10:0], in_data39};
        src40 <= {src40[10:0], in_data40};
        src41 <= {src41[10:0], in_data41};
        src42 <= {src42[10:0], in_data42};
        src43 <= {src43[10:0], in_data43};
        src44 <= {src44[10:0], in_data44};
        src45 <= {src45[10:0], in_data45};
        src46 <= {src46[10:0], in_data46};
        src47 <= {src47[10:0], in_data47};
        src48 <= {src48[10:0], in_data48};
        src49 <= {src49[10:0], in_data49};
        src50 <= {src50[10:0], in_data50};
        src51 <= {src51[10:0], in_data51};
        src52 <= {src52[10:0], in_data52};
        src53 <= {src53[10:0], in_data53};
        src54 <= {src54[10:0], in_data54};
        src55 <= {src55[10:0], in_data55};
        src56 <= {src56[10:0], in_data56};
        src57 <= {src57[10:0], in_data57};
        src58 <= {src58[10:0], in_data58};
        src59 <= {src59[10:0], in_data59};
        src60 <= {src60[10:0], in_data60};
        src61 <= {src61[10:0], in_data61};
        src62 <= {src62[10:0], in_data62};
        src63 <= {src63[10:0], in_data63};
        src64 <= {src64[10:0], in_data64};
        src65 <= {src65[10:0], in_data65};
        src66 <= {src66[10:0], in_data66};
        src67 <= {src67[10:0], in_data67};
        src68 <= {src68[10:0], in_data68};
        src69 <= {src69[10:0], in_data69};
        src70 <= {src70[10:0], in_data70};
        src71 <= {src71[10:0], in_data71};
        src72 <= {src72[10:0], in_data72};
        src73 <= {src73[10:0], in_data73};
        src74 <= {src74[10:0], in_data74};
        src75 <= {src75[10:0], in_data75};
        src76 <= {src76[10:0], in_data76};
        src77 <= {src77[10:0], in_data77};
        src78 <= {src78[10:0], in_data78};
        src79 <= {src79[10:0], in_data79};
        src80 <= {src80[10:0], in_data80};
        src81 <= {src81[10:0], in_data81};
        src82 <= {src82[10:0], in_data82};
        src83 <= {src83[10:0], in_data83};
        src84 <= {src84[10:0], in_data84};
        src85 <= {src85[10:0], in_data85};
        src86 <= {src86[10:0], in_data86};
        src87 <= {src87[10:0], in_data87};
        src88 <= {src88[10:0], in_data88};
        src89 <= {src89[10:0], in_data89};
        src90 <= {src90[10:0], in_data90};
        src91 <= {src91[10:0], in_data91};
        src92 <= {src92[10:0], in_data92};
        src93 <= {src93[10:0], in_data93};
        src94 <= {src94[10:0], in_data94};
        src95 <= {src95[10:0], in_data95};
        src96 <= {src96[10:0], in_data96};
        src97 <= {src97[10:0], in_data97};
        src98 <= {src98[10:0], in_data98};
        src99 <= {src99[10:0], in_data99};
        src100 <= {src100[10:0], in_data100};
        src101 <= {src101[10:0], in_data101};
        src102 <= {src102[10:0], in_data102};
        src103 <= {src103[10:0], in_data103};
        src104 <= {src104[10:0], in_data104};
        src105 <= {src105[10:0], in_data105};
        src106 <= {src106[10:0], in_data106};
        src107 <= {src107[10:0], in_data107};
        src108 <= {src108[10:0], in_data108};
        src109 <= {src109[10:0], in_data109};
        src110 <= {src110[10:0], in_data110};
        src111 <= {src111[10:0], in_data111};
        src112 <= {src112[10:0], in_data112};
        src113 <= {src113[10:0], in_data113};
        src114 <= {src114[10:0], in_data114};
        src115 <= {src115[10:0], in_data115};
        src116 <= {src116[10:0], in_data116};
        src117 <= {src117[10:0], in_data117};
        src118 <= {src118[10:0], in_data118};
        src119 <= {src119[10:0], in_data119};
        src120 <= {src120[10:0], in_data120};
        src121 <= {src121[10:0], in_data121};
        src122 <= {src122[10:0], in_data122};
        src123 <= {src123[10:0], in_data123};
        src124 <= {src124[10:0], in_data124};
        src125 <= {src125[10:0], in_data125};
        src126 <= {src126[10:0], in_data126};
        src127 <= {src127[10:0], in_data127};
        src128 <= {src128[10:0], in_data128};
        src129 <= {src129[10:0], in_data129};
        src130 <= {src130[10:0], in_data130};
        src131 <= {src131[10:0], in_data131};
        src132 <= {src132[10:0], in_data132};
        src133 <= {src133[10:0], in_data133};
        src134 <= {src134[10:0], in_data134};
        src135 <= {src135[10:0], in_data135};
        src136 <= {src136[10:0], in_data136};
        src137 <= {src137[10:0], in_data137};
        src138 <= {src138[10:0], in_data138};
        src139 <= {src139[10:0], in_data139};
        src140 <= {src140[10:0], in_data140};
        src141 <= {src141[10:0], in_data141};
        src142 <= {src142[10:0], in_data142};
        src143 <= {src143[10:0], in_data143};
        src144 <= {src144[10:0], in_data144};
        src145 <= {src145[10:0], in_data145};
        src146 <= {src146[10:0], in_data146};
        src147 <= {src147[10:0], in_data147};
        src148 <= {src148[10:0], in_data148};
        src149 <= {src149[10:0], in_data149};
        src150 <= {src150[10:0], in_data150};
        src151 <= {src151[10:0], in_data151};
        src152 <= {src152[10:0], in_data152};
        src153 <= {src153[10:0], in_data153};
        src154 <= {src154[10:0], in_data154};
        src155 <= {src155[10:0], in_data155};
        src156 <= {src156[10:0], in_data156};
        src157 <= {src157[10:0], in_data157};
        src158 <= {src158[10:0], in_data158};
        src159 <= {src159[10:0], in_data159};
        src160 <= {src160[10:0], in_data160};
        src161 <= {src161[10:0], in_data161};
    end
endmodule

module compressor2_1_162_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    input [11:0]src32,
    input [11:0]src33,
    input [11:0]src34,
    input [11:0]src35,
    input [11:0]src36,
    input [11:0]src37,
    input [11:0]src38,
    input [11:0]src39,
    input [11:0]src40,
    input [11:0]src41,
    input [11:0]src42,
    input [11:0]src43,
    input [11:0]src44,
    input [11:0]src45,
    input [11:0]src46,
    input [11:0]src47,
    input [11:0]src48,
    input [11:0]src49,
    input [11:0]src50,
    input [11:0]src51,
    input [11:0]src52,
    input [11:0]src53,
    input [11:0]src54,
    input [11:0]src55,
    input [11:0]src56,
    input [11:0]src57,
    input [11:0]src58,
    input [11:0]src59,
    input [11:0]src60,
    input [11:0]src61,
    input [11:0]src62,
    input [11:0]src63,
    input [11:0]src64,
    input [11:0]src65,
    input [11:0]src66,
    input [11:0]src67,
    input [11:0]src68,
    input [11:0]src69,
    input [11:0]src70,
    input [11:0]src71,
    input [11:0]src72,
    input [11:0]src73,
    input [11:0]src74,
    input [11:0]src75,
    input [11:0]src76,
    input [11:0]src77,
    input [11:0]src78,
    input [11:0]src79,
    input [11:0]src80,
    input [11:0]src81,
    input [11:0]src82,
    input [11:0]src83,
    input [11:0]src84,
    input [11:0]src85,
    input [11:0]src86,
    input [11:0]src87,
    input [11:0]src88,
    input [11:0]src89,
    input [11:0]src90,
    input [11:0]src91,
    input [11:0]src92,
    input [11:0]src93,
    input [11:0]src94,
    input [11:0]src95,
    input [11:0]src96,
    input [11:0]src97,
    input [11:0]src98,
    input [11:0]src99,
    input [11:0]src100,
    input [11:0]src101,
    input [11:0]src102,
    input [11:0]src103,
    input [11:0]src104,
    input [11:0]src105,
    input [11:0]src106,
    input [11:0]src107,
    input [11:0]src108,
    input [11:0]src109,
    input [11:0]src110,
    input [11:0]src111,
    input [11:0]src112,
    input [11:0]src113,
    input [11:0]src114,
    input [11:0]src115,
    input [11:0]src116,
    input [11:0]src117,
    input [11:0]src118,
    input [11:0]src119,
    input [11:0]src120,
    input [11:0]src121,
    input [11:0]src122,
    input [11:0]src123,
    input [11:0]src124,
    input [11:0]src125,
    input [11:0]src126,
    input [11:0]src127,
    input [11:0]src128,
    input [11:0]src129,
    input [11:0]src130,
    input [11:0]src131,
    input [11:0]src132,
    input [11:0]src133,
    input [11:0]src134,
    input [11:0]src135,
    input [11:0]src136,
    input [11:0]src137,
    input [11:0]src138,
    input [11:0]src139,
    input [11:0]src140,
    input [11:0]src141,
    input [11:0]src142,
    input [11:0]src143,
    input [11:0]src144,
    input [11:0]src145,
    input [11:0]src146,
    input [11:0]src147,
    input [11:0]src148,
    input [11:0]src149,
    input [11:0]src150,
    input [11:0]src151,
    input [11:0]src152,
    input [11:0]src153,
    input [11:0]src154,
    input [11:0]src155,
    input [11:0]src156,
    input [11:0]src157,
    input [11:0]src158,
    input [11:0]src159,
    input [11:0]src160,
    input [11:0]src161,
    output [19:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [0:0] comp_out18;
    wire [19:0] out;
    compressor compressor_inst(
        .src0({src161[0], src160[0], src159[0], src158[0], src157[0], src156[0], src155[0], src154[0], src153[0], src152[0], src151[0], src150[0], src149[0], src148[0], src147[0], src146[0], src145[0], src144[0], src143[0], src142[0], src141[0], src140[0], src139[0], src138[0], src137[0], src136[0], src135[0], src134[0], src133[0], src132[0], src131[0], src130[0], src129[0], src128[0], src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src161[1], src160[1], src159[1], src158[1], src157[1], src156[1], src155[1], src154[1], src153[1], src152[1], src151[1], src150[1], src149[1], src148[1], src147[1], src146[1], src145[1], src144[1], src143[1], src142[1], src141[1], src140[1], src139[1], src138[1], src137[1], src136[1], src135[1], src134[1], src133[1], src132[1], src131[1], src130[1], src129[1], src128[1], src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src161[2], src160[2], src159[2], src158[2], src157[2], src156[2], src155[2], src154[2], src153[2], src152[2], src151[2], src150[2], src149[2], src148[2], src147[2], src146[2], src145[2], src144[2], src143[2], src142[2], src141[2], src140[2], src139[2], src138[2], src137[2], src136[2], src135[2], src134[2], src133[2], src132[2], src131[2], src130[2], src129[2], src128[2], src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src161[3], src160[3], src159[3], src158[3], src157[3], src156[3], src155[3], src154[3], src153[3], src152[3], src151[3], src150[3], src149[3], src148[3], src147[3], src146[3], src145[3], src144[3], src143[3], src142[3], src141[3], src140[3], src139[3], src138[3], src137[3], src136[3], src135[3], src134[3], src133[3], src132[3], src131[3], src130[3], src129[3], src128[3], src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src161[4], src160[4], src159[4], src158[4], src157[4], src156[4], src155[4], src154[4], src153[4], src152[4], src151[4], src150[4], src149[4], src148[4], src147[4], src146[4], src145[4], src144[4], src143[4], src142[4], src141[4], src140[4], src139[4], src138[4], src137[4], src136[4], src135[4], src134[4], src133[4], src132[4], src131[4], src130[4], src129[4], src128[4], src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src161[5], src160[5], src159[5], src158[5], src157[5], src156[5], src155[5], src154[5], src153[5], src152[5], src151[5], src150[5], src149[5], src148[5], src147[5], src146[5], src145[5], src144[5], src143[5], src142[5], src141[5], src140[5], src139[5], src138[5], src137[5], src136[5], src135[5], src134[5], src133[5], src132[5], src131[5], src130[5], src129[5], src128[5], src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src161[6], src160[6], src159[6], src158[6], src157[6], src156[6], src155[6], src154[6], src153[6], src152[6], src151[6], src150[6], src149[6], src148[6], src147[6], src146[6], src145[6], src144[6], src143[6], src142[6], src141[6], src140[6], src139[6], src138[6], src137[6], src136[6], src135[6], src134[6], src133[6], src132[6], src131[6], src130[6], src129[6], src128[6], src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src161[7], src160[7], src159[7], src158[7], src157[7], src156[7], src155[7], src154[7], src153[7], src152[7], src151[7], src150[7], src149[7], src148[7], src147[7], src146[7], src145[7], src144[7], src143[7], src142[7], src141[7], src140[7], src139[7], src138[7], src137[7], src136[7], src135[7], src134[7], src133[7], src132[7], src131[7], src130[7], src129[7], src128[7], src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src161[8], src160[8], src159[8], src158[8], src157[8], src156[8], src155[8], src154[8], src153[8], src152[8], src151[8], src150[8], src149[8], src148[8], src147[8], src146[8], src145[8], src144[8], src143[8], src142[8], src141[8], src140[8], src139[8], src138[8], src137[8], src136[8], src135[8], src134[8], src133[8], src132[8], src131[8], src130[8], src129[8], src128[8], src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src161[9], src160[9], src159[9], src158[9], src157[9], src156[9], src155[9], src154[9], src153[9], src152[9], src151[9], src150[9], src149[9], src148[9], src147[9], src146[9], src145[9], src144[9], src143[9], src142[9], src141[9], src140[9], src139[9], src138[9], src137[9], src136[9], src135[9], src134[9], src133[9], src132[9], src131[9], src130[9], src129[9], src128[9], src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src161[10], src160[10], src159[10], src158[10], src157[10], src156[10], src155[10], src154[10], src153[10], src152[10], src151[10], src150[10], src149[10], src148[10], src147[10], src146[10], src145[10], src144[10], src143[10], src142[10], src141[10], src140[10], src139[10], src138[10], src137[10], src136[10], src135[10], src134[10], src133[10], src132[10], src131[10], src130[10], src129[10], src128[10], src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src161[11], src160[11], src159[11], src158[11], src157[11], src156[11], src155[11], src154[11], src153[11], src152[11], src151[11], src150[11], src149[11], src148[11], src147[11], src146[11], src145[11], src144[11], src143[11], src142[11], src141[11], src140[11], src139[11], src138[11], src137[11], src136[11], src135[11], src134[11], src133[11], src132[11], src131[11], src130[11], src129[11], src128[11], src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    rowadder2_1_19 rowadder2_1inst(
        .src0({comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[19:0];
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [0:0] dst18);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [51:0] stage1_0;
   wire [47:0] stage1_1;
   wire [53:0] stage1_2;
   wire [77:0] stage1_3;
   wire [75:0] stage1_4;
   wire [75:0] stage1_5;
   wire [73:0] stage1_6;
   wire [48:0] stage1_7;
   wire [75:0] stage1_8;
   wire [80:0] stage1_9;
   wire [53:0] stage1_10;
   wire [53:0] stage1_11;
   wire [53:0] stage1_12;
   wire [26:0] stage1_13;
   wire [46:0] stage2_0;
   wire [33:0] stage2_1;
   wire [21:0] stage2_2;
   wire [21:0] stage2_3;
   wire [33:0] stage2_4;
   wire [24:0] stage2_5;
   wire [35:0] stage2_6;
   wire [32:0] stage2_7;
   wire [25:0] stage2_8;
   wire [23:0] stage2_9;
   wire [31:0] stage2_10;
   wire [35:0] stage2_11;
   wire [20:0] stage2_12;
   wire [29:0] stage2_13;
   wire [9:0] stage2_14;
   wire [1:0] stage2_15;
   wire [9:0] stage3_0;
   wire [13:0] stage3_1;
   wire [17:0] stage3_2;
   wire [9:0] stage3_3;
   wire [18:0] stage3_4;
   wire [9:0] stage3_5;
   wire [9:0] stage3_6;
   wire [11:0] stage3_7;
   wire [18:0] stage3_8;
   wire [10:0] stage3_9;
   wire [11:0] stage3_10;
   wire [12:0] stage3_11;
   wire [19:0] stage3_12;
   wire [7:0] stage3_13;
   wire [10:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [9:0] stage4_0;
   wire [8:0] stage4_1;
   wire [3:0] stage4_2;
   wire [7:0] stage4_3;
   wire [4:0] stage4_4;
   wire [8:0] stage4_5;
   wire [5:0] stage4_6;
   wire [8:0] stage4_7;
   wire [3:0] stage4_8;
   wire [5:0] stage4_9;
   wire [5:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [10:0] stage4_13;
   wire [8:0] stage4_14;
   wire [4:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;
   wire [5:0] stage5_0;
   wire [3:0] stage5_1;
   wire [1:0] stage5_2;
   wire [2:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [1:0] stage5_6;
   wire [2:0] stage5_7;
   wire [4:0] stage5_8;
   wire [1:0] stage5_9;
   wire [6:0] stage5_10;
   wire [4:0] stage5_11;
   wire [0:0] stage5_12;
   wire [6:0] stage5_13;
   wire [4:0] stage5_14;
   wire [1:0] stage5_15;
   wire [3:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [0:0] stage6_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc615_5 gpc10 (
      {stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_1[24]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc615_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[25]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc615_5 gpc12 (
      {stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[26]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc615_5 gpc13 (
      {stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[27]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc615_5 gpc14 (
      {stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[28]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc615_5 gpc15 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[29]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc615_5 gpc16 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[30]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc615_5 gpc17 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_1[31]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc615_5 gpc18 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[32]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc615_5 gpc19 (
      {stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_1[33]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc615_5 gpc20 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[34]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[35]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_1[36]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[37]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc615_5 gpc24 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[38]},
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc615_5 gpc25 (
      {stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_1[39]},
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc615_5 gpc26 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136]},
      {stage0_1[40]},
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46]},
      {stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21]},
      {stage1_5[0],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52]},
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27]},
      {stage1_5[1],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[2],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[3],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[4],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[5],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[6],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[7],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[8],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[9],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[10],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[11],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[12],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[13],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[14],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[15],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[16],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[17],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154]},
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage1_5[18],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160]},
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135]},
      {stage1_5[19],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[20],stage1_4[47],stage1_3[47],stage1_2[47]}
   );
   gpc606_5 gpc48 (
      {stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[21],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc606_5 gpc49 (
      {stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[22],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc606_5 gpc50 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[23],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc606_5 gpc51 (
      {stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[24],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage0_3[136]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[25],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage0_3[137]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[26],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[7],stage1_5[27],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[8],stage1_5[28],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[9],stage1_5[29],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[10],stage1_5[30],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[11],stage1_5[31],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[12],stage1_5[32],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[13],stage1_5[33],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[14],stage1_5[34],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[15],stage1_5[35],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[16],stage1_5[36],stage1_4[63]}
   );
   gpc615_5 gpc64 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106]},
      {stage0_5[0]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[17],stage1_5[37],stage1_4[64]}
   );
   gpc615_5 gpc65 (
      {stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_5[1]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[18],stage1_5[38],stage1_4[65]}
   );
   gpc615_5 gpc66 (
      {stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116]},
      {stage0_5[2]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[19],stage1_5[39],stage1_4[66]}
   );
   gpc615_5 gpc67 (
      {stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_5[3]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[20],stage1_5[40],stage1_4[67]}
   );
   gpc615_5 gpc68 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_5[4]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[21],stage1_5[41],stage1_4[68]}
   );
   gpc615_5 gpc69 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_5[5]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[22],stage1_5[42],stage1_4[69]}
   );
   gpc615_5 gpc70 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136]},
      {stage0_5[6]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[23],stage1_5[43],stage1_4[70]}
   );
   gpc615_5 gpc71 (
      {stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_5[7]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[24],stage1_5[44],stage1_4[71]}
   );
   gpc615_5 gpc72 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146]},
      {stage0_5[8]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[25],stage1_5[45],stage1_4[72]}
   );
   gpc615_5 gpc73 (
      {stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_5[9]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[26],stage1_5[46],stage1_4[73]}
   );
   gpc615_5 gpc74 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156]},
      {stage0_5[10]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[20],stage1_6[27],stage1_5[47],stage1_4[74]}
   );
   gpc615_5 gpc75 (
      {stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_5[11]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[21],stage1_6[28],stage1_5[48],stage1_4[75]}
   );
   gpc606_5 gpc76 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[22],stage1_7[22],stage1_6[29],stage1_5[49]}
   );
   gpc606_5 gpc77 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[23],stage1_7[23],stage1_6[30],stage1_5[50]}
   );
   gpc606_5 gpc78 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[24],stage1_7[24],stage1_6[31],stage1_5[51]}
   );
   gpc606_5 gpc79 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[25],stage1_7[25],stage1_6[32],stage1_5[52]}
   );
   gpc606_5 gpc80 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[26],stage1_7[26],stage1_6[33],stage1_5[53]}
   );
   gpc606_5 gpc81 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[27],stage1_7[27],stage1_6[34],stage1_5[54]}
   );
   gpc606_5 gpc82 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[28],stage1_7[28],stage1_6[35],stage1_5[55]}
   );
   gpc606_5 gpc83 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[29],stage1_7[29],stage1_6[36],stage1_5[56]}
   );
   gpc606_5 gpc84 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[30],stage1_7[30],stage1_6[37],stage1_5[57]}
   );
   gpc606_5 gpc85 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[31],stage1_7[31],stage1_6[38],stage1_5[58]}
   );
   gpc606_5 gpc86 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[32],stage1_7[32],stage1_6[39],stage1_5[59]}
   );
   gpc606_5 gpc87 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[33],stage1_7[33],stage1_6[40],stage1_5[60]}
   );
   gpc606_5 gpc88 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[34],stage1_7[34],stage1_6[41],stage1_5[61]}
   );
   gpc606_5 gpc89 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[35],stage1_7[35],stage1_6[42],stage1_5[62]}
   );
   gpc606_5 gpc90 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[36],stage1_7[36],stage1_6[43],stage1_5[63]}
   );
   gpc615_5 gpc91 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106]},
      {stage0_6[132]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[37],stage1_7[37],stage1_6[44],stage1_5[64]}
   );
   gpc615_5 gpc92 (
      {stage0_5[107], stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111]},
      {stage0_6[133]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[38],stage1_7[38],stage1_6[45],stage1_5[65]}
   );
   gpc615_5 gpc93 (
      {stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116]},
      {stage0_6[134]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[39],stage1_7[39],stage1_6[46],stage1_5[66]}
   );
   gpc615_5 gpc94 (
      {stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121]},
      {stage0_6[135]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[40],stage1_7[40],stage1_6[47],stage1_5[67]}
   );
   gpc615_5 gpc95 (
      {stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126]},
      {stage0_6[136]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[41],stage1_7[41],stage1_6[48],stage1_5[68]}
   );
   gpc615_5 gpc96 (
      {stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_6[137]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[42],stage1_7[42],stage1_6[49],stage1_5[69]}
   );
   gpc615_5 gpc97 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136]},
      {stage0_6[138]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[43],stage1_7[43],stage1_6[50],stage1_5[70]}
   );
   gpc615_5 gpc98 (
      {stage0_5[137], stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141]},
      {stage0_6[139]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[44],stage1_7[44],stage1_6[51],stage1_5[71]}
   );
   gpc615_5 gpc99 (
      {stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145], stage0_5[146]},
      {stage0_6[140]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[45],stage1_7[45],stage1_6[52],stage1_5[72]}
   );
   gpc615_5 gpc100 (
      {stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_6[141]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[46],stage1_7[46],stage1_6[53],stage1_5[73]}
   );
   gpc615_5 gpc101 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156]},
      {stage0_6[142]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[47],stage1_7[47],stage1_6[54],stage1_5[74]}
   );
   gpc615_5 gpc102 (
      {stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_6[143]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[48],stage1_7[48],stage1_6[55],stage1_5[75]}
   );
   gpc606_5 gpc103 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[27],stage1_8[49]}
   );
   gpc606_5 gpc104 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[1],stage1_9[28],stage1_8[50]}
   );
   gpc606_5 gpc105 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[2],stage1_9[29],stage1_8[51]}
   );
   gpc606_5 gpc106 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[3],stage1_9[30],stage1_8[52]}
   );
   gpc606_5 gpc107 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[4],stage1_9[31],stage1_8[53]}
   );
   gpc606_5 gpc108 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[5],stage1_9[32],stage1_8[54]}
   );
   gpc606_5 gpc109 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[6],stage1_9[33],stage1_8[55]}
   );
   gpc606_5 gpc110 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[7],stage1_9[34],stage1_8[56]}
   );
   gpc606_5 gpc111 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[8],stage1_9[35],stage1_8[57]}
   );
   gpc606_5 gpc112 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[9],stage1_9[36],stage1_8[58]}
   );
   gpc606_5 gpc113 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[10],stage1_9[37],stage1_8[59]}
   );
   gpc606_5 gpc114 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[11],stage1_9[38],stage1_8[60]}
   );
   gpc606_5 gpc115 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[12],stage1_9[39],stage1_8[61]}
   );
   gpc606_5 gpc116 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[13],stage1_9[40],stage1_8[62]}
   );
   gpc606_5 gpc117 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[14],stage1_9[41],stage1_8[63]}
   );
   gpc606_5 gpc118 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[15],stage1_9[42],stage1_8[64]}
   );
   gpc606_5 gpc119 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[16],stage1_9[43],stage1_8[65]}
   );
   gpc606_5 gpc120 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[17],stage1_9[44],stage1_8[66]}
   );
   gpc606_5 gpc121 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[18],stage1_9[45],stage1_8[67]}
   );
   gpc606_5 gpc122 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[19],stage1_9[46],stage1_8[68]}
   );
   gpc606_5 gpc123 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[20],stage1_9[47],stage1_8[69]}
   );
   gpc606_5 gpc124 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[21],stage1_10[21],stage1_9[48],stage1_8[70]}
   );
   gpc606_5 gpc125 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[22],stage1_10[22],stage1_9[49],stage1_8[71]}
   );
   gpc606_5 gpc126 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[23],stage1_10[23],stage1_9[50],stage1_8[72]}
   );
   gpc606_5 gpc127 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[24],stage1_10[24],stage1_9[51],stage1_8[73]}
   );
   gpc606_5 gpc128 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[25],stage1_10[25],stage1_9[52],stage1_8[74]}
   );
   gpc606_5 gpc129 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[26],stage1_10[26],stage1_9[53],stage1_8[75]}
   );
   gpc606_5 gpc130 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[27],stage1_11[27],stage1_10[27],stage1_9[54]}
   );
   gpc606_5 gpc131 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[28],stage1_11[28],stage1_10[28],stage1_9[55]}
   );
   gpc606_5 gpc132 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[29],stage1_11[29],stage1_10[29],stage1_9[56]}
   );
   gpc606_5 gpc133 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[30],stage1_11[30],stage1_10[30],stage1_9[57]}
   );
   gpc606_5 gpc134 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[31],stage1_11[31],stage1_10[31],stage1_9[58]}
   );
   gpc606_5 gpc135 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[32],stage1_11[32],stage1_10[32],stage1_9[59]}
   );
   gpc606_5 gpc136 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[33],stage1_11[33],stage1_10[33],stage1_9[60]}
   );
   gpc606_5 gpc137 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[34],stage1_11[34],stage1_10[34],stage1_9[61]}
   );
   gpc606_5 gpc138 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[35],stage1_11[35],stage1_10[35],stage1_9[62]}
   );
   gpc606_5 gpc139 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[36],stage1_11[36],stage1_10[36],stage1_9[63]}
   );
   gpc606_5 gpc140 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[37],stage1_11[37],stage1_10[37],stage1_9[64]}
   );
   gpc606_5 gpc141 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[38],stage1_11[38],stage1_10[38],stage1_9[65]}
   );
   gpc606_5 gpc142 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[39],stage1_11[39],stage1_10[39],stage1_9[66]}
   );
   gpc606_5 gpc143 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[40],stage1_11[40],stage1_10[40],stage1_9[67]}
   );
   gpc606_5 gpc144 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[41],stage1_11[41],stage1_10[41],stage1_9[68]}
   );
   gpc606_5 gpc145 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[42],stage1_11[42],stage1_10[42],stage1_9[69]}
   );
   gpc606_5 gpc146 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[43],stage1_11[43],stage1_10[43],stage1_9[70]}
   );
   gpc606_5 gpc147 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[44],stage1_11[44],stage1_10[44],stage1_9[71]}
   );
   gpc606_5 gpc148 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[45],stage1_11[45],stage1_10[45],stage1_9[72]}
   );
   gpc606_5 gpc149 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[46],stage1_11[46],stage1_10[46],stage1_9[73]}
   );
   gpc606_5 gpc150 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[47],stage1_11[47],stage1_10[47],stage1_9[74]}
   );
   gpc606_5 gpc151 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[48],stage1_11[48],stage1_10[48],stage1_9[75]}
   );
   gpc606_5 gpc152 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[49],stage1_11[49],stage1_10[49],stage1_9[76]}
   );
   gpc606_5 gpc153 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[50],stage1_11[50],stage1_10[50],stage1_9[77]}
   );
   gpc606_5 gpc154 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[51],stage1_11[51],stage1_10[51],stage1_9[78]}
   );
   gpc606_5 gpc155 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[52],stage1_11[52],stage1_10[52],stage1_9[79]}
   );
   gpc606_5 gpc156 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[53],stage1_11[53],stage1_10[53],stage1_9[80]}
   );
   gpc1_1 gpc157 (
      {stage0_0[137]},
      {stage1_0[27]}
   );
   gpc1_1 gpc158 (
      {stage0_0[138]},
      {stage1_0[28]}
   );
   gpc1_1 gpc159 (
      {stage0_0[139]},
      {stage1_0[29]}
   );
   gpc1_1 gpc160 (
      {stage0_0[140]},
      {stage1_0[30]}
   );
   gpc1_1 gpc161 (
      {stage0_0[141]},
      {stage1_0[31]}
   );
   gpc1_1 gpc162 (
      {stage0_0[142]},
      {stage1_0[32]}
   );
   gpc1_1 gpc163 (
      {stage0_0[143]},
      {stage1_0[33]}
   );
   gpc1_1 gpc164 (
      {stage0_0[144]},
      {stage1_0[34]}
   );
   gpc1_1 gpc165 (
      {stage0_0[145]},
      {stage1_0[35]}
   );
   gpc1_1 gpc166 (
      {stage0_0[146]},
      {stage1_0[36]}
   );
   gpc1_1 gpc167 (
      {stage0_0[147]},
      {stage1_0[37]}
   );
   gpc1_1 gpc168 (
      {stage0_0[148]},
      {stage1_0[38]}
   );
   gpc1_1 gpc169 (
      {stage0_0[149]},
      {stage1_0[39]}
   );
   gpc1_1 gpc170 (
      {stage0_0[150]},
      {stage1_0[40]}
   );
   gpc1_1 gpc171 (
      {stage0_0[151]},
      {stage1_0[41]}
   );
   gpc1_1 gpc172 (
      {stage0_0[152]},
      {stage1_0[42]}
   );
   gpc1_1 gpc173 (
      {stage0_0[153]},
      {stage1_0[43]}
   );
   gpc1_1 gpc174 (
      {stage0_0[154]},
      {stage1_0[44]}
   );
   gpc1_1 gpc175 (
      {stage0_0[155]},
      {stage1_0[45]}
   );
   gpc1_1 gpc176 (
      {stage0_0[156]},
      {stage1_0[46]}
   );
   gpc1_1 gpc177 (
      {stage0_0[157]},
      {stage1_0[47]}
   );
   gpc1_1 gpc178 (
      {stage0_0[158]},
      {stage1_0[48]}
   );
   gpc1_1 gpc179 (
      {stage0_0[159]},
      {stage1_0[49]}
   );
   gpc1_1 gpc180 (
      {stage0_0[160]},
      {stage1_0[50]}
   );
   gpc1_1 gpc181 (
      {stage0_0[161]},
      {stage1_0[51]}
   );
   gpc1_1 gpc182 (
      {stage0_1[161]},
      {stage1_1[47]}
   );
   gpc1_1 gpc183 (
      {stage0_3[138]},
      {stage1_3[54]}
   );
   gpc1_1 gpc184 (
      {stage0_3[139]},
      {stage1_3[55]}
   );
   gpc1_1 gpc185 (
      {stage0_3[140]},
      {stage1_3[56]}
   );
   gpc1_1 gpc186 (
      {stage0_3[141]},
      {stage1_3[57]}
   );
   gpc1_1 gpc187 (
      {stage0_3[142]},
      {stage1_3[58]}
   );
   gpc1_1 gpc188 (
      {stage0_3[143]},
      {stage1_3[59]}
   );
   gpc1_1 gpc189 (
      {stage0_3[144]},
      {stage1_3[60]}
   );
   gpc1_1 gpc190 (
      {stage0_3[145]},
      {stage1_3[61]}
   );
   gpc1_1 gpc191 (
      {stage0_3[146]},
      {stage1_3[62]}
   );
   gpc1_1 gpc192 (
      {stage0_3[147]},
      {stage1_3[63]}
   );
   gpc1_1 gpc193 (
      {stage0_3[148]},
      {stage1_3[64]}
   );
   gpc1_1 gpc194 (
      {stage0_3[149]},
      {stage1_3[65]}
   );
   gpc1_1 gpc195 (
      {stage0_3[150]},
      {stage1_3[66]}
   );
   gpc1_1 gpc196 (
      {stage0_3[151]},
      {stage1_3[67]}
   );
   gpc1_1 gpc197 (
      {stage0_3[152]},
      {stage1_3[68]}
   );
   gpc1_1 gpc198 (
      {stage0_3[153]},
      {stage1_3[69]}
   );
   gpc1_1 gpc199 (
      {stage0_3[154]},
      {stage1_3[70]}
   );
   gpc1_1 gpc200 (
      {stage0_3[155]},
      {stage1_3[71]}
   );
   gpc1_1 gpc201 (
      {stage0_3[156]},
      {stage1_3[72]}
   );
   gpc1_1 gpc202 (
      {stage0_3[157]},
      {stage1_3[73]}
   );
   gpc1_1 gpc203 (
      {stage0_3[158]},
      {stage1_3[74]}
   );
   gpc1_1 gpc204 (
      {stage0_3[159]},
      {stage1_3[75]}
   );
   gpc1_1 gpc205 (
      {stage0_3[160]},
      {stage1_3[76]}
   );
   gpc1_1 gpc206 (
      {stage0_3[161]},
      {stage1_3[77]}
   );
   gpc1_1 gpc207 (
      {stage0_6[144]},
      {stage1_6[56]}
   );
   gpc1_1 gpc208 (
      {stage0_6[145]},
      {stage1_6[57]}
   );
   gpc1_1 gpc209 (
      {stage0_6[146]},
      {stage1_6[58]}
   );
   gpc1_1 gpc210 (
      {stage0_6[147]},
      {stage1_6[59]}
   );
   gpc1_1 gpc211 (
      {stage0_6[148]},
      {stage1_6[60]}
   );
   gpc1_1 gpc212 (
      {stage0_6[149]},
      {stage1_6[61]}
   );
   gpc1_1 gpc213 (
      {stage0_6[150]},
      {stage1_6[62]}
   );
   gpc1_1 gpc214 (
      {stage0_6[151]},
      {stage1_6[63]}
   );
   gpc1_1 gpc215 (
      {stage0_6[152]},
      {stage1_6[64]}
   );
   gpc1_1 gpc216 (
      {stage0_6[153]},
      {stage1_6[65]}
   );
   gpc1_1 gpc217 (
      {stage0_6[154]},
      {stage1_6[66]}
   );
   gpc1_1 gpc218 (
      {stage0_6[155]},
      {stage1_6[67]}
   );
   gpc1_1 gpc219 (
      {stage0_6[156]},
      {stage1_6[68]}
   );
   gpc1_1 gpc220 (
      {stage0_6[157]},
      {stage1_6[69]}
   );
   gpc1_1 gpc221 (
      {stage0_6[158]},
      {stage1_6[70]}
   );
   gpc1_1 gpc222 (
      {stage0_6[159]},
      {stage1_6[71]}
   );
   gpc1_1 gpc223 (
      {stage0_6[160]},
      {stage1_6[72]}
   );
   gpc1_1 gpc224 (
      {stage0_6[161]},
      {stage1_6[73]}
   );
   gpc606_5 gpc225 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc226 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc227 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc228 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc229 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc230 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc606_5 gpc231 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[5],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc232 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[6],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc233 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[7],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc606_5 gpc234 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[8],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc235 (
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage1_4[36]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[6],stage2_5[9],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc236 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[37]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[7],stage2_5[10],stage2_4[11],stage2_3[11]}
   );
   gpc615_5 gpc237 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage1_4[38]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[8],stage2_5[11],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc238 (
      {stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage1_4[39]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[9],stage2_5[12],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc239 (
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage1_4[40]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[10],stage2_5[13],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc240 (
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage1_4[41]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[11],stage2_5[14],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc241 (
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52]},
      {stage1_4[42]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[12],stage2_5[15],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc242 (
      {stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage1_4[43]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[13],stage2_5[16],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc243 (
      {stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62]},
      {stage1_4[44]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[14],stage2_5[17],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc244 (
      {stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage1_4[45]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[15],stage2_5[18],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc245 (
      {stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72]},
      {stage1_4[46]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[16],stage2_5[19],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc246 (
      {stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage1_4[47]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[17],stage2_5[20],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc247 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52]},
      {stage1_5[72]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[12],stage2_6[18],stage2_5[21],stage2_4[22]}
   );
   gpc615_5 gpc248 (
      {stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_5[73]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[13],stage2_6[19],stage2_5[22],stage2_4[23]}
   );
   gpc615_5 gpc249 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_5[74]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[14],stage2_6[20],stage2_5[23],stage2_4[24]}
   );
   gpc615_5 gpc250 (
      {stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67]},
      {stage1_5[75]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[15],stage2_6[21],stage2_5[24],stage2_4[25]}
   );
   gpc615_5 gpc251 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28]},
      {stage1_7[0]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[4],stage2_7[16],stage2_6[22]}
   );
   gpc615_5 gpc252 (
      {stage1_6[29], stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33]},
      {stage1_7[1]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[5],stage2_7[17],stage2_6[23]}
   );
   gpc615_5 gpc253 (
      {stage1_6[34], stage1_6[35], stage1_6[36], stage1_6[37], stage1_6[38]},
      {stage1_7[2]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[6],stage2_7[18],stage2_6[24]}
   );
   gpc615_5 gpc254 (
      {stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42], stage1_6[43]},
      {stage1_7[3]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[3],stage2_8[7],stage2_7[19],stage2_6[25]}
   );
   gpc615_5 gpc255 (
      {stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage1_7[4]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[4],stage2_8[8],stage2_7[20],stage2_6[26]}
   );
   gpc615_5 gpc256 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_7[5]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[5],stage2_8[9],stage2_7[21],stage2_6[27]}
   );
   gpc615_5 gpc257 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58]},
      {stage1_7[6]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[6],stage2_8[10],stage2_7[22],stage2_6[28]}
   );
   gpc615_5 gpc258 (
      {stage1_6[59], stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63]},
      {stage1_7[7]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[7],stage2_8[11],stage2_7[23],stage2_6[29]}
   );
   gpc615_5 gpc259 (
      {stage1_6[64], stage1_6[65], stage1_6[66], stage1_6[67], stage1_6[68]},
      {stage1_7[8]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[8],stage2_8[12],stage2_7[24],stage2_6[30]}
   );
   gpc615_5 gpc260 (
      {stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage1_8[54]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[9],stage2_9[9],stage2_8[13],stage2_7[25]}
   );
   gpc615_5 gpc261 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage1_8[55]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[10],stage2_9[10],stage2_8[14],stage2_7[26]}
   );
   gpc615_5 gpc262 (
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_8[56]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[11],stage2_9[11],stage2_8[15],stage2_7[27]}
   );
   gpc615_5 gpc263 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[57]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[12],stage2_9[12],stage2_8[16],stage2_7[28]}
   );
   gpc615_5 gpc264 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[58]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[13],stage2_9[13],stage2_8[17],stage2_7[29]}
   );
   gpc615_5 gpc265 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[59]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[14],stage2_9[14],stage2_8[18],stage2_7[30]}
   );
   gpc615_5 gpc266 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[60]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[15],stage2_9[15],stage2_8[19],stage2_7[31]}
   );
   gpc615_5 gpc267 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[61]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[16],stage2_9[16],stage2_8[20],stage2_7[32]}
   );
   gpc2135_5 gpc268 (
      {stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_9[48], stage1_9[49], stage1_9[50]},
      {stage1_10[0]},
      {stage1_11[0], stage1_11[1]},
      {stage2_12[0],stage2_11[8],stage2_10[17],stage2_9[17],stage2_8[21]}
   );
   gpc606_5 gpc269 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[9],stage2_10[18],stage2_9[18],stage2_8[22]}
   );
   gpc606_5 gpc270 (
      {stage1_9[51], stage1_9[52], stage1_9[53], stage1_9[54], stage1_9[55], stage1_9[56]},
      {stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7]},
      {stage2_13[0],stage2_12[2],stage2_11[10],stage2_10[19],stage2_9[19]}
   );
   gpc606_5 gpc271 (
      {stage1_9[57], stage1_9[58], stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62]},
      {stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage2_13[1],stage2_12[3],stage2_11[11],stage2_10[20],stage2_9[20]}
   );
   gpc606_5 gpc272 (
      {stage1_9[63], stage1_9[64], stage1_9[65], stage1_9[66], stage1_9[67], stage1_9[68]},
      {stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage2_13[2],stage2_12[4],stage2_11[12],stage2_10[21],stage2_9[21]}
   );
   gpc606_5 gpc273 (
      {stage1_9[69], stage1_9[70], stage1_9[71], stage1_9[72], stage1_9[73], stage1_9[74]},
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25]},
      {stage2_13[3],stage2_12[5],stage2_11[13],stage2_10[22],stage2_9[22]}
   );
   gpc606_5 gpc274 (
      {stage1_9[75], stage1_9[76], stage1_9[77], stage1_9[78], stage1_9[79], stage1_9[80]},
      {stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30], stage1_11[31]},
      {stage2_13[4],stage2_12[6],stage2_11[14],stage2_10[23],stage2_9[23]}
   );
   gpc606_5 gpc275 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[5],stage2_12[7],stage2_11[15],stage2_10[24]}
   );
   gpc606_5 gpc276 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[6],stage2_12[8],stage2_11[16],stage2_10[25]}
   );
   gpc606_5 gpc277 (
      {stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[7],stage2_12[9],stage2_11[17],stage2_10[26]}
   );
   gpc606_5 gpc278 (
      {stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[8],stage2_12[10],stage2_11[18],stage2_10[27]}
   );
   gpc606_5 gpc279 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[9],stage2_12[11],stage2_11[19],stage2_10[28]}
   );
   gpc606_5 gpc280 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[10],stage2_12[12],stage2_11[20],stage2_10[29]}
   );
   gpc606_5 gpc281 (
      {stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[11],stage2_12[13],stage2_11[21],stage2_10[30]}
   );
   gpc615_5 gpc282 (
      {stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_11[32]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[12],stage2_12[14],stage2_11[22],stage2_10[31]}
   );
   gpc615_5 gpc283 (
      {stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37]},
      {stage1_12[48]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[8],stage2_13[13],stage2_12[15],stage2_11[23]}
   );
   gpc615_5 gpc284 (
      {stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_12[49]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[9],stage2_13[14],stage2_12[16],stage2_11[24]}
   );
   gpc1_1 gpc285 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc286 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc287 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc288 (
      {stage1_0[9]},
      {stage2_0[4]}
   );
   gpc1_1 gpc289 (
      {stage1_0[10]},
      {stage2_0[5]}
   );
   gpc1_1 gpc290 (
      {stage1_0[11]},
      {stage2_0[6]}
   );
   gpc1_1 gpc291 (
      {stage1_0[12]},
      {stage2_0[7]}
   );
   gpc1_1 gpc292 (
      {stage1_0[13]},
      {stage2_0[8]}
   );
   gpc1_1 gpc293 (
      {stage1_0[14]},
      {stage2_0[9]}
   );
   gpc1_1 gpc294 (
      {stage1_0[15]},
      {stage2_0[10]}
   );
   gpc1_1 gpc295 (
      {stage1_0[16]},
      {stage2_0[11]}
   );
   gpc1_1 gpc296 (
      {stage1_0[17]},
      {stage2_0[12]}
   );
   gpc1_1 gpc297 (
      {stage1_0[18]},
      {stage2_0[13]}
   );
   gpc1_1 gpc298 (
      {stage1_0[19]},
      {stage2_0[14]}
   );
   gpc1_1 gpc299 (
      {stage1_0[20]},
      {stage2_0[15]}
   );
   gpc1_1 gpc300 (
      {stage1_0[21]},
      {stage2_0[16]}
   );
   gpc1_1 gpc301 (
      {stage1_0[22]},
      {stage2_0[17]}
   );
   gpc1_1 gpc302 (
      {stage1_0[23]},
      {stage2_0[18]}
   );
   gpc1_1 gpc303 (
      {stage1_0[24]},
      {stage2_0[19]}
   );
   gpc1_1 gpc304 (
      {stage1_0[25]},
      {stage2_0[20]}
   );
   gpc1_1 gpc305 (
      {stage1_0[26]},
      {stage2_0[21]}
   );
   gpc1_1 gpc306 (
      {stage1_0[27]},
      {stage2_0[22]}
   );
   gpc1_1 gpc307 (
      {stage1_0[28]},
      {stage2_0[23]}
   );
   gpc1_1 gpc308 (
      {stage1_0[29]},
      {stage2_0[24]}
   );
   gpc1_1 gpc309 (
      {stage1_0[30]},
      {stage2_0[25]}
   );
   gpc1_1 gpc310 (
      {stage1_0[31]},
      {stage2_0[26]}
   );
   gpc1_1 gpc311 (
      {stage1_0[32]},
      {stage2_0[27]}
   );
   gpc1_1 gpc312 (
      {stage1_0[33]},
      {stage2_0[28]}
   );
   gpc1_1 gpc313 (
      {stage1_0[34]},
      {stage2_0[29]}
   );
   gpc1_1 gpc314 (
      {stage1_0[35]},
      {stage2_0[30]}
   );
   gpc1_1 gpc315 (
      {stage1_0[36]},
      {stage2_0[31]}
   );
   gpc1_1 gpc316 (
      {stage1_0[37]},
      {stage2_0[32]}
   );
   gpc1_1 gpc317 (
      {stage1_0[38]},
      {stage2_0[33]}
   );
   gpc1_1 gpc318 (
      {stage1_0[39]},
      {stage2_0[34]}
   );
   gpc1_1 gpc319 (
      {stage1_0[40]},
      {stage2_0[35]}
   );
   gpc1_1 gpc320 (
      {stage1_0[41]},
      {stage2_0[36]}
   );
   gpc1_1 gpc321 (
      {stage1_0[42]},
      {stage2_0[37]}
   );
   gpc1_1 gpc322 (
      {stage1_0[43]},
      {stage2_0[38]}
   );
   gpc1_1 gpc323 (
      {stage1_0[44]},
      {stage2_0[39]}
   );
   gpc1_1 gpc324 (
      {stage1_0[45]},
      {stage2_0[40]}
   );
   gpc1_1 gpc325 (
      {stage1_0[46]},
      {stage2_0[41]}
   );
   gpc1_1 gpc326 (
      {stage1_0[47]},
      {stage2_0[42]}
   );
   gpc1_1 gpc327 (
      {stage1_0[48]},
      {stage2_0[43]}
   );
   gpc1_1 gpc328 (
      {stage1_0[49]},
      {stage2_0[44]}
   );
   gpc1_1 gpc329 (
      {stage1_0[50]},
      {stage2_0[45]}
   );
   gpc1_1 gpc330 (
      {stage1_0[51]},
      {stage2_0[46]}
   );
   gpc1_1 gpc331 (
      {stage1_1[18]},
      {stage2_1[4]}
   );
   gpc1_1 gpc332 (
      {stage1_1[19]},
      {stage2_1[5]}
   );
   gpc1_1 gpc333 (
      {stage1_1[20]},
      {stage2_1[6]}
   );
   gpc1_1 gpc334 (
      {stage1_1[21]},
      {stage2_1[7]}
   );
   gpc1_1 gpc335 (
      {stage1_1[22]},
      {stage2_1[8]}
   );
   gpc1_1 gpc336 (
      {stage1_1[23]},
      {stage2_1[9]}
   );
   gpc1_1 gpc337 (
      {stage1_1[24]},
      {stage2_1[10]}
   );
   gpc1_1 gpc338 (
      {stage1_1[25]},
      {stage2_1[11]}
   );
   gpc1_1 gpc339 (
      {stage1_1[26]},
      {stage2_1[12]}
   );
   gpc1_1 gpc340 (
      {stage1_1[27]},
      {stage2_1[13]}
   );
   gpc1_1 gpc341 (
      {stage1_1[28]},
      {stage2_1[14]}
   );
   gpc1_1 gpc342 (
      {stage1_1[29]},
      {stage2_1[15]}
   );
   gpc1_1 gpc343 (
      {stage1_1[30]},
      {stage2_1[16]}
   );
   gpc1_1 gpc344 (
      {stage1_1[31]},
      {stage2_1[17]}
   );
   gpc1_1 gpc345 (
      {stage1_1[32]},
      {stage2_1[18]}
   );
   gpc1_1 gpc346 (
      {stage1_1[33]},
      {stage2_1[19]}
   );
   gpc1_1 gpc347 (
      {stage1_1[34]},
      {stage2_1[20]}
   );
   gpc1_1 gpc348 (
      {stage1_1[35]},
      {stage2_1[21]}
   );
   gpc1_1 gpc349 (
      {stage1_1[36]},
      {stage2_1[22]}
   );
   gpc1_1 gpc350 (
      {stage1_1[37]},
      {stage2_1[23]}
   );
   gpc1_1 gpc351 (
      {stage1_1[38]},
      {stage2_1[24]}
   );
   gpc1_1 gpc352 (
      {stage1_1[39]},
      {stage2_1[25]}
   );
   gpc1_1 gpc353 (
      {stage1_1[40]},
      {stage2_1[26]}
   );
   gpc1_1 gpc354 (
      {stage1_1[41]},
      {stage2_1[27]}
   );
   gpc1_1 gpc355 (
      {stage1_1[42]},
      {stage2_1[28]}
   );
   gpc1_1 gpc356 (
      {stage1_1[43]},
      {stage2_1[29]}
   );
   gpc1_1 gpc357 (
      {stage1_1[44]},
      {stage2_1[30]}
   );
   gpc1_1 gpc358 (
      {stage1_1[45]},
      {stage2_1[31]}
   );
   gpc1_1 gpc359 (
      {stage1_1[46]},
      {stage2_1[32]}
   );
   gpc1_1 gpc360 (
      {stage1_1[47]},
      {stage2_1[33]}
   );
   gpc1_1 gpc361 (
      {stage1_2[42]},
      {stage2_2[10]}
   );
   gpc1_1 gpc362 (
      {stage1_2[43]},
      {stage2_2[11]}
   );
   gpc1_1 gpc363 (
      {stage1_2[44]},
      {stage2_2[12]}
   );
   gpc1_1 gpc364 (
      {stage1_2[45]},
      {stage2_2[13]}
   );
   gpc1_1 gpc365 (
      {stage1_2[46]},
      {stage2_2[14]}
   );
   gpc1_1 gpc366 (
      {stage1_2[47]},
      {stage2_2[15]}
   );
   gpc1_1 gpc367 (
      {stage1_2[48]},
      {stage2_2[16]}
   );
   gpc1_1 gpc368 (
      {stage1_2[49]},
      {stage2_2[17]}
   );
   gpc1_1 gpc369 (
      {stage1_2[50]},
      {stage2_2[18]}
   );
   gpc1_1 gpc370 (
      {stage1_2[51]},
      {stage2_2[19]}
   );
   gpc1_1 gpc371 (
      {stage1_2[52]},
      {stage2_2[20]}
   );
   gpc1_1 gpc372 (
      {stage1_2[53]},
      {stage2_2[21]}
   );
   gpc1_1 gpc373 (
      {stage1_4[68]},
      {stage2_4[26]}
   );
   gpc1_1 gpc374 (
      {stage1_4[69]},
      {stage2_4[27]}
   );
   gpc1_1 gpc375 (
      {stage1_4[70]},
      {stage2_4[28]}
   );
   gpc1_1 gpc376 (
      {stage1_4[71]},
      {stage2_4[29]}
   );
   gpc1_1 gpc377 (
      {stage1_4[72]},
      {stage2_4[30]}
   );
   gpc1_1 gpc378 (
      {stage1_4[73]},
      {stage2_4[31]}
   );
   gpc1_1 gpc379 (
      {stage1_4[74]},
      {stage2_4[32]}
   );
   gpc1_1 gpc380 (
      {stage1_4[75]},
      {stage2_4[33]}
   );
   gpc1_1 gpc381 (
      {stage1_6[69]},
      {stage2_6[31]}
   );
   gpc1_1 gpc382 (
      {stage1_6[70]},
      {stage2_6[32]}
   );
   gpc1_1 gpc383 (
      {stage1_6[71]},
      {stage2_6[33]}
   );
   gpc1_1 gpc384 (
      {stage1_6[72]},
      {stage2_6[34]}
   );
   gpc1_1 gpc385 (
      {stage1_6[73]},
      {stage2_6[35]}
   );
   gpc1_1 gpc386 (
      {stage1_8[73]},
      {stage2_8[23]}
   );
   gpc1_1 gpc387 (
      {stage1_8[74]},
      {stage2_8[24]}
   );
   gpc1_1 gpc388 (
      {stage1_8[75]},
      {stage2_8[25]}
   );
   gpc1_1 gpc389 (
      {stage1_11[43]},
      {stage2_11[25]}
   );
   gpc1_1 gpc390 (
      {stage1_11[44]},
      {stage2_11[26]}
   );
   gpc1_1 gpc391 (
      {stage1_11[45]},
      {stage2_11[27]}
   );
   gpc1_1 gpc392 (
      {stage1_11[46]},
      {stage2_11[28]}
   );
   gpc1_1 gpc393 (
      {stage1_11[47]},
      {stage2_11[29]}
   );
   gpc1_1 gpc394 (
      {stage1_11[48]},
      {stage2_11[30]}
   );
   gpc1_1 gpc395 (
      {stage1_11[49]},
      {stage2_11[31]}
   );
   gpc1_1 gpc396 (
      {stage1_11[50]},
      {stage2_11[32]}
   );
   gpc1_1 gpc397 (
      {stage1_11[51]},
      {stage2_11[33]}
   );
   gpc1_1 gpc398 (
      {stage1_11[52]},
      {stage2_11[34]}
   );
   gpc1_1 gpc399 (
      {stage1_11[53]},
      {stage2_11[35]}
   );
   gpc1_1 gpc400 (
      {stage1_12[50]},
      {stage2_12[17]}
   );
   gpc1_1 gpc401 (
      {stage1_12[51]},
      {stage2_12[18]}
   );
   gpc1_1 gpc402 (
      {stage1_12[52]},
      {stage2_12[19]}
   );
   gpc1_1 gpc403 (
      {stage1_12[53]},
      {stage2_12[20]}
   );
   gpc1_1 gpc404 (
      {stage1_13[12]},
      {stage2_13[15]}
   );
   gpc1_1 gpc405 (
      {stage1_13[13]},
      {stage2_13[16]}
   );
   gpc1_1 gpc406 (
      {stage1_13[14]},
      {stage2_13[17]}
   );
   gpc1_1 gpc407 (
      {stage1_13[15]},
      {stage2_13[18]}
   );
   gpc1_1 gpc408 (
      {stage1_13[16]},
      {stage2_13[19]}
   );
   gpc1_1 gpc409 (
      {stage1_13[17]},
      {stage2_13[20]}
   );
   gpc1_1 gpc410 (
      {stage1_13[18]},
      {stage2_13[21]}
   );
   gpc1_1 gpc411 (
      {stage1_13[19]},
      {stage2_13[22]}
   );
   gpc1_1 gpc412 (
      {stage1_13[20]},
      {stage2_13[23]}
   );
   gpc1_1 gpc413 (
      {stage1_13[21]},
      {stage2_13[24]}
   );
   gpc1_1 gpc414 (
      {stage1_13[22]},
      {stage2_13[25]}
   );
   gpc1_1 gpc415 (
      {stage1_13[23]},
      {stage2_13[26]}
   );
   gpc1_1 gpc416 (
      {stage1_13[24]},
      {stage2_13[27]}
   );
   gpc1_1 gpc417 (
      {stage1_13[25]},
      {stage2_13[28]}
   );
   gpc1_1 gpc418 (
      {stage1_13[26]},
      {stage2_13[29]}
   );
   gpc2135_5 gpc419 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc2135_5 gpc420 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[1]},
      {stage2_3[2], stage2_3[3]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc2135_5 gpc421 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_2[2]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc2135_5 gpc422 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19]},
      {stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[3]},
      {stage2_3[6], stage2_3[7]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc2135_5 gpc423 (
      {stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24]},
      {stage2_1[12], stage2_1[13], stage2_1[14]},
      {stage2_2[4]},
      {stage2_3[8], stage2_3[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc2135_5 gpc424 (
      {stage2_0[25], stage2_0[26], stage2_0[27], stage2_0[28], stage2_0[29]},
      {stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[5]},
      {stage2_3[10], stage2_3[11]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc2135_5 gpc425 (
      {stage2_0[30], stage2_0[31], stage2_0[32], stage2_0[33], stage2_0[34]},
      {stage2_1[18], stage2_1[19], stage2_1[20]},
      {stage2_2[6]},
      {stage2_3[12], stage2_3[13]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc2135_5 gpc426 (
      {stage2_0[35], stage2_0[36], stage2_0[37], stage2_0[38], stage2_0[39]},
      {stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[7]},
      {stage2_3[14], stage2_3[15]},
      {stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7],stage3_0[7]}
   );
   gpc606_5 gpc427 (
      {stage2_0[40], stage2_0[41], stage2_0[42], stage2_0[43], stage2_0[44], stage2_0[45]},
      {stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13]},
      {stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8],stage3_0[8]}
   );
   gpc606_5 gpc428 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21]},
      {stage3_5[0],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc2135_5 gpc429 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage2_7[0], stage2_7[1]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[10]}
   );
   gpc606_5 gpc430 (
      {stage2_4[5], stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[1],stage3_7[1],stage3_6[1],stage3_5[2],stage3_4[11]}
   );
   gpc615_5 gpc431 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[3]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[2],stage3_7[2],stage3_6[2],stage3_5[3],stage3_4[12]}
   );
   gpc615_5 gpc432 (
      {stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_5[4]},
      {stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18]},
      {stage3_8[3],stage3_7[3],stage3_6[3],stage3_5[4],stage3_4[13]}
   );
   gpc615_5 gpc433 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[5]},
      {stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24]},
      {stage3_8[4],stage3_7[4],stage3_6[4],stage3_5[5],stage3_4[14]}
   );
   gpc615_5 gpc434 (
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30]},
      {stage2_5[6]},
      {stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage3_8[5],stage3_7[5],stage3_6[5],stage3_5[6],stage3_4[15]}
   );
   gpc606_5 gpc435 (
      {stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6], stage2_7[7]},
      {stage3_9[0],stage3_8[6],stage3_7[6],stage3_6[6],stage3_5[7]}
   );
   gpc606_5 gpc436 (
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18]},
      {stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage3_9[1],stage3_8[7],stage3_7[7],stage3_6[7],stage3_5[8]}
   );
   gpc606_5 gpc437 (
      {stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24]},
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19]},
      {stage3_9[2],stage3_8[8],stage3_7[8],stage3_6[8],stage3_5[9]}
   );
   gpc2135_5 gpc438 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[3],stage3_8[9],stage3_7[9],stage3_6[9]}
   );
   gpc615_5 gpc439 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[1]},
      {stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7]},
      {stage3_11[0],stage3_10[1],stage3_9[4],stage3_8[10],stage3_7[10]}
   );
   gpc615_5 gpc440 (
      {stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[2]},
      {stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13]},
      {stage3_11[1],stage3_10[2],stage3_9[5],stage3_8[11],stage3_7[11]}
   );
   gpc615_5 gpc441 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_9[14]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[3],stage3_9[6],stage3_8[12]}
   );
   gpc615_5 gpc442 (
      {stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12]},
      {stage2_9[15]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[4],stage3_9[7],stage3_8[13]}
   );
   gpc615_5 gpc443 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage2_9[16]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[4],stage3_10[5],stage3_9[8],stage3_8[14]}
   );
   gpc615_5 gpc444 (
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22]},
      {stage2_9[17]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[5],stage3_10[6],stage3_9[9],stage3_8[15]}
   );
   gpc606_5 gpc445 (
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[4],stage3_11[6],stage3_10[7],stage3_9[10]}
   );
   gpc615_5 gpc446 (
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28]},
      {stage2_11[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[5],stage3_11[7],stage3_10[8]}
   );
   gpc606_5 gpc447 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[6],stage3_11[8]}
   );
   gpc606_5 gpc448 (
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[2],stage3_13[3],stage3_12[7],stage3_11[9]}
   );
   gpc606_5 gpc449 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[3],stage3_13[4],stage3_12[8],stage3_11[10]}
   );
   gpc606_5 gpc450 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[4],stage3_13[5],stage3_12[9],stage3_11[11]}
   );
   gpc615_5 gpc451 (
      {stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage2_12[6]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[5],stage3_13[6],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc452 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[6],stage3_13[7],stage3_12[11]}
   );
   gpc1_1 gpc453 (
      {stage2_0[46]},
      {stage3_0[9]}
   );
   gpc1_1 gpc454 (
      {stage2_1[30]},
      {stage3_1[10]}
   );
   gpc1_1 gpc455 (
      {stage2_1[31]},
      {stage3_1[11]}
   );
   gpc1_1 gpc456 (
      {stage2_1[32]},
      {stage3_1[12]}
   );
   gpc1_1 gpc457 (
      {stage2_1[33]},
      {stage3_1[13]}
   );
   gpc1_1 gpc458 (
      {stage2_2[14]},
      {stage3_2[10]}
   );
   gpc1_1 gpc459 (
      {stage2_2[15]},
      {stage3_2[11]}
   );
   gpc1_1 gpc460 (
      {stage2_2[16]},
      {stage3_2[12]}
   );
   gpc1_1 gpc461 (
      {stage2_2[17]},
      {stage3_2[13]}
   );
   gpc1_1 gpc462 (
      {stage2_2[18]},
      {stage3_2[14]}
   );
   gpc1_1 gpc463 (
      {stage2_2[19]},
      {stage3_2[15]}
   );
   gpc1_1 gpc464 (
      {stage2_2[20]},
      {stage3_2[16]}
   );
   gpc1_1 gpc465 (
      {stage2_2[21]},
      {stage3_2[17]}
   );
   gpc1_1 gpc466 (
      {stage2_4[31]},
      {stage3_4[16]}
   );
   gpc1_1 gpc467 (
      {stage2_4[32]},
      {stage3_4[17]}
   );
   gpc1_1 gpc468 (
      {stage2_4[33]},
      {stage3_4[18]}
   );
   gpc1_1 gpc469 (
      {stage2_8[23]},
      {stage3_8[16]}
   );
   gpc1_1 gpc470 (
      {stage2_8[24]},
      {stage3_8[17]}
   );
   gpc1_1 gpc471 (
      {stage2_8[25]},
      {stage3_8[18]}
   );
   gpc1_1 gpc472 (
      {stage2_10[29]},
      {stage3_10[9]}
   );
   gpc1_1 gpc473 (
      {stage2_10[30]},
      {stage3_10[10]}
   );
   gpc1_1 gpc474 (
      {stage2_10[31]},
      {stage3_10[11]}
   );
   gpc1_1 gpc475 (
      {stage2_12[13]},
      {stage3_12[12]}
   );
   gpc1_1 gpc476 (
      {stage2_12[14]},
      {stage3_12[13]}
   );
   gpc1_1 gpc477 (
      {stage2_12[15]},
      {stage3_12[14]}
   );
   gpc1_1 gpc478 (
      {stage2_12[16]},
      {stage3_12[15]}
   );
   gpc1_1 gpc479 (
      {stage2_12[17]},
      {stage3_12[16]}
   );
   gpc1_1 gpc480 (
      {stage2_12[18]},
      {stage3_12[17]}
   );
   gpc1_1 gpc481 (
      {stage2_12[19]},
      {stage3_12[18]}
   );
   gpc1_1 gpc482 (
      {stage2_12[20]},
      {stage3_12[19]}
   );
   gpc1_1 gpc483 (
      {stage2_14[6]},
      {stage3_14[7]}
   );
   gpc1_1 gpc484 (
      {stage2_14[7]},
      {stage3_14[8]}
   );
   gpc1_1 gpc485 (
      {stage2_14[8]},
      {stage3_14[9]}
   );
   gpc1_1 gpc486 (
      {stage2_14[9]},
      {stage3_14[10]}
   );
   gpc1_1 gpc487 (
      {stage2_15[0]},
      {stage3_15[6]}
   );
   gpc1_1 gpc488 (
      {stage2_15[1]},
      {stage3_15[7]}
   );
   gpc606_5 gpc489 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc490 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc606_5 gpc491 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc492 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc1406_5 gpc493 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[3],stage4_5[4]}
   );
   gpc615_5 gpc494 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[4]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6]},
      {stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1],stage4_6[4]}
   );
   gpc615_5 gpc495 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[5]},
      {stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12]},
      {stage4_10[1],stage4_9[2],stage4_8[2],stage4_7[2],stage4_6[5]}
   );
   gpc606_5 gpc496 (
      {stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17], stage3_8[18]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[2],stage4_9[3],stage4_8[3]}
   );
   gpc606_5 gpc497 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[1],stage4_10[3],stage4_9[4]}
   );
   gpc615_5 gpc498 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[6]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[2],stage4_11[2],stage4_10[4],stage4_9[5]}
   );
   gpc615_5 gpc499 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[3],stage4_11[3],stage4_10[5]}
   );
   gpc207_4 gpc500 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[1],stage4_13[3],stage4_12[4]}
   );
   gpc207_4 gpc501 (
      {stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18], stage3_12[19]},
      {stage3_14[2], stage3_14[3]},
      {stage4_15[1],stage4_14[2],stage4_13[4],stage4_12[5]}
   );
   gpc623_5 gpc502 (
      {stage3_13[0], stage3_13[1], stage3_13[2]},
      {stage3_14[4], stage3_14[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[2],stage4_14[3],stage4_13[5]}
   );
   gpc1_1 gpc503 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc504 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc505 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc506 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc507 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc508 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc509 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc510 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc511 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc512 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc513 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc514 (
      {stage3_1[7]},
      {stage4_1[2]}
   );
   gpc1_1 gpc515 (
      {stage3_1[8]},
      {stage4_1[3]}
   );
   gpc1_1 gpc516 (
      {stage3_1[9]},
      {stage4_1[4]}
   );
   gpc1_1 gpc517 (
      {stage3_1[10]},
      {stage4_1[5]}
   );
   gpc1_1 gpc518 (
      {stage3_1[11]},
      {stage4_1[6]}
   );
   gpc1_1 gpc519 (
      {stage3_1[12]},
      {stage4_1[7]}
   );
   gpc1_1 gpc520 (
      {stage3_1[13]},
      {stage4_1[8]}
   );
   gpc1_1 gpc521 (
      {stage3_3[6]},
      {stage4_3[4]}
   );
   gpc1_1 gpc522 (
      {stage3_3[7]},
      {stage4_3[5]}
   );
   gpc1_1 gpc523 (
      {stage3_3[8]},
      {stage4_3[6]}
   );
   gpc1_1 gpc524 (
      {stage3_3[9]},
      {stage4_3[7]}
   );
   gpc1_1 gpc525 (
      {stage3_4[18]},
      {stage4_4[4]}
   );
   gpc1_1 gpc526 (
      {stage3_5[6]},
      {stage4_5[5]}
   );
   gpc1_1 gpc527 (
      {stage3_5[7]},
      {stage4_5[6]}
   );
   gpc1_1 gpc528 (
      {stage3_5[8]},
      {stage4_5[7]}
   );
   gpc1_1 gpc529 (
      {stage3_5[9]},
      {stage4_5[8]}
   );
   gpc1_1 gpc530 (
      {stage3_7[6]},
      {stage4_7[3]}
   );
   gpc1_1 gpc531 (
      {stage3_7[7]},
      {stage4_7[4]}
   );
   gpc1_1 gpc532 (
      {stage3_7[8]},
      {stage4_7[5]}
   );
   gpc1_1 gpc533 (
      {stage3_7[9]},
      {stage4_7[6]}
   );
   gpc1_1 gpc534 (
      {stage3_7[10]},
      {stage4_7[7]}
   );
   gpc1_1 gpc535 (
      {stage3_7[11]},
      {stage4_7[8]}
   );
   gpc1_1 gpc536 (
      {stage3_13[3]},
      {stage4_13[6]}
   );
   gpc1_1 gpc537 (
      {stage3_13[4]},
      {stage4_13[7]}
   );
   gpc1_1 gpc538 (
      {stage3_13[5]},
      {stage4_13[8]}
   );
   gpc1_1 gpc539 (
      {stage3_13[6]},
      {stage4_13[9]}
   );
   gpc1_1 gpc540 (
      {stage3_13[7]},
      {stage4_13[10]}
   );
   gpc1_1 gpc541 (
      {stage3_14[6]},
      {stage4_14[4]}
   );
   gpc1_1 gpc542 (
      {stage3_14[7]},
      {stage4_14[5]}
   );
   gpc1_1 gpc543 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc544 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc545 (
      {stage3_14[10]},
      {stage4_14[8]}
   );
   gpc1_1 gpc546 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc547 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc1_1 gpc548 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
   gpc1325_5 gpc549 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1]},
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc615_5 gpc550 (
      {stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_2[3]},
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc623_5 gpc551 (
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0], stage4_5[1]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[2]}
   );
   gpc1406_5 gpc552 (
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[2]}
   );
   gpc615_5 gpc553 (
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7], stage4_7[8]},
      {stage4_8[1]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2]}
   );
   gpc606_5 gpc554 (
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[0]}
   );
   gpc606_5 gpc555 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], 1'b0},
      {stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1],stage5_13[1]}
   );
   gpc1_1 gpc556 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc557 (
      {stage4_0[6]},
      {stage5_0[2]}
   );
   gpc1_1 gpc558 (
      {stage4_0[7]},
      {stage5_0[3]}
   );
   gpc1_1 gpc559 (
      {stage4_0[8]},
      {stage5_0[4]}
   );
   gpc1_1 gpc560 (
      {stage4_0[9]},
      {stage5_0[5]}
   );
   gpc1_1 gpc561 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc562 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc563 (
      {stage4_3[7]},
      {stage5_3[2]}
   );
   gpc1_1 gpc564 (
      {stage4_4[3]},
      {stage5_4[3]}
   );
   gpc1_1 gpc565 (
      {stage4_4[4]},
      {stage5_4[4]}
   );
   gpc1_1 gpc566 (
      {stage4_5[8]},
      {stage5_5[3]}
   );
   gpc1_1 gpc567 (
      {stage4_8[2]},
      {stage5_8[3]}
   );
   gpc1_1 gpc568 (
      {stage4_8[3]},
      {stage5_8[4]}
   );
   gpc1_1 gpc569 (
      {stage4_10[0]},
      {stage5_10[1]}
   );
   gpc1_1 gpc570 (
      {stage4_10[1]},
      {stage5_10[2]}
   );
   gpc1_1 gpc571 (
      {stage4_10[2]},
      {stage5_10[3]}
   );
   gpc1_1 gpc572 (
      {stage4_10[3]},
      {stage5_10[4]}
   );
   gpc1_1 gpc573 (
      {stage4_10[4]},
      {stage5_10[5]}
   );
   gpc1_1 gpc574 (
      {stage4_10[5]},
      {stage5_10[6]}
   );
   gpc1_1 gpc575 (
      {stage4_11[0]},
      {stage5_11[1]}
   );
   gpc1_1 gpc576 (
      {stage4_11[1]},
      {stage5_11[2]}
   );
   gpc1_1 gpc577 (
      {stage4_11[2]},
      {stage5_11[3]}
   );
   gpc1_1 gpc578 (
      {stage4_11[3]},
      {stage5_11[4]}
   );
   gpc1_1 gpc579 (
      {stage4_13[6]},
      {stage5_13[2]}
   );
   gpc1_1 gpc580 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc581 (
      {stage4_13[8]},
      {stage5_13[4]}
   );
   gpc1_1 gpc582 (
      {stage4_13[9]},
      {stage5_13[5]}
   );
   gpc1_1 gpc583 (
      {stage4_13[10]},
      {stage5_13[6]}
   );
   gpc1_1 gpc584 (
      {stage4_14[6]},
      {stage5_14[2]}
   );
   gpc1_1 gpc585 (
      {stage4_14[7]},
      {stage5_14[3]}
   );
   gpc1_1 gpc586 (
      {stage4_14[8]},
      {stage5_14[4]}
   );
   gpc1_1 gpc587 (
      {stage4_16[0]},
      {stage5_16[2]}
   );
   gpc1_1 gpc588 (
      {stage4_16[1]},
      {stage5_16[3]}
   );
   gpc1_1 gpc589 (
      {stage4_17[0]},
      {stage5_17[1]}
   );
   gpc2135_5 gpc590 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0]},
      {stage5_3[0], stage5_3[1]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc2135_5 gpc591 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4]},
      {stage5_5[0], stage5_5[1], stage5_5[2]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[1]}
   );
   gpc615_5 gpc592 (
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4]},
      {stage5_9[0]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc615_5 gpc593 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1325_5 gpc594 (
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1]}
   );
   gpc1_1 gpc595 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc596 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc597 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc598 (
      {stage5_3[2]},
      {stage6_3[1]}
   );
   gpc1_1 gpc599 (
      {stage5_5[3]},
      {stage6_5[1]}
   );
   gpc1_1 gpc600 (
      {stage5_6[1]},
      {stage6_6[1]}
   );
   gpc1_1 gpc601 (
      {stage5_7[2]},
      {stage6_7[1]}
   );
   gpc1_1 gpc602 (
      {stage5_9[1]},
      {stage6_9[1]}
   );
   gpc1_1 gpc603 (
      {stage5_10[6]},
      {stage6_10[1]}
   );
   gpc1_1 gpc604 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc605 (
      {stage5_16[3]},
      {stage6_16[1]}
   );
   gpc1_1 gpc606 (
      {stage5_17[1]},
      {stage6_17[1]}
   );
endmodule
module rowadder2_1_19(input [18:0] src0, input [18:0] src1, output [19:0] dst0);
    wire [18:0] gene;
    wire [18:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[18:16]}),
        .S({1'h0, prop[18:16]})
    );
    assign dst0 = {carryout[18], out[18:0]};
endmodule


module comp2_1test_162_12_162_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [11:0] src64;
    reg [11:0] src65;
    reg [11:0] src66;
    reg [11:0] src67;
    reg [11:0] src68;
    reg [11:0] src69;
    reg [11:0] src70;
    reg [11:0] src71;
    reg [11:0] src72;
    reg [11:0] src73;
    reg [11:0] src74;
    reg [11:0] src75;
    reg [11:0] src76;
    reg [11:0] src77;
    reg [11:0] src78;
    reg [11:0] src79;
    reg [11:0] src80;
    reg [11:0] src81;
    reg [11:0] src82;
    reg [11:0] src83;
    reg [11:0] src84;
    reg [11:0] src85;
    reg [11:0] src86;
    reg [11:0] src87;
    reg [11:0] src88;
    reg [11:0] src89;
    reg [11:0] src90;
    reg [11:0] src91;
    reg [11:0] src92;
    reg [11:0] src93;
    reg [11:0] src94;
    reg [11:0] src95;
    reg [11:0] src96;
    reg [11:0] src97;
    reg [11:0] src98;
    reg [11:0] src99;
    reg [11:0] src100;
    reg [11:0] src101;
    reg [11:0] src102;
    reg [11:0] src103;
    reg [11:0] src104;
    reg [11:0] src105;
    reg [11:0] src106;
    reg [11:0] src107;
    reg [11:0] src108;
    reg [11:0] src109;
    reg [11:0] src110;
    reg [11:0] src111;
    reg [11:0] src112;
    reg [11:0] src113;
    reg [11:0] src114;
    reg [11:0] src115;
    reg [11:0] src116;
    reg [11:0] src117;
    reg [11:0] src118;
    reg [11:0] src119;
    reg [11:0] src120;
    reg [11:0] src121;
    reg [11:0] src122;
    reg [11:0] src123;
    reg [11:0] src124;
    reg [11:0] src125;
    reg [11:0] src126;
    reg [11:0] src127;
    reg [11:0] src128;
    reg [11:0] src129;
    reg [11:0] src130;
    reg [11:0] src131;
    reg [11:0] src132;
    reg [11:0] src133;
    reg [11:0] src134;
    reg [11:0] src135;
    reg [11:0] src136;
    reg [11:0] src137;
    reg [11:0] src138;
    reg [11:0] src139;
    reg [11:0] src140;
    reg [11:0] src141;
    reg [11:0] src142;
    reg [11:0] src143;
    reg [11:0] src144;
    reg [11:0] src145;
    reg [11:0] src146;
    reg [11:0] src147;
    reg [11:0] src148;
    reg [11:0] src149;
    reg [11:0] src150;
    reg [11:0] src151;
    reg [11:0] src152;
    reg [11:0] src153;
    reg [11:0] src154;
    reg [11:0] src155;
    reg [11:0] src156;
    reg [11:0] src157;
    reg [11:0] src158;
    reg [11:0] src159;
    reg [11:0] src160;
    reg [11:0] src161;
    reg [19:0] exp;
    wire [19:0] dst;
    assign test = dst == exp;
    compressor2_1_162_12 compressor2_1_162_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .src128(src128),
        .src129(src129),
        .src130(src130),
        .src131(src131),
        .src132(src132),
        .src133(src133),
        .src134(src134),
        .src135(src135),
        .src136(src136),
        .src137(src137),
        .src138(src138),
        .src139(src139),
        .src140(src140),
        .src141(src141),
        .src142(src142),
        .src143(src143),
        .src144(src144),
        .src145(src145),
        .src146(src146),
        .src147(src147),
        .src148(src148),
        .src149(src149),
        .src150(src150),
        .src151(src151),
        .src152(src152),
        .src153(src153),
        .src154(src154),
        .src155(src155),
        .src156(src156),
        .src157(src157),
        .src158(src158),
        .src159(src159),
        .src160(src160),
        .src161(src161),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, src128, src129, src130, src131, src132, src133, src134, src135, src136, src137, src138, src139, src140, src141, src142, src143, src144, src145, src146, src147, src148, src149, src150, src151, src152, src153, src154, src155, src156, src157, src158, src159, src160, src161, dst, exp, test);
        src0 <= 12'hf3;
        src1 <= 12'h124;
        src2 <= 12'hf9a;
        src3 <= 12'h11e;
        src4 <= 12'hd16;
        src5 <= 12'h45a;
        src6 <= 12'hca9;
        src7 <= 12'h21d;
        src8 <= 12'h644;
        src9 <= 12'h1b9;
        src10 <= 12'hcff;
        src11 <= 12'ha0;
        src12 <= 12'h127;
        src13 <= 12'h4ba;
        src14 <= 12'hefa;
        src15 <= 12'h142;
        src16 <= 12'h492;
        src17 <= 12'h12a;
        src18 <= 12'h254;
        src19 <= 12'heaf;
        src20 <= 12'h70f;
        src21 <= 12'h83d;
        src22 <= 12'h7f9;
        src23 <= 12'ha21;
        src24 <= 12'he99;
        src25 <= 12'h78;
        src26 <= 12'hfa1;
        src27 <= 12'h2ce;
        src28 <= 12'h79f;
        src29 <= 12'haa7;
        src30 <= 12'ha8c;
        src31 <= 12'hb71;
        src32 <= 12'h27;
        src33 <= 12'h8d6;
        src34 <= 12'h6df;
        src35 <= 12'hcb6;
        src36 <= 12'h305;
        src37 <= 12'ha78;
        src38 <= 12'h2cf;
        src39 <= 12'hcb6;
        src40 <= 12'h4b9;
        src41 <= 12'h844;
        src42 <= 12'hef4;
        src43 <= 12'h26c;
        src44 <= 12'he82;
        src45 <= 12'h27e;
        src46 <= 12'h7e3;
        src47 <= 12'h4c3;
        src48 <= 12'hfa8;
        src49 <= 12'h985;
        src50 <= 12'hfa;
        src51 <= 12'h2e9;
        src52 <= 12'h972;
        src53 <= 12'h12d;
        src54 <= 12'hef0;
        src55 <= 12'h1a6;
        src56 <= 12'hdba;
        src57 <= 12'h456;
        src58 <= 12'h2e7;
        src59 <= 12'h534;
        src60 <= 12'h4b3;
        src61 <= 12'h278;
        src62 <= 12'ha2f;
        src63 <= 12'hcf3;
        src64 <= 12'hd68;
        src65 <= 12'h8d7;
        src66 <= 12'hc87;
        src67 <= 12'h750;
        src68 <= 12'hb65;
        src69 <= 12'hdcb;
        src70 <= 12'h407;
        src71 <= 12'h36a;
        src72 <= 12'h40b;
        src73 <= 12'ha0c;
        src74 <= 12'h3c4;
        src75 <= 12'h380;
        src76 <= 12'hb40;
        src77 <= 12'hcb2;
        src78 <= 12'h27;
        src79 <= 12'h39c;
        src80 <= 12'h455;
        src81 <= 12'h85f;
        src82 <= 12'h6c3;
        src83 <= 12'h6e2;
        src84 <= 12'h6ca;
        src85 <= 12'hb0a;
        src86 <= 12'hfb5;
        src87 <= 12'hde0;
        src88 <= 12'he02;
        src89 <= 12'he17;
        src90 <= 12'h7e8;
        src91 <= 12'h85f;
        src92 <= 12'h660;
        src93 <= 12'h3e3;
        src94 <= 12'h312;
        src95 <= 12'hadb;
        src96 <= 12'h49a;
        src97 <= 12'ha2;
        src98 <= 12'hab0;
        src99 <= 12'h548;
        src100 <= 12'h616;
        src101 <= 12'h3f2;
        src102 <= 12'h6d6;
        src103 <= 12'h167;
        src104 <= 12'had5;
        src105 <= 12'h83f;
        src106 <= 12'h60f;
        src107 <= 12'hdf6;
        src108 <= 12'h925;
        src109 <= 12'h9d4;
        src110 <= 12'hfff;
        src111 <= 12'h717;
        src112 <= 12'hff7;
        src113 <= 12'hf73;
        src114 <= 12'he91;
        src115 <= 12'hc55;
        src116 <= 12'hb40;
        src117 <= 12'he78;
        src118 <= 12'h251;
        src119 <= 12'hcab;
        src120 <= 12'h1b2;
        src121 <= 12'h6e1;
        src122 <= 12'hff7;
        src123 <= 12'ha7d;
        src124 <= 12'h5c6;
        src125 <= 12'h92e;
        src126 <= 12'hed6;
        src127 <= 12'hba;
        src128 <= 12'hfa8;
        src129 <= 12'he50;
        src130 <= 12'hc0;
        src131 <= 12'h51b;
        src132 <= 12'h658;
        src133 <= 12'h9b5;
        src134 <= 12'h604;
        src135 <= 12'haea;
        src136 <= 12'h975;
        src137 <= 12'hedb;
        src138 <= 12'hf19;
        src139 <= 12'h19;
        src140 <= 12'h560;
        src141 <= 12'hea9;
        src142 <= 12'he04;
        src143 <= 12'h37f;
        src144 <= 12'h395;
        src145 <= 12'h1de;
        src146 <= 12'ha5b;
        src147 <= 12'hb78;
        src148 <= 12'h1e1;
        src149 <= 12'h5;
        src150 <= 12'hf39;
        src151 <= 12'heb2;
        src152 <= 12'h94e;
        src153 <= 12'ha52;
        src154 <= 12'hafa;
        src155 <= 12'h5;
        src156 <= 12'h5f0;
        src157 <= 12'h6e3;
        src158 <= 12'h87c;
        src159 <= 12'hcb5;
        src160 <= 12'hb4b;
        src161 <= 12'h321;
        exp <= 20'h50a45;
        #1
        src0 <= 12'h676;
        src1 <= 12'h937;
        src2 <= 12'hfb;
        src3 <= 12'h734;
        src4 <= 12'hd85;
        src5 <= 12'hedd;
        src6 <= 12'h6fa;
        src7 <= 12'hb23;
        src8 <= 12'h8a8;
        src9 <= 12'h538;
        src10 <= 12'h72e;
        src11 <= 12'h4fc;
        src12 <= 12'hea0;
        src13 <= 12'h90;
        src14 <= 12'hb4d;
        src15 <= 12'h430;
        src16 <= 12'hdb1;
        src17 <= 12'h15;
        src18 <= 12'he9f;
        src19 <= 12'h91a;
        src20 <= 12'hef1;
        src21 <= 12'hf4a;
        src22 <= 12'hdd3;
        src23 <= 12'h261;
        src24 <= 12'hc30;
        src25 <= 12'h24c;
        src26 <= 12'hfb8;
        src27 <= 12'h9f;
        src28 <= 12'hb5a;
        src29 <= 12'h467;
        src30 <= 12'hd2b;
        src31 <= 12'h2dc;
        src32 <= 12'hf53;
        src33 <= 12'hbaa;
        src34 <= 12'h1b5;
        src35 <= 12'hab9;
        src36 <= 12'h355;
        src37 <= 12'haae;
        src38 <= 12'hb44;
        src39 <= 12'ha45;
        src40 <= 12'h5c8;
        src41 <= 12'h734;
        src42 <= 12'h465;
        src43 <= 12'hb53;
        src44 <= 12'h4a7;
        src45 <= 12'haa3;
        src46 <= 12'h3c9;
        src47 <= 12'h1a4;
        src48 <= 12'h161;
        src49 <= 12'hdde;
        src50 <= 12'h5a3;
        src51 <= 12'h8b8;
        src52 <= 12'h7cc;
        src53 <= 12'h8fa;
        src54 <= 12'ha0f;
        src55 <= 12'h5bd;
        src56 <= 12'he2d;
        src57 <= 12'h4f2;
        src58 <= 12'hb18;
        src59 <= 12'hedf;
        src60 <= 12'hfd0;
        src61 <= 12'he8b;
        src62 <= 12'h871;
        src63 <= 12'he8f;
        src64 <= 12'h2a5;
        src65 <= 12'h551;
        src66 <= 12'h66;
        src67 <= 12'h289;
        src68 <= 12'hf4;
        src69 <= 12'h264;
        src70 <= 12'hba4;
        src71 <= 12'h3ff;
        src72 <= 12'hb3c;
        src73 <= 12'h1d0;
        src74 <= 12'h193;
        src75 <= 12'h2ad;
        src76 <= 12'h5a;
        src77 <= 12'h572;
        src78 <= 12'h124;
        src79 <= 12'hcff;
        src80 <= 12'h39a;
        src81 <= 12'hdaa;
        src82 <= 12'hb0c;
        src83 <= 12'h673;
        src84 <= 12'hd88;
        src85 <= 12'h92c;
        src86 <= 12'hb13;
        src87 <= 12'hed2;
        src88 <= 12'h183;
        src89 <= 12'h314;
        src90 <= 12'h450;
        src91 <= 12'h74c;
        src92 <= 12'h4bb;
        src93 <= 12'hbaa;
        src94 <= 12'h73c;
        src95 <= 12'h260;
        src96 <= 12'h1b2;
        src97 <= 12'h3df;
        src98 <= 12'h4b2;
        src99 <= 12'habc;
        src100 <= 12'h8ce;
        src101 <= 12'ha3d;
        src102 <= 12'h860;
        src103 <= 12'h19e;
        src104 <= 12'h93f;
        src105 <= 12'ha6f;
        src106 <= 12'h982;
        src107 <= 12'h68d;
        src108 <= 12'he3;
        src109 <= 12'h533;
        src110 <= 12'h9d9;
        src111 <= 12'h2e8;
        src112 <= 12'he52;
        src113 <= 12'hc8b;
        src114 <= 12'h240;
        src115 <= 12'h2e7;
        src116 <= 12'h17f;
        src117 <= 12'h14e;
        src118 <= 12'had2;
        src119 <= 12'h72b;
        src120 <= 12'h73;
        src121 <= 12'hd75;
        src122 <= 12'h9fc;
        src123 <= 12'haf4;
        src124 <= 12'h913;
        src125 <= 12'h5f4;
        src126 <= 12'hbe0;
        src127 <= 12'hc91;
        src128 <= 12'ha12;
        src129 <= 12'h3c6;
        src130 <= 12'h652;
        src131 <= 12'h2ec;
        src132 <= 12'h75b;
        src133 <= 12'he72;
        src134 <= 12'hb72;
        src135 <= 12'h3a1;
        src136 <= 12'hbab;
        src137 <= 12'h571;
        src138 <= 12'hb21;
        src139 <= 12'hfc1;
        src140 <= 12'hdde;
        src141 <= 12'h349;
        src142 <= 12'he81;
        src143 <= 12'h3f;
        src144 <= 12'he8b;
        src145 <= 12'h313;
        src146 <= 12'hdcd;
        src147 <= 12'hfc9;
        src148 <= 12'h664;
        src149 <= 12'h9fa;
        src150 <= 12'hf9c;
        src151 <= 12'ha1;
        src152 <= 12'hdec;
        src153 <= 12'h7ff;
        src154 <= 12'h978;
        src155 <= 12'h6de;
        src156 <= 12'hb64;
        src157 <= 12'hf46;
        src158 <= 12'hf8;
        src159 <= 12'hc13;
        src160 <= 12'h3da;
        src161 <= 12'h90c;
        exp <= 20'h50985;
        #1
        src0 <= 12'h695;
        src1 <= 12'hd4e;
        src2 <= 12'h73e;
        src3 <= 12'ha53;
        src4 <= 12'h596;
        src5 <= 12'h226;
        src6 <= 12'h962;
        src7 <= 12'h8c4;
        src8 <= 12'h773;
        src9 <= 12'hd24;
        src10 <= 12'h25d;
        src11 <= 12'h3aa;
        src12 <= 12'hb26;
        src13 <= 12'h1ac;
        src14 <= 12'h3d;
        src15 <= 12'h923;
        src16 <= 12'hc59;
        src17 <= 12'he97;
        src18 <= 12'hd01;
        src19 <= 12'he72;
        src20 <= 12'hdc8;
        src21 <= 12'h8bf;
        src22 <= 12'h159;
        src23 <= 12'h4b5;
        src24 <= 12'h94;
        src25 <= 12'hcca;
        src26 <= 12'hc29;
        src27 <= 12'hfcb;
        src28 <= 12'he58;
        src29 <= 12'ha67;
        src30 <= 12'h492;
        src31 <= 12'h421;
        src32 <= 12'h34;
        src33 <= 12'h293;
        src34 <= 12'hf01;
        src35 <= 12'he0;
        src36 <= 12'hdc4;
        src37 <= 12'ha13;
        src38 <= 12'h8cc;
        src39 <= 12'h523;
        src40 <= 12'h22a;
        src41 <= 12'h1b4;
        src42 <= 12'h64d;
        src43 <= 12'he67;
        src44 <= 12'h574;
        src45 <= 12'h74d;
        src46 <= 12'h954;
        src47 <= 12'hf5a;
        src48 <= 12'h259;
        src49 <= 12'h1de;
        src50 <= 12'h62d;
        src51 <= 12'hb63;
        src52 <= 12'ha05;
        src53 <= 12'h73c;
        src54 <= 12'ha5c;
        src55 <= 12'h5f9;
        src56 <= 12'h326;
        src57 <= 12'he21;
        src58 <= 12'h6da;
        src59 <= 12'hae;
        src60 <= 12'h966;
        src61 <= 12'h222;
        src62 <= 12'h19c;
        src63 <= 12'hae0;
        src64 <= 12'h566;
        src65 <= 12'hee0;
        src66 <= 12'h6aa;
        src67 <= 12'hb27;
        src68 <= 12'had9;
        src69 <= 12'hfec;
        src70 <= 12'h4e0;
        src71 <= 12'hf58;
        src72 <= 12'h36c;
        src73 <= 12'h706;
        src74 <= 12'hfde;
        src75 <= 12'hd62;
        src76 <= 12'he4;
        src77 <= 12'hcb6;
        src78 <= 12'h995;
        src79 <= 12'hea2;
        src80 <= 12'h3da;
        src81 <= 12'h6c8;
        src82 <= 12'h6aa;
        src83 <= 12'h1a7;
        src84 <= 12'h3e6;
        src85 <= 12'h79;
        src86 <= 12'hc2e;
        src87 <= 12'h36b;
        src88 <= 12'h6f3;
        src89 <= 12'hdf0;
        src90 <= 12'hc64;
        src91 <= 12'hd33;
        src92 <= 12'h9b9;
        src93 <= 12'h3ce;
        src94 <= 12'h1f0;
        src95 <= 12'h2b1;
        src96 <= 12'h181;
        src97 <= 12'hb5c;
        src98 <= 12'h4c9;
        src99 <= 12'hdc8;
        src100 <= 12'h0;
        src101 <= 12'hc7c;
        src102 <= 12'hfaf;
        src103 <= 12'hbcd;
        src104 <= 12'hbb;
        src105 <= 12'h69d;
        src106 <= 12'h19c;
        src107 <= 12'h6ec;
        src108 <= 12'hfbd;
        src109 <= 12'h66e;
        src110 <= 12'h78;
        src111 <= 12'h543;
        src112 <= 12'h1a4;
        src113 <= 12'hab;
        src114 <= 12'h847;
        src115 <= 12'hb6d;
        src116 <= 12'hc96;
        src117 <= 12'h12d;
        src118 <= 12'heb7;
        src119 <= 12'h986;
        src120 <= 12'hc56;
        src121 <= 12'h6f5;
        src122 <= 12'he47;
        src123 <= 12'h7b;
        src124 <= 12'h6c2;
        src125 <= 12'he8b;
        src126 <= 12'h758;
        src127 <= 12'hc57;
        src128 <= 12'h7c4;
        src129 <= 12'hdde;
        src130 <= 12'h64d;
        src131 <= 12'hf86;
        src132 <= 12'hba2;
        src133 <= 12'h40c;
        src134 <= 12'h8ab;
        src135 <= 12'h4c0;
        src136 <= 12'h946;
        src137 <= 12'h98d;
        src138 <= 12'h23e;
        src139 <= 12'h18a;
        src140 <= 12'h903;
        src141 <= 12'h624;
        src142 <= 12'hc2e;
        src143 <= 12'he6a;
        src144 <= 12'hebf;
        src145 <= 12'h3e3;
        src146 <= 12'h7a8;
        src147 <= 12'hd35;
        src148 <= 12'h53b;
        src149 <= 12'ha5e;
        src150 <= 12'h2a1;
        src151 <= 12'hd9d;
        src152 <= 12'h414;
        src153 <= 12'h6dd;
        src154 <= 12'h88b;
        src155 <= 12'h176;
        src156 <= 12'h5c;
        src157 <= 12'hcd0;
        src158 <= 12'h2be;
        src159 <= 12'hd50;
        src160 <= 12'hf01;
        src161 <= 12'h3a5;
        exp <= 20'h505ed;
        #1
        src0 <= 12'h3f9;
        src1 <= 12'h23c;
        src2 <= 12'hbb5;
        src3 <= 12'h258;
        src4 <= 12'h16e;
        src5 <= 12'h672;
        src6 <= 12'hdf2;
        src7 <= 12'hfd3;
        src8 <= 12'hf7d;
        src9 <= 12'hff7;
        src10 <= 12'hde2;
        src11 <= 12'hf89;
        src12 <= 12'hfca;
        src13 <= 12'hfce;
        src14 <= 12'h1a9;
        src15 <= 12'hd5f;
        src16 <= 12'h7e;
        src17 <= 12'hf99;
        src18 <= 12'h7b6;
        src19 <= 12'h6b3;
        src20 <= 12'h9ab;
        src21 <= 12'ha32;
        src22 <= 12'ha4f;
        src23 <= 12'h38c;
        src24 <= 12'h7d9;
        src25 <= 12'h601;
        src26 <= 12'hdb8;
        src27 <= 12'h222;
        src28 <= 12'h9e6;
        src29 <= 12'h822;
        src30 <= 12'h224;
        src31 <= 12'hccb;
        src32 <= 12'h5f3;
        src33 <= 12'h3b9;
        src34 <= 12'h891;
        src35 <= 12'h87b;
        src36 <= 12'ha22;
        src37 <= 12'hac9;
        src38 <= 12'hfe9;
        src39 <= 12'hf62;
        src40 <= 12'hc5d;
        src41 <= 12'h26a;
        src42 <= 12'he47;
        src43 <= 12'hc00;
        src44 <= 12'h57e;
        src45 <= 12'h62c;
        src46 <= 12'hfb2;
        src47 <= 12'hf45;
        src48 <= 12'h64b;
        src49 <= 12'h8ae;
        src50 <= 12'h14;
        src51 <= 12'h4b4;
        src52 <= 12'h4b7;
        src53 <= 12'h53b;
        src54 <= 12'h54a;
        src55 <= 12'hcd2;
        src56 <= 12'h97e;
        src57 <= 12'h1c;
        src58 <= 12'h209;
        src59 <= 12'hbdc;
        src60 <= 12'h12;
        src61 <= 12'hda7;
        src62 <= 12'h868;
        src63 <= 12'h6e4;
        src64 <= 12'h23e;
        src65 <= 12'h7d0;
        src66 <= 12'h1ae;
        src67 <= 12'h211;
        src68 <= 12'hbed;
        src69 <= 12'h6f6;
        src70 <= 12'hb88;
        src71 <= 12'ha0b;
        src72 <= 12'h3d9;
        src73 <= 12'h7a9;
        src74 <= 12'h898;
        src75 <= 12'h906;
        src76 <= 12'h745;
        src77 <= 12'hedf;
        src78 <= 12'he0e;
        src79 <= 12'h546;
        src80 <= 12'h454;
        src81 <= 12'hbab;
        src82 <= 12'h52c;
        src83 <= 12'hdd4;
        src84 <= 12'h766;
        src85 <= 12'he35;
        src86 <= 12'hbc1;
        src87 <= 12'h4b5;
        src88 <= 12'h7a8;
        src89 <= 12'h475;
        src90 <= 12'hd4a;
        src91 <= 12'h932;
        src92 <= 12'h71f;
        src93 <= 12'hac1;
        src94 <= 12'heee;
        src95 <= 12'h846;
        src96 <= 12'hc64;
        src97 <= 12'h2e;
        src98 <= 12'h8b3;
        src99 <= 12'h13c;
        src100 <= 12'hf5c;
        src101 <= 12'hd8a;
        src102 <= 12'h21a;
        src103 <= 12'he73;
        src104 <= 12'he4c;
        src105 <= 12'hfe1;
        src106 <= 12'hdee;
        src107 <= 12'hfd4;
        src108 <= 12'h918;
        src109 <= 12'hc5f;
        src110 <= 12'h378;
        src111 <= 12'h4f1;
        src112 <= 12'h982;
        src113 <= 12'he8e;
        src114 <= 12'hba1;
        src115 <= 12'hca4;
        src116 <= 12'h670;
        src117 <= 12'ha68;
        src118 <= 12'h457;
        src119 <= 12'h9f7;
        src120 <= 12'h686;
        src121 <= 12'h5ce;
        src122 <= 12'h978;
        src123 <= 12'h98f;
        src124 <= 12'h303;
        src125 <= 12'h9aa;
        src126 <= 12'h2a8;
        src127 <= 12'hf2f;
        src128 <= 12'h941;
        src129 <= 12'h2b9;
        src130 <= 12'h3a8;
        src131 <= 12'h9bd;
        src132 <= 12'hdd9;
        src133 <= 12'hc07;
        src134 <= 12'hadf;
        src135 <= 12'hd29;
        src136 <= 12'h8e0;
        src137 <= 12'h990;
        src138 <= 12'h723;
        src139 <= 12'ha07;
        src140 <= 12'ha4;
        src141 <= 12'hfcc;
        src142 <= 12'h3bc;
        src143 <= 12'hf20;
        src144 <= 12'hb0;
        src145 <= 12'h407;
        src146 <= 12'ha6c;
        src147 <= 12'h235;
        src148 <= 12'h170;
        src149 <= 12'h97f;
        src150 <= 12'h2d6;
        src151 <= 12'h784;
        src152 <= 12'h33;
        src153 <= 12'h630;
        src154 <= 12'h522;
        src155 <= 12'h9d4;
        src156 <= 12'h8d3;
        src157 <= 12'h37b;
        src158 <= 12'he9e;
        src159 <= 12'h142;
        src160 <= 12'ha7a;
        src161 <= 12'hbe8;
        exp <= 20'h568a5;
        #1
        src0 <= 12'h344;
        src1 <= 12'h92b;
        src2 <= 12'hae6;
        src3 <= 12'h52e;
        src4 <= 12'h547;
        src5 <= 12'h9a1;
        src6 <= 12'hd8a;
        src7 <= 12'hce1;
        src8 <= 12'h88f;
        src9 <= 12'h3f1;
        src10 <= 12'hc13;
        src11 <= 12'h2fa;
        src12 <= 12'h9c1;
        src13 <= 12'hb5e;
        src14 <= 12'h1;
        src15 <= 12'hece;
        src16 <= 12'ha6a;
        src17 <= 12'hbcc;
        src18 <= 12'h996;
        src19 <= 12'ha47;
        src20 <= 12'h452;
        src21 <= 12'h3eb;
        src22 <= 12'h26b;
        src23 <= 12'hb73;
        src24 <= 12'h642;
        src25 <= 12'he51;
        src26 <= 12'h82f;
        src27 <= 12'h58e;
        src28 <= 12'ha05;
        src29 <= 12'h2da;
        src30 <= 12'h762;
        src31 <= 12'ha16;
        src32 <= 12'h4e9;
        src33 <= 12'h7f6;
        src34 <= 12'h192;
        src35 <= 12'hd49;
        src36 <= 12'hf49;
        src37 <= 12'hf98;
        src38 <= 12'h438;
        src39 <= 12'h583;
        src40 <= 12'hd56;
        src41 <= 12'h1d0;
        src42 <= 12'h3ac;
        src43 <= 12'h83f;
        src44 <= 12'h728;
        src45 <= 12'h9cb;
        src46 <= 12'hbe4;
        src47 <= 12'h7c5;
        src48 <= 12'hecc;
        src49 <= 12'h805;
        src50 <= 12'h2c1;
        src51 <= 12'h954;
        src52 <= 12'h9de;
        src53 <= 12'ha84;
        src54 <= 12'hfb9;
        src55 <= 12'h733;
        src56 <= 12'hd45;
        src57 <= 12'h8a7;
        src58 <= 12'h308;
        src59 <= 12'h978;
        src60 <= 12'h293;
        src61 <= 12'h140;
        src62 <= 12'h8f6;
        src63 <= 12'h895;
        src64 <= 12'he53;
        src65 <= 12'h956;
        src66 <= 12'he35;
        src67 <= 12'he45;
        src68 <= 12'h7e0;
        src69 <= 12'ha63;
        src70 <= 12'h7e;
        src71 <= 12'ha68;
        src72 <= 12'h6d0;
        src73 <= 12'hd63;
        src74 <= 12'h624;
        src75 <= 12'hee3;
        src76 <= 12'h741;
        src77 <= 12'h6f6;
        src78 <= 12'h44c;
        src79 <= 12'hfa7;
        src80 <= 12'h868;
        src81 <= 12'h460;
        src82 <= 12'h8c2;
        src83 <= 12'h5f6;
        src84 <= 12'hbd7;
        src85 <= 12'hfac;
        src86 <= 12'hdba;
        src87 <= 12'h98e;
        src88 <= 12'hb98;
        src89 <= 12'h6f5;
        src90 <= 12'h7da;
        src91 <= 12'ha21;
        src92 <= 12'h309;
        src93 <= 12'h369;
        src94 <= 12'h355;
        src95 <= 12'hd7f;
        src96 <= 12'h6ee;
        src97 <= 12'h8aa;
        src98 <= 12'hed;
        src99 <= 12'hf04;
        src100 <= 12'h5b;
        src101 <= 12'h849;
        src102 <= 12'hcee;
        src103 <= 12'hd;
        src104 <= 12'h930;
        src105 <= 12'hf7d;
        src106 <= 12'hfaa;
        src107 <= 12'hc0;
        src108 <= 12'h44b;
        src109 <= 12'hbd6;
        src110 <= 12'h8d2;
        src111 <= 12'h3d4;
        src112 <= 12'hb3e;
        src113 <= 12'h80;
        src114 <= 12'h698;
        src115 <= 12'h833;
        src116 <= 12'hc15;
        src117 <= 12'h5de;
        src118 <= 12'hed3;
        src119 <= 12'hba1;
        src120 <= 12'hf2c;
        src121 <= 12'ha1f;
        src122 <= 12'h409;
        src123 <= 12'h906;
        src124 <= 12'h400;
        src125 <= 12'h1a5;
        src126 <= 12'ha29;
        src127 <= 12'h857;
        src128 <= 12'h82f;
        src129 <= 12'h1a;
        src130 <= 12'h23f;
        src131 <= 12'h2a3;
        src132 <= 12'h62e;
        src133 <= 12'h98b;
        src134 <= 12'h2f;
        src135 <= 12'h3b4;
        src136 <= 12'h4a4;
        src137 <= 12'h796;
        src138 <= 12'hd6b;
        src139 <= 12'h25;
        src140 <= 12'h985;
        src141 <= 12'hfe5;
        src142 <= 12'h478;
        src143 <= 12'h77c;
        src144 <= 12'h818;
        src145 <= 12'h373;
        src146 <= 12'h35;
        src147 <= 12'h441;
        src148 <= 12'h551;
        src149 <= 12'hcc7;
        src150 <= 12'h440;
        src151 <= 12'h4da;
        src152 <= 12'h67c;
        src153 <= 12'h61e;
        src154 <= 12'h3f5;
        src155 <= 12'h978;
        src156 <= 12'h292;
        src157 <= 12'ha54;
        src158 <= 12'h440;
        src159 <= 12'h167;
        src160 <= 12'h2c7;
        src161 <= 12'h27a;
        exp <= 20'h4f45c;
        #1
        src0 <= 12'h5ca;
        src1 <= 12'hb0d;
        src2 <= 12'ha47;
        src3 <= 12'ha64;
        src4 <= 12'h4ab;
        src5 <= 12'hdd7;
        src6 <= 12'hcf9;
        src7 <= 12'hdc8;
        src8 <= 12'h2df;
        src9 <= 12'h99b;
        src10 <= 12'hc4;
        src11 <= 12'h2c1;
        src12 <= 12'h31b;
        src13 <= 12'h19e;
        src14 <= 12'h8ee;
        src15 <= 12'h73d;
        src16 <= 12'h2b9;
        src17 <= 12'h663;
        src18 <= 12'h718;
        src19 <= 12'h34b;
        src20 <= 12'h6bf;
        src21 <= 12'haf1;
        src22 <= 12'h307;
        src23 <= 12'hc1e;
        src24 <= 12'h38b;
        src25 <= 12'h31b;
        src26 <= 12'hef0;
        src27 <= 12'h266;
        src28 <= 12'hb1d;
        src29 <= 12'hcc6;
        src30 <= 12'h6d2;
        src31 <= 12'h843;
        src32 <= 12'h59a;
        src33 <= 12'h480;
        src34 <= 12'hb5e;
        src35 <= 12'ha06;
        src36 <= 12'h544;
        src37 <= 12'hdd0;
        src38 <= 12'h290;
        src39 <= 12'h782;
        src40 <= 12'hb62;
        src41 <= 12'hd62;
        src42 <= 12'h585;
        src43 <= 12'h413;
        src44 <= 12'haaf;
        src45 <= 12'h699;
        src46 <= 12'hc18;
        src47 <= 12'hafa;
        src48 <= 12'hb77;
        src49 <= 12'h365;
        src50 <= 12'h964;
        src51 <= 12'h927;
        src52 <= 12'hc6;
        src53 <= 12'hf72;
        src54 <= 12'h8da;
        src55 <= 12'ha91;
        src56 <= 12'h220;
        src57 <= 12'h11c;
        src58 <= 12'h8c9;
        src59 <= 12'haf4;
        src60 <= 12'hb0;
        src61 <= 12'hb46;
        src62 <= 12'h23c;
        src63 <= 12'h74f;
        src64 <= 12'h1f6;
        src65 <= 12'hc5;
        src66 <= 12'hd74;
        src67 <= 12'hb1b;
        src68 <= 12'h567;
        src69 <= 12'hd16;
        src70 <= 12'haa;
        src71 <= 12'hecf;
        src72 <= 12'h2ef;
        src73 <= 12'h62e;
        src74 <= 12'h510;
        src75 <= 12'hb65;
        src76 <= 12'h140;
        src77 <= 12'h4fd;
        src78 <= 12'h7d5;
        src79 <= 12'hfb0;
        src80 <= 12'h3a7;
        src81 <= 12'h3ea;
        src82 <= 12'h83b;
        src83 <= 12'h747;
        src84 <= 12'hd12;
        src85 <= 12'h56a;
        src86 <= 12'hf17;
        src87 <= 12'h20e;
        src88 <= 12'h7cb;
        src89 <= 12'h48d;
        src90 <= 12'ha75;
        src91 <= 12'hf46;
        src92 <= 12'h220;
        src93 <= 12'h1e6;
        src94 <= 12'hbf8;
        src95 <= 12'h4c4;
        src96 <= 12'h63e;
        src97 <= 12'h8cd;
        src98 <= 12'h1e6;
        src99 <= 12'h53f;
        src100 <= 12'h282;
        src101 <= 12'h395;
        src102 <= 12'h98a;
        src103 <= 12'h49f;
        src104 <= 12'hafc;
        src105 <= 12'heb1;
        src106 <= 12'h93b;
        src107 <= 12'hc0a;
        src108 <= 12'hc89;
        src109 <= 12'h3ca;
        src110 <= 12'h911;
        src111 <= 12'hcfe;
        src112 <= 12'hf3b;
        src113 <= 12'hada;
        src114 <= 12'h73f;
        src115 <= 12'h674;
        src116 <= 12'ha5d;
        src117 <= 12'h762;
        src118 <= 12'h1c6;
        src119 <= 12'hee2;
        src120 <= 12'h822;
        src121 <= 12'he40;
        src122 <= 12'h78;
        src123 <= 12'hcba;
        src124 <= 12'h64f;
        src125 <= 12'hf5a;
        src126 <= 12'ha2e;
        src127 <= 12'h5b2;
        src128 <= 12'h915;
        src129 <= 12'h597;
        src130 <= 12'h714;
        src131 <= 12'h48d;
        src132 <= 12'hecd;
        src133 <= 12'h461;
        src134 <= 12'h33b;
        src135 <= 12'had3;
        src136 <= 12'ha85;
        src137 <= 12'h1bd;
        src138 <= 12'hce4;
        src139 <= 12'hbb1;
        src140 <= 12'hc87;
        src141 <= 12'h639;
        src142 <= 12'h565;
        src143 <= 12'hf0a;
        src144 <= 12'h2d6;
        src145 <= 12'h47c;
        src146 <= 12'hf60;
        src147 <= 12'h201;
        src148 <= 12'h700;
        src149 <= 12'h95b;
        src150 <= 12'h598;
        src151 <= 12'ha1c;
        src152 <= 12'hc57;
        src153 <= 12'h425;
        src154 <= 12'heda;
        src155 <= 12'h5b;
        src156 <= 12'h4b7;
        src157 <= 12'h306;
        src158 <= 12'h999;
        src159 <= 12'h7fe;
        src160 <= 12'h5e1;
        src161 <= 12'hf34;
        exp <= 20'h4ef66;
        #1
        src0 <= 12'hbfa;
        src1 <= 12'hb3e;
        src2 <= 12'h559;
        src3 <= 12'h76;
        src4 <= 12'hb9e;
        src5 <= 12'h4d3;
        src6 <= 12'ha12;
        src7 <= 12'h96b;
        src8 <= 12'h388;
        src9 <= 12'hb4b;
        src10 <= 12'h815;
        src11 <= 12'h386;
        src12 <= 12'h29;
        src13 <= 12'h328;
        src14 <= 12'h8b9;
        src15 <= 12'h9b9;
        src16 <= 12'h6db;
        src17 <= 12'hfa6;
        src18 <= 12'hfe2;
        src19 <= 12'h155;
        src20 <= 12'h3ae;
        src21 <= 12'h390;
        src22 <= 12'h2d9;
        src23 <= 12'h482;
        src24 <= 12'h179;
        src25 <= 12'h29a;
        src26 <= 12'h658;
        src27 <= 12'h384;
        src28 <= 12'hb90;
        src29 <= 12'ha8b;
        src30 <= 12'h227;
        src31 <= 12'h7ad;
        src32 <= 12'he78;
        src33 <= 12'h259;
        src34 <= 12'h4ca;
        src35 <= 12'h98d;
        src36 <= 12'h6dd;
        src37 <= 12'h2e7;
        src38 <= 12'haca;
        src39 <= 12'hb5b;
        src40 <= 12'h5f4;
        src41 <= 12'hced;
        src42 <= 12'h8e5;
        src43 <= 12'h6a1;
        src44 <= 12'hfdc;
        src45 <= 12'h11e;
        src46 <= 12'h3df;
        src47 <= 12'hd31;
        src48 <= 12'he66;
        src49 <= 12'h610;
        src50 <= 12'h538;
        src51 <= 12'h8f0;
        src52 <= 12'h422;
        src53 <= 12'h6d5;
        src54 <= 12'h828;
        src55 <= 12'h83a;
        src56 <= 12'h926;
        src57 <= 12'hef;
        src58 <= 12'h16;
        src59 <= 12'had2;
        src60 <= 12'h66c;
        src61 <= 12'hf7b;
        src62 <= 12'h922;
        src63 <= 12'h94a;
        src64 <= 12'h51a;
        src65 <= 12'h227;
        src66 <= 12'hd9f;
        src67 <= 12'h7e4;
        src68 <= 12'hd08;
        src69 <= 12'hff0;
        src70 <= 12'h1f2;
        src71 <= 12'h8da;
        src72 <= 12'ha63;
        src73 <= 12'ha5e;
        src74 <= 12'hc7a;
        src75 <= 12'he64;
        src76 <= 12'h170;
        src77 <= 12'he94;
        src78 <= 12'h45f;
        src79 <= 12'hb95;
        src80 <= 12'h76f;
        src81 <= 12'h18a;
        src82 <= 12'hef6;
        src83 <= 12'hec9;
        src84 <= 12'h515;
        src85 <= 12'h784;
        src86 <= 12'hb1b;
        src87 <= 12'hfdd;
        src88 <= 12'h790;
        src89 <= 12'h184;
        src90 <= 12'hbf7;
        src91 <= 12'h181;
        src92 <= 12'h96e;
        src93 <= 12'hc1;
        src94 <= 12'ha47;
        src95 <= 12'h15d;
        src96 <= 12'h3c1;
        src97 <= 12'hc35;
        src98 <= 12'h620;
        src99 <= 12'h5c7;
        src100 <= 12'h2d4;
        src101 <= 12'h31c;
        src102 <= 12'h334;
        src103 <= 12'h5da;
        src104 <= 12'hf40;
        src105 <= 12'h2bc;
        src106 <= 12'h283;
        src107 <= 12'hae9;
        src108 <= 12'hca3;
        src109 <= 12'h56f;
        src110 <= 12'h2a7;
        src111 <= 12'h862;
        src112 <= 12'h757;
        src113 <= 12'h24f;
        src114 <= 12'h450;
        src115 <= 12'h589;
        src116 <= 12'h33f;
        src117 <= 12'h6a9;
        src118 <= 12'h13c;
        src119 <= 12'had7;
        src120 <= 12'h9f9;
        src121 <= 12'hce2;
        src122 <= 12'h5a5;
        src123 <= 12'h40c;
        src124 <= 12'h6fb;
        src125 <= 12'hd30;
        src126 <= 12'hb2f;
        src127 <= 12'hf99;
        src128 <= 12'hded;
        src129 <= 12'hb6d;
        src130 <= 12'had8;
        src131 <= 12'h759;
        src132 <= 12'h40a;
        src133 <= 12'h93;
        src134 <= 12'h442;
        src135 <= 12'h586;
        src136 <= 12'hc5d;
        src137 <= 12'h5bd;
        src138 <= 12'h37d;
        src139 <= 12'h39e;
        src140 <= 12'h153;
        src141 <= 12'h828;
        src142 <= 12'hc87;
        src143 <= 12'h20c;
        src144 <= 12'hc3e;
        src145 <= 12'hd33;
        src146 <= 12'h27c;
        src147 <= 12'ha62;
        src148 <= 12'he7e;
        src149 <= 12'h36a;
        src150 <= 12'h177;
        src151 <= 12'h481;
        src152 <= 12'h22c;
        src153 <= 12'h107;
        src154 <= 12'he4c;
        src155 <= 12'hd2a;
        src156 <= 12'hdf4;
        src157 <= 12'hf34;
        src158 <= 12'h536;
        src159 <= 12'hfbb;
        src160 <= 12'h51e;
        src161 <= 12'hb7d;
        exp <= 20'h4cdfb;
        #1
        src0 <= 12'h373;
        src1 <= 12'h8f;
        src2 <= 12'h359;
        src3 <= 12'hf72;
        src4 <= 12'h19f;
        src5 <= 12'haee;
        src6 <= 12'h2c2;
        src7 <= 12'h302;
        src8 <= 12'h4f3;
        src9 <= 12'h248;
        src10 <= 12'h7c0;
        src11 <= 12'h559;
        src12 <= 12'hc17;
        src13 <= 12'hd5;
        src14 <= 12'h2cc;
        src15 <= 12'h849;
        src16 <= 12'h2c7;
        src17 <= 12'hdac;
        src18 <= 12'h7bd;
        src19 <= 12'hccb;
        src20 <= 12'he93;
        src21 <= 12'hd25;
        src22 <= 12'h35b;
        src23 <= 12'hfde;
        src24 <= 12'h13b;
        src25 <= 12'hf8c;
        src26 <= 12'hc4b;
        src27 <= 12'h46f;
        src28 <= 12'h6fe;
        src29 <= 12'h4f0;
        src30 <= 12'h9e6;
        src31 <= 12'he42;
        src32 <= 12'h294;
        src33 <= 12'h61f;
        src34 <= 12'h805;
        src35 <= 12'h9a7;
        src36 <= 12'he3d;
        src37 <= 12'h8e6;
        src38 <= 12'h97c;
        src39 <= 12'hd5b;
        src40 <= 12'h75c;
        src41 <= 12'ha33;
        src42 <= 12'h461;
        src43 <= 12'ha31;
        src44 <= 12'h9e6;
        src45 <= 12'hc1;
        src46 <= 12'h185;
        src47 <= 12'hf2b;
        src48 <= 12'h218;
        src49 <= 12'ha82;
        src50 <= 12'h4b2;
        src51 <= 12'h403;
        src52 <= 12'hdd0;
        src53 <= 12'h76d;
        src54 <= 12'h139;
        src55 <= 12'h2fd;
        src56 <= 12'h678;
        src57 <= 12'hc0;
        src58 <= 12'h7d9;
        src59 <= 12'h582;
        src60 <= 12'h65f;
        src61 <= 12'hb6d;
        src62 <= 12'h345;
        src63 <= 12'h599;
        src64 <= 12'h6d;
        src65 <= 12'h2bb;
        src66 <= 12'h158;
        src67 <= 12'hc0c;
        src68 <= 12'h243;
        src69 <= 12'haad;
        src70 <= 12'hb7f;
        src71 <= 12'hee8;
        src72 <= 12'hcde;
        src73 <= 12'haba;
        src74 <= 12'h514;
        src75 <= 12'hb24;
        src76 <= 12'h40c;
        src77 <= 12'h81a;
        src78 <= 12'h541;
        src79 <= 12'h741;
        src80 <= 12'h20f;
        src81 <= 12'h9;
        src82 <= 12'h227;
        src83 <= 12'h5f7;
        src84 <= 12'h7d;
        src85 <= 12'h7d3;
        src86 <= 12'h925;
        src87 <= 12'h1d5;
        src88 <= 12'h606;
        src89 <= 12'h637;
        src90 <= 12'ha91;
        src91 <= 12'h4ac;
        src92 <= 12'hbba;
        src93 <= 12'h893;
        src94 <= 12'h390;
        src95 <= 12'hb3a;
        src96 <= 12'h2f4;
        src97 <= 12'h88f;
        src98 <= 12'hf63;
        src99 <= 12'h724;
        src100 <= 12'h838;
        src101 <= 12'h91d;
        src102 <= 12'hc81;
        src103 <= 12'hfa4;
        src104 <= 12'h451;
        src105 <= 12'h98a;
        src106 <= 12'hdd7;
        src107 <= 12'h9f1;
        src108 <= 12'hbcc;
        src109 <= 12'hecb;
        src110 <= 12'hf4;
        src111 <= 12'hb29;
        src112 <= 12'h865;
        src113 <= 12'he7b;
        src114 <= 12'h686;
        src115 <= 12'hebf;
        src116 <= 12'h74b;
        src117 <= 12'hd37;
        src118 <= 12'h620;
        src119 <= 12'h152;
        src120 <= 12'hb96;
        src121 <= 12'h9c4;
        src122 <= 12'ha02;
        src123 <= 12'h2d8;
        src124 <= 12'h8d3;
        src125 <= 12'h396;
        src126 <= 12'h163;
        src127 <= 12'hb8d;
        src128 <= 12'h13;
        src129 <= 12'hc04;
        src130 <= 12'h620;
        src131 <= 12'hc81;
        src132 <= 12'h828;
        src133 <= 12'hc4c;
        src134 <= 12'hcec;
        src135 <= 12'hb95;
        src136 <= 12'haf3;
        src137 <= 12'h609;
        src138 <= 12'hc6d;
        src139 <= 12'haa1;
        src140 <= 12'h543;
        src141 <= 12'h608;
        src142 <= 12'h687;
        src143 <= 12'hbd7;
        src144 <= 12'h4c;
        src145 <= 12'h6c1;
        src146 <= 12'h2ea;
        src147 <= 12'h58a;
        src148 <= 12'hde9;
        src149 <= 12'h36b;
        src150 <= 12'h92d;
        src151 <= 12'h3ca;
        src152 <= 12'hae7;
        src153 <= 12'hd87;
        src154 <= 12'h20f;
        src155 <= 12'h3f7;
        src156 <= 12'hf52;
        src157 <= 12'h567;
        src158 <= 12'h7fd;
        src159 <= 12'he28;
        src160 <= 12'h19;
        src161 <= 12'h4d5;
        exp <= 20'h4d21f;
        #1
        src0 <= 12'h45;
        src1 <= 12'h728;
        src2 <= 12'hdfe;
        src3 <= 12'h7aa;
        src4 <= 12'h255;
        src5 <= 12'hb69;
        src6 <= 12'h307;
        src7 <= 12'hb4a;
        src8 <= 12'hf8d;
        src9 <= 12'h143;
        src10 <= 12'h64c;
        src11 <= 12'hb1f;
        src12 <= 12'hf49;
        src13 <= 12'h878;
        src14 <= 12'h19e;
        src15 <= 12'h140;
        src16 <= 12'h62d;
        src17 <= 12'h583;
        src18 <= 12'hb9a;
        src19 <= 12'h8d4;
        src20 <= 12'h910;
        src21 <= 12'hef;
        src22 <= 12'h6a8;
        src23 <= 12'h674;
        src24 <= 12'h437;
        src25 <= 12'h620;
        src26 <= 12'h9f3;
        src27 <= 12'h49;
        src28 <= 12'he9d;
        src29 <= 12'h8af;
        src30 <= 12'h35b;
        src31 <= 12'hc2b;
        src32 <= 12'h4a9;
        src33 <= 12'h5d7;
        src34 <= 12'h540;
        src35 <= 12'h651;
        src36 <= 12'he80;
        src37 <= 12'h5e9;
        src38 <= 12'hfa3;
        src39 <= 12'hc01;
        src40 <= 12'h5a8;
        src41 <= 12'hb95;
        src42 <= 12'hf71;
        src43 <= 12'hfb0;
        src44 <= 12'haf4;
        src45 <= 12'h3d6;
        src46 <= 12'hdb0;
        src47 <= 12'h7ab;
        src48 <= 12'h892;
        src49 <= 12'hdd9;
        src50 <= 12'h694;
        src51 <= 12'h579;
        src52 <= 12'haa4;
        src53 <= 12'hb2c;
        src54 <= 12'h753;
        src55 <= 12'h296;
        src56 <= 12'h717;
        src57 <= 12'ha4a;
        src58 <= 12'h38;
        src59 <= 12'h4f6;
        src60 <= 12'hc20;
        src61 <= 12'h16a;
        src62 <= 12'hdf4;
        src63 <= 12'h65a;
        src64 <= 12'hb54;
        src65 <= 12'he26;
        src66 <= 12'hac5;
        src67 <= 12'h134;
        src68 <= 12'h888;
        src69 <= 12'h88;
        src70 <= 12'hdb6;
        src71 <= 12'hbb7;
        src72 <= 12'h924;
        src73 <= 12'h943;
        src74 <= 12'he93;
        src75 <= 12'haba;
        src76 <= 12'h59c;
        src77 <= 12'ha56;
        src78 <= 12'h87f;
        src79 <= 12'h113;
        src80 <= 12'hbd4;
        src81 <= 12'h12e;
        src82 <= 12'h7b1;
        src83 <= 12'h62d;
        src84 <= 12'h935;
        src85 <= 12'h842;
        src86 <= 12'hd7a;
        src87 <= 12'h1f0;
        src88 <= 12'hef2;
        src89 <= 12'h496;
        src90 <= 12'h501;
        src91 <= 12'h70e;
        src92 <= 12'h385;
        src93 <= 12'h9cb;
        src94 <= 12'h7f2;
        src95 <= 12'hcf9;
        src96 <= 12'h7c7;
        src97 <= 12'h176;
        src98 <= 12'hba8;
        src99 <= 12'he67;
        src100 <= 12'hcf6;
        src101 <= 12'h62a;
        src102 <= 12'h711;
        src103 <= 12'hbe1;
        src104 <= 12'h3de;
        src105 <= 12'h695;
        src106 <= 12'hcf;
        src107 <= 12'h46e;
        src108 <= 12'he9f;
        src109 <= 12'hea9;
        src110 <= 12'hd9b;
        src111 <= 12'h5f1;
        src112 <= 12'h20;
        src113 <= 12'h19b;
        src114 <= 12'hd6b;
        src115 <= 12'h324;
        src116 <= 12'h4a4;
        src117 <= 12'hff2;
        src118 <= 12'hcf2;
        src119 <= 12'hd84;
        src120 <= 12'ha9b;
        src121 <= 12'h5c1;
        src122 <= 12'he1c;
        src123 <= 12'h2eb;
        src124 <= 12'h7e;
        src125 <= 12'h3b9;
        src126 <= 12'h413;
        src127 <= 12'hc5b;
        src128 <= 12'h850;
        src129 <= 12'hbf8;
        src130 <= 12'h111;
        src131 <= 12'hef3;
        src132 <= 12'hfa0;
        src133 <= 12'h23d;
        src134 <= 12'h3c3;
        src135 <= 12'h4b8;
        src136 <= 12'h4db;
        src137 <= 12'h773;
        src138 <= 12'h793;
        src139 <= 12'hdc0;
        src140 <= 12'h791;
        src141 <= 12'he4f;
        src142 <= 12'h8f5;
        src143 <= 12'h785;
        src144 <= 12'h570;
        src145 <= 12'ha36;
        src146 <= 12'hd9b;
        src147 <= 12'habb;
        src148 <= 12'h7b5;
        src149 <= 12'h45a;
        src150 <= 12'h147;
        src151 <= 12'h142;
        src152 <= 12'h565;
        src153 <= 12'h697;
        src154 <= 12'hbe5;
        src155 <= 12'hc6b;
        src156 <= 12'h838;
        src157 <= 12'h4a0;
        src158 <= 12'h353;
        src159 <= 12'h121;
        src160 <= 12'h494;
        src161 <= 12'hc38;
        exp <= 20'h50d67;
        #1
        src0 <= 12'ha9b;
        src1 <= 12'h18f;
        src2 <= 12'hd03;
        src3 <= 12'he9e;
        src4 <= 12'h984;
        src5 <= 12'h598;
        src6 <= 12'h21d;
        src7 <= 12'h649;
        src8 <= 12'h2e2;
        src9 <= 12'h582;
        src10 <= 12'hb15;
        src11 <= 12'h39f;
        src12 <= 12'h565;
        src13 <= 12'h88e;
        src14 <= 12'hcd;
        src15 <= 12'h66b;
        src16 <= 12'h33e;
        src17 <= 12'h8dd;
        src18 <= 12'h3ad;
        src19 <= 12'h42d;
        src20 <= 12'hc28;
        src21 <= 12'hba1;
        src22 <= 12'h706;
        src23 <= 12'h86e;
        src24 <= 12'h9d0;
        src25 <= 12'h6cd;
        src26 <= 12'hb07;
        src27 <= 12'h506;
        src28 <= 12'h857;
        src29 <= 12'hed6;
        src30 <= 12'h43b;
        src31 <= 12'h76;
        src32 <= 12'hc42;
        src33 <= 12'hadc;
        src34 <= 12'h250;
        src35 <= 12'hc7c;
        src36 <= 12'h835;
        src37 <= 12'hd7c;
        src38 <= 12'hb4a;
        src39 <= 12'hb17;
        src40 <= 12'h26e;
        src41 <= 12'h77e;
        src42 <= 12'hbbd;
        src43 <= 12'h87c;
        src44 <= 12'hd01;
        src45 <= 12'h726;
        src46 <= 12'h8e7;
        src47 <= 12'h490;
        src48 <= 12'h49d;
        src49 <= 12'h145;
        src50 <= 12'hb7c;
        src51 <= 12'hc9a;
        src52 <= 12'h8a;
        src53 <= 12'hcec;
        src54 <= 12'h4a4;
        src55 <= 12'ha79;
        src56 <= 12'hbe2;
        src57 <= 12'hd7e;
        src58 <= 12'h20e;
        src59 <= 12'h92e;
        src60 <= 12'heb5;
        src61 <= 12'h741;
        src62 <= 12'heae;
        src63 <= 12'h82c;
        src64 <= 12'h123;
        src65 <= 12'h839;
        src66 <= 12'h8ca;
        src67 <= 12'hbe5;
        src68 <= 12'h7fc;
        src69 <= 12'hc1b;
        src70 <= 12'h8a;
        src71 <= 12'h992;
        src72 <= 12'hee7;
        src73 <= 12'h2;
        src74 <= 12'he94;
        src75 <= 12'h9c1;
        src76 <= 12'hb1b;
        src77 <= 12'hb7c;
        src78 <= 12'h2d1;
        src79 <= 12'hd1;
        src80 <= 12'h3ba;
        src81 <= 12'h90c;
        src82 <= 12'hcfe;
        src83 <= 12'hfad;
        src84 <= 12'h3b0;
        src85 <= 12'hd18;
        src86 <= 12'ha78;
        src87 <= 12'h8b6;
        src88 <= 12'hca3;
        src89 <= 12'hbc0;
        src90 <= 12'h18b;
        src91 <= 12'h6c5;
        src92 <= 12'h8d3;
        src93 <= 12'he42;
        src94 <= 12'h449;
        src95 <= 12'hb2;
        src96 <= 12'hf21;
        src97 <= 12'h60b;
        src98 <= 12'hdff;
        src99 <= 12'hd;
        src100 <= 12'hc31;
        src101 <= 12'h898;
        src102 <= 12'h745;
        src103 <= 12'h87b;
        src104 <= 12'h758;
        src105 <= 12'h30d;
        src106 <= 12'hed;
        src107 <= 12'ha8b;
        src108 <= 12'hbb9;
        src109 <= 12'hea4;
        src110 <= 12'he67;
        src111 <= 12'he8;
        src112 <= 12'h301;
        src113 <= 12'hf51;
        src114 <= 12'h67;
        src115 <= 12'ha9b;
        src116 <= 12'haba;
        src117 <= 12'h4db;
        src118 <= 12'h209;
        src119 <= 12'h95d;
        src120 <= 12'h846;
        src121 <= 12'hbd7;
        src122 <= 12'h7a3;
        src123 <= 12'hafa;
        src124 <= 12'h198;
        src125 <= 12'hc4c;
        src126 <= 12'h4ee;
        src127 <= 12'h875;
        src128 <= 12'h97e;
        src129 <= 12'hb0b;
        src130 <= 12'h421;
        src131 <= 12'h9b5;
        src132 <= 12'h8d7;
        src133 <= 12'h6cc;
        src134 <= 12'hc73;
        src135 <= 12'hfde;
        src136 <= 12'hb6f;
        src137 <= 12'hc90;
        src138 <= 12'h759;
        src139 <= 12'ha5f;
        src140 <= 12'h5f5;
        src141 <= 12'hdc3;
        src142 <= 12'hb87;
        src143 <= 12'hea2;
        src144 <= 12'hd4f;
        src145 <= 12'h434;
        src146 <= 12'h324;
        src147 <= 12'h699;
        src148 <= 12'hb08;
        src149 <= 12'hd16;
        src150 <= 12'h91c;
        src151 <= 12'h862;
        src152 <= 12'hc4e;
        src153 <= 12'h571;
        src154 <= 12'h1f3;
        src155 <= 12'ha89;
        src156 <= 12'h99d;
        src157 <= 12'hd62;
        src158 <= 12'h41c;
        src159 <= 12'hbf5;
        src160 <= 12'hd61;
        src161 <= 12'h509;
        exp <= 20'h54cf5;
        #1
        src0 <= 12'hdbd;
        src1 <= 12'h751;
        src2 <= 12'h7a9;
        src3 <= 12'hb1c;
        src4 <= 12'hbd5;
        src5 <= 12'h5bb;
        src6 <= 12'h820;
        src7 <= 12'hc4;
        src8 <= 12'haed;
        src9 <= 12'h345;
        src10 <= 12'h7fe;
        src11 <= 12'h293;
        src12 <= 12'h1a9;
        src13 <= 12'h94;
        src14 <= 12'h3d1;
        src15 <= 12'hf83;
        src16 <= 12'heae;
        src17 <= 12'h7f4;
        src18 <= 12'h323;
        src19 <= 12'hdac;
        src20 <= 12'h116;
        src21 <= 12'h42;
        src22 <= 12'h56e;
        src23 <= 12'h25b;
        src24 <= 12'hb99;
        src25 <= 12'hdcd;
        src26 <= 12'hb31;
        src27 <= 12'h398;
        src28 <= 12'hdc;
        src29 <= 12'h1f3;
        src30 <= 12'hb78;
        src31 <= 12'h72;
        src32 <= 12'hb74;
        src33 <= 12'hc83;
        src34 <= 12'h60a;
        src35 <= 12'h75c;
        src36 <= 12'h7fc;
        src37 <= 12'h466;
        src38 <= 12'he50;
        src39 <= 12'h142;
        src40 <= 12'hf75;
        src41 <= 12'hb34;
        src42 <= 12'h51f;
        src43 <= 12'hbf7;
        src44 <= 12'hb45;
        src45 <= 12'h175;
        src46 <= 12'h8f7;
        src47 <= 12'h5b9;
        src48 <= 12'he0b;
        src49 <= 12'hac4;
        src50 <= 12'h307;
        src51 <= 12'h535;
        src52 <= 12'hf45;
        src53 <= 12'ha59;
        src54 <= 12'hed3;
        src55 <= 12'hdd8;
        src56 <= 12'h7b2;
        src57 <= 12'h1ef;
        src58 <= 12'h1eb;
        src59 <= 12'ha72;
        src60 <= 12'hcbd;
        src61 <= 12'ha1e;
        src62 <= 12'h8b9;
        src63 <= 12'h5f3;
        src64 <= 12'h933;
        src65 <= 12'h38a;
        src66 <= 12'hfbc;
        src67 <= 12'h3d7;
        src68 <= 12'haed;
        src69 <= 12'hd52;
        src70 <= 12'h5b4;
        src71 <= 12'hca2;
        src72 <= 12'hce4;
        src73 <= 12'h28b;
        src74 <= 12'h355;
        src75 <= 12'h538;
        src76 <= 12'h26e;
        src77 <= 12'hb64;
        src78 <= 12'h5ca;
        src79 <= 12'h6d;
        src80 <= 12'h8e8;
        src81 <= 12'h986;
        src82 <= 12'hb78;
        src83 <= 12'h6ba;
        src84 <= 12'h86e;
        src85 <= 12'hab8;
        src86 <= 12'h6ae;
        src87 <= 12'hc23;
        src88 <= 12'h703;
        src89 <= 12'hd87;
        src90 <= 12'hf22;
        src91 <= 12'h657;
        src92 <= 12'h5f3;
        src93 <= 12'h7ce;
        src94 <= 12'hfa9;
        src95 <= 12'hee8;
        src96 <= 12'h285;
        src97 <= 12'hb44;
        src98 <= 12'h32f;
        src99 <= 12'hcb5;
        src100 <= 12'ha6d;
        src101 <= 12'h21e;
        src102 <= 12'hb2f;
        src103 <= 12'h3b;
        src104 <= 12'ha5;
        src105 <= 12'hff1;
        src106 <= 12'h9a8;
        src107 <= 12'hcb3;
        src108 <= 12'h28d;
        src109 <= 12'he7;
        src110 <= 12'hee3;
        src111 <= 12'h774;
        src112 <= 12'h50f;
        src113 <= 12'h7ce;
        src114 <= 12'hd35;
        src115 <= 12'ha3a;
        src116 <= 12'hef0;
        src117 <= 12'h3c2;
        src118 <= 12'h4fc;
        src119 <= 12'h542;
        src120 <= 12'h3cc;
        src121 <= 12'he63;
        src122 <= 12'h648;
        src123 <= 12'h3a;
        src124 <= 12'hac;
        src125 <= 12'hdbb;
        src126 <= 12'h53;
        src127 <= 12'hca3;
        src128 <= 12'hca0;
        src129 <= 12'hcc9;
        src130 <= 12'h384;
        src131 <= 12'h661;
        src132 <= 12'he25;
        src133 <= 12'h15;
        src134 <= 12'h2dd;
        src135 <= 12'h1d9;
        src136 <= 12'h193;
        src137 <= 12'h9ae;
        src138 <= 12'h59e;
        src139 <= 12'haa6;
        src140 <= 12'h2ee;
        src141 <= 12'h102;
        src142 <= 12'h9e0;
        src143 <= 12'h246;
        src144 <= 12'he04;
        src145 <= 12'hd6a;
        src146 <= 12'hc1d;
        src147 <= 12'h4a5;
        src148 <= 12'hd11;
        src149 <= 12'h934;
        src150 <= 12'h5e;
        src151 <= 12'hd8d;
        src152 <= 12'h523;
        src153 <= 12'h940;
        src154 <= 12'hfb7;
        src155 <= 12'h203;
        src156 <= 12'h49c;
        src157 <= 12'hf50;
        src158 <= 12'hb6d;
        src159 <= 12'h5d8;
        src160 <= 12'h17b;
        src161 <= 12'h201;
        exp <= 20'h4f1e9;
        #1
        src0 <= 12'hc3f;
        src1 <= 12'h5ee;
        src2 <= 12'h50e;
        src3 <= 12'hfb5;
        src4 <= 12'he31;
        src5 <= 12'h272;
        src6 <= 12'h8d0;
        src7 <= 12'h4a8;
        src8 <= 12'hf0;
        src9 <= 12'h3d6;
        src10 <= 12'hf36;
        src11 <= 12'h18f;
        src12 <= 12'hc9c;
        src13 <= 12'h363;
        src14 <= 12'hd4f;
        src15 <= 12'h65a;
        src16 <= 12'h863;
        src17 <= 12'h46;
        src18 <= 12'ha31;
        src19 <= 12'hb88;
        src20 <= 12'hf15;
        src21 <= 12'h9e6;
        src22 <= 12'h314;
        src23 <= 12'he7a;
        src24 <= 12'hbd;
        src25 <= 12'h168;
        src26 <= 12'h594;
        src27 <= 12'h7b5;
        src28 <= 12'h23d;
        src29 <= 12'heec;
        src30 <= 12'h7c0;
        src31 <= 12'hc1e;
        src32 <= 12'hbe3;
        src33 <= 12'hfe5;
        src34 <= 12'h87a;
        src35 <= 12'h52f;
        src36 <= 12'hdd5;
        src37 <= 12'haf;
        src38 <= 12'h418;
        src39 <= 12'h671;
        src40 <= 12'hd92;
        src41 <= 12'h3eb;
        src42 <= 12'hdc2;
        src43 <= 12'h4aa;
        src44 <= 12'h542;
        src45 <= 12'he32;
        src46 <= 12'hd76;
        src47 <= 12'h265;
        src48 <= 12'h230;
        src49 <= 12'hdf1;
        src50 <= 12'h972;
        src51 <= 12'hdf5;
        src52 <= 12'hd6b;
        src53 <= 12'h2b0;
        src54 <= 12'h921;
        src55 <= 12'h88a;
        src56 <= 12'h8fa;
        src57 <= 12'hbea;
        src58 <= 12'he0a;
        src59 <= 12'he26;
        src60 <= 12'h2f;
        src61 <= 12'hec5;
        src62 <= 12'h2;
        src63 <= 12'h5e0;
        src64 <= 12'hecc;
        src65 <= 12'hf41;
        src66 <= 12'h3b7;
        src67 <= 12'h711;
        src68 <= 12'hd05;
        src69 <= 12'h3ed;
        src70 <= 12'h31c;
        src71 <= 12'h5f4;
        src72 <= 12'had0;
        src73 <= 12'he0d;
        src74 <= 12'h1d5;
        src75 <= 12'h544;
        src76 <= 12'h49f;
        src77 <= 12'hd5;
        src78 <= 12'hc8a;
        src79 <= 12'hb8b;
        src80 <= 12'h2f1;
        src81 <= 12'ha22;
        src82 <= 12'h75c;
        src83 <= 12'h3e0;
        src84 <= 12'h357;
        src85 <= 12'h8ba;
        src86 <= 12'hf6f;
        src87 <= 12'h76b;
        src88 <= 12'h7ad;
        src89 <= 12'h617;
        src90 <= 12'h3e2;
        src91 <= 12'h59a;
        src92 <= 12'hccf;
        src93 <= 12'h79c;
        src94 <= 12'haae;
        src95 <= 12'hbe4;
        src96 <= 12'h577;
        src97 <= 12'hbf9;
        src98 <= 12'h4eb;
        src99 <= 12'hf7;
        src100 <= 12'haf3;
        src101 <= 12'hc90;
        src102 <= 12'h601;
        src103 <= 12'hd7e;
        src104 <= 12'h740;
        src105 <= 12'hf31;
        src106 <= 12'h6be;
        src107 <= 12'hf89;
        src108 <= 12'h885;
        src109 <= 12'h245;
        src110 <= 12'h766;
        src111 <= 12'hc45;
        src112 <= 12'h2bd;
        src113 <= 12'he2d;
        src114 <= 12'h9fc;
        src115 <= 12'h363;
        src116 <= 12'hf9d;
        src117 <= 12'h5d2;
        src118 <= 12'h481;
        src119 <= 12'h12e;
        src120 <= 12'hb53;
        src121 <= 12'h58c;
        src122 <= 12'h610;
        src123 <= 12'hf2e;
        src124 <= 12'h202;
        src125 <= 12'he62;
        src126 <= 12'hb6;
        src127 <= 12'h1cd;
        src128 <= 12'hbea;
        src129 <= 12'h393;
        src130 <= 12'he93;
        src131 <= 12'h9ce;
        src132 <= 12'h8be;
        src133 <= 12'hb47;
        src134 <= 12'ha0;
        src135 <= 12'h91c;
        src136 <= 12'h27c;
        src137 <= 12'h673;
        src138 <= 12'h447;
        src139 <= 12'hf36;
        src140 <= 12'h66e;
        src141 <= 12'h4e0;
        src142 <= 12'h988;
        src143 <= 12'ha77;
        src144 <= 12'h980;
        src145 <= 12'hae8;
        src146 <= 12'h6a4;
        src147 <= 12'hf5b;
        src148 <= 12'h91b;
        src149 <= 12'hbed;
        src150 <= 12'h7ac;
        src151 <= 12'hd37;
        src152 <= 12'hc56;
        src153 <= 12'h680;
        src154 <= 12'h19f;
        src155 <= 12'h171;
        src156 <= 12'ha71;
        src157 <= 12'h207;
        src158 <= 12'h2d9;
        src159 <= 12'h4ae;
        src160 <= 12'h909;
        src161 <= 12'h7dc;
        exp <= 20'h522b9;
        #1
        src0 <= 12'hcad;
        src1 <= 12'h6e;
        src2 <= 12'h63b;
        src3 <= 12'hc2c;
        src4 <= 12'hd65;
        src5 <= 12'h6b0;
        src6 <= 12'hb38;
        src7 <= 12'h1db;
        src8 <= 12'h7c1;
        src9 <= 12'h48e;
        src10 <= 12'h47;
        src11 <= 12'h312;
        src12 <= 12'h1be;
        src13 <= 12'ha34;
        src14 <= 12'h5ef;
        src15 <= 12'h63e;
        src16 <= 12'ha8b;
        src17 <= 12'h4a7;
        src18 <= 12'he77;
        src19 <= 12'h8de;
        src20 <= 12'hf00;
        src21 <= 12'hc41;
        src22 <= 12'h105;
        src23 <= 12'h973;
        src24 <= 12'hb81;
        src25 <= 12'h133;
        src26 <= 12'h45e;
        src27 <= 12'h3ea;
        src28 <= 12'h429;
        src29 <= 12'hb92;
        src30 <= 12'h9a0;
        src31 <= 12'h7fd;
        src32 <= 12'ha0b;
        src33 <= 12'hbae;
        src34 <= 12'hc2;
        src35 <= 12'hb10;
        src36 <= 12'h44d;
        src37 <= 12'ha35;
        src38 <= 12'he4b;
        src39 <= 12'he94;
        src40 <= 12'h90f;
        src41 <= 12'h273;
        src42 <= 12'ha3c;
        src43 <= 12'hac4;
        src44 <= 12'h1e9;
        src45 <= 12'h2e9;
        src46 <= 12'hbff;
        src47 <= 12'hd76;
        src48 <= 12'h680;
        src49 <= 12'h947;
        src50 <= 12'h2c4;
        src51 <= 12'had9;
        src52 <= 12'hdd7;
        src53 <= 12'hd81;
        src54 <= 12'h6c1;
        src55 <= 12'hf54;
        src56 <= 12'h3a2;
        src57 <= 12'hf21;
        src58 <= 12'h8d4;
        src59 <= 12'h757;
        src60 <= 12'hf4f;
        src61 <= 12'h41d;
        src62 <= 12'hc50;
        src63 <= 12'hbe3;
        src64 <= 12'h399;
        src65 <= 12'h882;
        src66 <= 12'h3fb;
        src67 <= 12'hf2d;
        src68 <= 12'h6ea;
        src69 <= 12'he2b;
        src70 <= 12'h260;
        src71 <= 12'h88f;
        src72 <= 12'h3c7;
        src73 <= 12'hdd1;
        src74 <= 12'h6fe;
        src75 <= 12'h88;
        src76 <= 12'h6d9;
        src77 <= 12'h207;
        src78 <= 12'he65;
        src79 <= 12'hd66;
        src80 <= 12'h518;
        src81 <= 12'h872;
        src82 <= 12'h9df;
        src83 <= 12'hc12;
        src84 <= 12'h2f3;
        src85 <= 12'h222;
        src86 <= 12'h950;
        src87 <= 12'h8ad;
        src88 <= 12'he07;
        src89 <= 12'h7bc;
        src90 <= 12'h61f;
        src91 <= 12'hbac;
        src92 <= 12'h528;
        src93 <= 12'hc9f;
        src94 <= 12'he3d;
        src95 <= 12'h3d1;
        src96 <= 12'h31d;
        src97 <= 12'hf3b;
        src98 <= 12'h66a;
        src99 <= 12'h9a7;
        src100 <= 12'hbb2;
        src101 <= 12'h426;
        src102 <= 12'heff;
        src103 <= 12'h790;
        src104 <= 12'h160;
        src105 <= 12'h874;
        src106 <= 12'h120;
        src107 <= 12'h125;
        src108 <= 12'h554;
        src109 <= 12'hb00;
        src110 <= 12'hade;
        src111 <= 12'hcb3;
        src112 <= 12'hfdc;
        src113 <= 12'h8cc;
        src114 <= 12'h870;
        src115 <= 12'h1c8;
        src116 <= 12'h2ed;
        src117 <= 12'h976;
        src118 <= 12'hbd5;
        src119 <= 12'h67c;
        src120 <= 12'h3be;
        src121 <= 12'h6e0;
        src122 <= 12'hb2d;
        src123 <= 12'hc6d;
        src124 <= 12'h9c;
        src125 <= 12'hd23;
        src126 <= 12'hd17;
        src127 <= 12'hdc4;
        src128 <= 12'h379;
        src129 <= 12'hcaa;
        src130 <= 12'h2af;
        src131 <= 12'h390;
        src132 <= 12'h104;
        src133 <= 12'hc25;
        src134 <= 12'hcec;
        src135 <= 12'h826;
        src136 <= 12'h5a3;
        src137 <= 12'h39a;
        src138 <= 12'h6b;
        src139 <= 12'h7c4;
        src140 <= 12'h450;
        src141 <= 12'hcfa;
        src142 <= 12'hfe4;
        src143 <= 12'h5e7;
        src144 <= 12'h12f;
        src145 <= 12'haee;
        src146 <= 12'h100;
        src147 <= 12'h5bc;
        src148 <= 12'h76a;
        src149 <= 12'h802;
        src150 <= 12'h7d;
        src151 <= 12'hf05;
        src152 <= 12'hc17;
        src153 <= 12'h441;
        src154 <= 12'h179;
        src155 <= 12'h75d;
        src156 <= 12'h917;
        src157 <= 12'h1e0;
        src158 <= 12'h81b;
        src159 <= 12'h62a;
        src160 <= 12'hf05;
        src161 <= 12'ha73;
        exp <= 20'h50f13;
        #1
        src0 <= 12'hdbe;
        src1 <= 12'h101;
        src2 <= 12'hfee;
        src3 <= 12'h358;
        src4 <= 12'h5f9;
        src5 <= 12'ha0d;
        src6 <= 12'h85d;
        src7 <= 12'h616;
        src8 <= 12'h45;
        src9 <= 12'hf53;
        src10 <= 12'h6ca;
        src11 <= 12'hcb9;
        src12 <= 12'hff0;
        src13 <= 12'h456;
        src14 <= 12'hb30;
        src15 <= 12'h215;
        src16 <= 12'h390;
        src17 <= 12'hc1f;
        src18 <= 12'h866;
        src19 <= 12'h762;
        src20 <= 12'h9a5;
        src21 <= 12'h927;
        src22 <= 12'hab4;
        src23 <= 12'h30d;
        src24 <= 12'hc70;
        src25 <= 12'h12e;
        src26 <= 12'h106;
        src27 <= 12'h6b8;
        src28 <= 12'hbc3;
        src29 <= 12'h9ba;
        src30 <= 12'h3b5;
        src31 <= 12'hc53;
        src32 <= 12'hd88;
        src33 <= 12'hb67;
        src34 <= 12'h862;
        src35 <= 12'h563;
        src36 <= 12'h82d;
        src37 <= 12'hd4a;
        src38 <= 12'hd3c;
        src39 <= 12'h7c2;
        src40 <= 12'h74d;
        src41 <= 12'hd38;
        src42 <= 12'h2f;
        src43 <= 12'he47;
        src44 <= 12'h4a3;
        src45 <= 12'h470;
        src46 <= 12'hd1f;
        src47 <= 12'hc;
        src48 <= 12'h730;
        src49 <= 12'hd50;
        src50 <= 12'h49;
        src51 <= 12'h610;
        src52 <= 12'hd37;
        src53 <= 12'h97c;
        src54 <= 12'h637;
        src55 <= 12'hd86;
        src56 <= 12'hd04;
        src57 <= 12'h16c;
        src58 <= 12'h2c7;
        src59 <= 12'h278;
        src60 <= 12'h3e3;
        src61 <= 12'h52a;
        src62 <= 12'h4f2;
        src63 <= 12'hfa7;
        src64 <= 12'h948;
        src65 <= 12'he1a;
        src66 <= 12'h6ee;
        src67 <= 12'h873;
        src68 <= 12'h350;
        src69 <= 12'hf57;
        src70 <= 12'h7a0;
        src71 <= 12'hfd9;
        src72 <= 12'hc4d;
        src73 <= 12'h70a;
        src74 <= 12'h1a9;
        src75 <= 12'h52;
        src76 <= 12'h775;
        src77 <= 12'h5a7;
        src78 <= 12'hd08;
        src79 <= 12'h561;
        src80 <= 12'hea6;
        src81 <= 12'h57d;
        src82 <= 12'hdbc;
        src83 <= 12'h2f3;
        src84 <= 12'h654;
        src85 <= 12'hc5c;
        src86 <= 12'hce9;
        src87 <= 12'hc67;
        src88 <= 12'hee4;
        src89 <= 12'ha15;
        src90 <= 12'h239;
        src91 <= 12'h5d4;
        src92 <= 12'hfaf;
        src93 <= 12'h3e7;
        src94 <= 12'h45;
        src95 <= 12'hb7f;
        src96 <= 12'hcfc;
        src97 <= 12'hb26;
        src98 <= 12'h90;
        src99 <= 12'h4fe;
        src100 <= 12'h85b;
        src101 <= 12'hd08;
        src102 <= 12'h701;
        src103 <= 12'hf77;
        src104 <= 12'habe;
        src105 <= 12'h5b9;
        src106 <= 12'h67d;
        src107 <= 12'hd53;
        src108 <= 12'hb9d;
        src109 <= 12'he3f;
        src110 <= 12'h3df;
        src111 <= 12'hc56;
        src112 <= 12'hd28;
        src113 <= 12'hd43;
        src114 <= 12'h581;
        src115 <= 12'h9c0;
        src116 <= 12'hc1b;
        src117 <= 12'h92;
        src118 <= 12'hc0c;
        src119 <= 12'h5ae;
        src120 <= 12'ha77;
        src121 <= 12'h54f;
        src122 <= 12'h62e;
        src123 <= 12'hae0;
        src124 <= 12'ha4f;
        src125 <= 12'hd15;
        src126 <= 12'hcf9;
        src127 <= 12'h6ae;
        src128 <= 12'h4bf;
        src129 <= 12'h21a;
        src130 <= 12'ha9a;
        src131 <= 12'h974;
        src132 <= 12'hdaa;
        src133 <= 12'h388;
        src134 <= 12'h5cc;
        src135 <= 12'h146;
        src136 <= 12'h1ea;
        src137 <= 12'hbfc;
        src138 <= 12'hbfa;
        src139 <= 12'h6c5;
        src140 <= 12'h702;
        src141 <= 12'h678;
        src142 <= 12'h251;
        src143 <= 12'hd31;
        src144 <= 12'h43d;
        src145 <= 12'h56c;
        src146 <= 12'h822;
        src147 <= 12'hc4e;
        src148 <= 12'h849;
        src149 <= 12'ha46;
        src150 <= 12'h88d;
        src151 <= 12'he88;
        src152 <= 12'hf51;
        src153 <= 12'h5a0;
        src154 <= 12'h968;
        src155 <= 12'h476;
        src156 <= 12'h55b;
        src157 <= 12'hba8;
        src158 <= 12'h6e7;
        src159 <= 12'ha50;
        src160 <= 12'h5a5;
        src161 <= 12'hb84;
        exp <= 20'h55285;
        #1
        src0 <= 12'h33e;
        src1 <= 12'h86b;
        src2 <= 12'hb65;
        src3 <= 12'ha78;
        src4 <= 12'ha7a;
        src5 <= 12'h6a9;
        src6 <= 12'haab;
        src7 <= 12'hc95;
        src8 <= 12'hd42;
        src9 <= 12'h441;
        src10 <= 12'h6;
        src11 <= 12'h929;
        src12 <= 12'heed;
        src13 <= 12'h382;
        src14 <= 12'h7b8;
        src15 <= 12'h9fc;
        src16 <= 12'h9a5;
        src17 <= 12'h75d;
        src18 <= 12'h157;
        src19 <= 12'h79;
        src20 <= 12'h68b;
        src21 <= 12'hfac;
        src22 <= 12'h830;
        src23 <= 12'heb9;
        src24 <= 12'h8;
        src25 <= 12'h658;
        src26 <= 12'h105;
        src27 <= 12'hc26;
        src28 <= 12'h738;
        src29 <= 12'h133;
        src30 <= 12'h8e2;
        src31 <= 12'h42a;
        src32 <= 12'h582;
        src33 <= 12'h5d6;
        src34 <= 12'hf52;
        src35 <= 12'h48;
        src36 <= 12'h9f;
        src37 <= 12'h78f;
        src38 <= 12'h420;
        src39 <= 12'h454;
        src40 <= 12'hffa;
        src41 <= 12'h82c;
        src42 <= 12'hb8d;
        src43 <= 12'h839;
        src44 <= 12'hb3;
        src45 <= 12'h36e;
        src46 <= 12'h506;
        src47 <= 12'hda1;
        src48 <= 12'h927;
        src49 <= 12'ha7a;
        src50 <= 12'ha4;
        src51 <= 12'h826;
        src52 <= 12'h6d;
        src53 <= 12'h248;
        src54 <= 12'h182;
        src55 <= 12'h222;
        src56 <= 12'hd90;
        src57 <= 12'h8eb;
        src58 <= 12'h2fb;
        src59 <= 12'h48b;
        src60 <= 12'hd26;
        src61 <= 12'h8c8;
        src62 <= 12'h1e0;
        src63 <= 12'hd24;
        src64 <= 12'h1cb;
        src65 <= 12'hd69;
        src66 <= 12'hd51;
        src67 <= 12'ha6;
        src68 <= 12'h696;
        src69 <= 12'h3a3;
        src70 <= 12'hbe2;
        src71 <= 12'hbf7;
        src72 <= 12'hb9;
        src73 <= 12'hec6;
        src74 <= 12'he0f;
        src75 <= 12'hb63;
        src76 <= 12'h214;
        src77 <= 12'ha31;
        src78 <= 12'hb13;
        src79 <= 12'h5a5;
        src80 <= 12'ha43;
        src81 <= 12'he9;
        src82 <= 12'he42;
        src83 <= 12'h1d5;
        src84 <= 12'ha29;
        src85 <= 12'h7d8;
        src86 <= 12'hbf8;
        src87 <= 12'he4;
        src88 <= 12'h3c8;
        src89 <= 12'h15f;
        src90 <= 12'hdaf;
        src91 <= 12'h25f;
        src92 <= 12'hb9;
        src93 <= 12'h17f;
        src94 <= 12'hddd;
        src95 <= 12'h48f;
        src96 <= 12'hfbe;
        src97 <= 12'h4c9;
        src98 <= 12'h7b9;
        src99 <= 12'hcff;
        src100 <= 12'h8c3;
        src101 <= 12'h8f7;
        src102 <= 12'h492;
        src103 <= 12'h317;
        src104 <= 12'h584;
        src105 <= 12'hb7c;
        src106 <= 12'h643;
        src107 <= 12'hba2;
        src108 <= 12'h87a;
        src109 <= 12'h163;
        src110 <= 12'h519;
        src111 <= 12'h5a2;
        src112 <= 12'h74f;
        src113 <= 12'h866;
        src114 <= 12'h9b9;
        src115 <= 12'h72c;
        src116 <= 12'h103;
        src117 <= 12'hc71;
        src118 <= 12'ha76;
        src119 <= 12'h1a;
        src120 <= 12'h656;
        src121 <= 12'hd96;
        src122 <= 12'h88c;
        src123 <= 12'hd1f;
        src124 <= 12'hdae;
        src125 <= 12'hf1;
        src126 <= 12'hb98;
        src127 <= 12'hd5f;
        src128 <= 12'h4b5;
        src129 <= 12'h98c;
        src130 <= 12'h90a;
        src131 <= 12'he9d;
        src132 <= 12'he02;
        src133 <= 12'h24b;
        src134 <= 12'hef4;
        src135 <= 12'h3b9;
        src136 <= 12'h2d4;
        src137 <= 12'hf40;
        src138 <= 12'h274;
        src139 <= 12'he6b;
        src140 <= 12'hd5a;
        src141 <= 12'hda2;
        src142 <= 12'h422;
        src143 <= 12'h676;
        src144 <= 12'hcac;
        src145 <= 12'h6cb;
        src146 <= 12'h942;
        src147 <= 12'h5c7;
        src148 <= 12'h8eb;
        src149 <= 12'h1a2;
        src150 <= 12'h396;
        src151 <= 12'h6a0;
        src152 <= 12'h266;
        src153 <= 12'he16;
        src154 <= 12'hed1;
        src155 <= 12'hf51;
        src156 <= 12'hd3;
        src157 <= 12'h364;
        src158 <= 12'h11d;
        src159 <= 12'h23a;
        src160 <= 12'hfab;
        src161 <= 12'heb9;
        exp <= 20'h4cffb;
        #1
        src0 <= 12'h540;
        src1 <= 12'h9d2;
        src2 <= 12'ha9b;
        src3 <= 12'h73c;
        src4 <= 12'h581;
        src5 <= 12'h529;
        src6 <= 12'hc2e;
        src7 <= 12'ha9c;
        src8 <= 12'hcac;
        src9 <= 12'haf8;
        src10 <= 12'h33e;
        src11 <= 12'h426;
        src12 <= 12'h257;
        src13 <= 12'hb03;
        src14 <= 12'ha6a;
        src15 <= 12'hf49;
        src16 <= 12'hce3;
        src17 <= 12'hde;
        src18 <= 12'h358;
        src19 <= 12'ha93;
        src20 <= 12'h18d;
        src21 <= 12'hb7d;
        src22 <= 12'h56b;
        src23 <= 12'ha98;
        src24 <= 12'h47f;
        src25 <= 12'hc57;
        src26 <= 12'h51f;
        src27 <= 12'h145;
        src28 <= 12'h2d9;
        src29 <= 12'h639;
        src30 <= 12'h7eb;
        src31 <= 12'h52f;
        src32 <= 12'h700;
        src33 <= 12'hb04;
        src34 <= 12'h49f;
        src35 <= 12'h6e6;
        src36 <= 12'h4af;
        src37 <= 12'h215;
        src38 <= 12'h966;
        src39 <= 12'he9b;
        src40 <= 12'h26b;
        src41 <= 12'ha23;
        src42 <= 12'he74;
        src43 <= 12'h278;
        src44 <= 12'h761;
        src45 <= 12'h687;
        src46 <= 12'h100;
        src47 <= 12'h8bb;
        src48 <= 12'hc9a;
        src49 <= 12'h63;
        src50 <= 12'hee6;
        src51 <= 12'h3d6;
        src52 <= 12'hff8;
        src53 <= 12'h83f;
        src54 <= 12'h80f;
        src55 <= 12'hef1;
        src56 <= 12'he14;
        src57 <= 12'hed2;
        src58 <= 12'h124;
        src59 <= 12'h1d7;
        src60 <= 12'h20b;
        src61 <= 12'h415;
        src62 <= 12'hdca;
        src63 <= 12'h8ef;
        src64 <= 12'h65d;
        src65 <= 12'ha18;
        src66 <= 12'h4cf;
        src67 <= 12'hd27;
        src68 <= 12'h234;
        src69 <= 12'h708;
        src70 <= 12'hdf4;
        src71 <= 12'h515;
        src72 <= 12'h434;
        src73 <= 12'h2be;
        src74 <= 12'hd18;
        src75 <= 12'hcb3;
        src76 <= 12'h5ba;
        src77 <= 12'h3af;
        src78 <= 12'hb55;
        src79 <= 12'h7a4;
        src80 <= 12'h9ef;
        src81 <= 12'h9bf;
        src82 <= 12'h212;
        src83 <= 12'h858;
        src84 <= 12'h7a;
        src85 <= 12'had4;
        src86 <= 12'he46;
        src87 <= 12'hb2f;
        src88 <= 12'h704;
        src89 <= 12'h8f6;
        src90 <= 12'h83d;
        src91 <= 12'hb17;
        src92 <= 12'h688;
        src93 <= 12'h2c8;
        src94 <= 12'h6ba;
        src95 <= 12'h860;
        src96 <= 12'h7d8;
        src97 <= 12'h782;
        src98 <= 12'h63;
        src99 <= 12'h9d8;
        src100 <= 12'h198;
        src101 <= 12'h5b8;
        src102 <= 12'h687;
        src103 <= 12'hd40;
        src104 <= 12'h1f0;
        src105 <= 12'hdc1;
        src106 <= 12'h1be;
        src107 <= 12'hc4b;
        src108 <= 12'h1c6;
        src109 <= 12'h61;
        src110 <= 12'ha18;
        src111 <= 12'hd65;
        src112 <= 12'hee8;
        src113 <= 12'h2c6;
        src114 <= 12'h240;
        src115 <= 12'hbb1;
        src116 <= 12'h98d;
        src117 <= 12'h134;
        src118 <= 12'hcd9;
        src119 <= 12'h6d5;
        src120 <= 12'hc36;
        src121 <= 12'hac5;
        src122 <= 12'h4b7;
        src123 <= 12'he81;
        src124 <= 12'h4df;
        src125 <= 12'h21f;
        src126 <= 12'hee2;
        src127 <= 12'h1c2;
        src128 <= 12'h8f3;
        src129 <= 12'hedb;
        src130 <= 12'h70e;
        src131 <= 12'h5be;
        src132 <= 12'h1a;
        src133 <= 12'hedd;
        src134 <= 12'hee7;
        src135 <= 12'h2;
        src136 <= 12'h7e3;
        src137 <= 12'h39f;
        src138 <= 12'h610;
        src139 <= 12'h6a8;
        src140 <= 12'h5a;
        src141 <= 12'hc93;
        src142 <= 12'h483;
        src143 <= 12'h8dd;
        src144 <= 12'h78d;
        src145 <= 12'haaf;
        src146 <= 12'h178;
        src147 <= 12'h480;
        src148 <= 12'h39f;
        src149 <= 12'h638;
        src150 <= 12'h594;
        src151 <= 12'hd2b;
        src152 <= 12'h785;
        src153 <= 12'h490;
        src154 <= 12'hfdc;
        src155 <= 12'h92a;
        src156 <= 12'h514;
        src157 <= 12'h881;
        src158 <= 12'h90e;
        src159 <= 12'hd2d;
        src160 <= 12'h8a1;
        src161 <= 12'h3b5;
        exp <= 20'h4d101;
        #1
        src0 <= 12'hd12;
        src1 <= 12'hcfb;
        src2 <= 12'hfb8;
        src3 <= 12'h70a;
        src4 <= 12'h8f7;
        src5 <= 12'h9e1;
        src6 <= 12'h379;
        src7 <= 12'h369;
        src8 <= 12'h38;
        src9 <= 12'h335;
        src10 <= 12'h3d2;
        src11 <= 12'h838;
        src12 <= 12'h485;
        src13 <= 12'h6bb;
        src14 <= 12'haa4;
        src15 <= 12'h33b;
        src16 <= 12'ha38;
        src17 <= 12'h57;
        src18 <= 12'h1b2;
        src19 <= 12'hec3;
        src20 <= 12'hb10;
        src21 <= 12'h907;
        src22 <= 12'h98f;
        src23 <= 12'h325;
        src24 <= 12'h127;
        src25 <= 12'h8bc;
        src26 <= 12'hab;
        src27 <= 12'he2f;
        src28 <= 12'h77e;
        src29 <= 12'h40b;
        src30 <= 12'hdcf;
        src31 <= 12'hb6b;
        src32 <= 12'h457;
        src33 <= 12'h43d;
        src34 <= 12'h587;
        src35 <= 12'he22;
        src36 <= 12'hf3b;
        src37 <= 12'h807;
        src38 <= 12'h66f;
        src39 <= 12'h824;
        src40 <= 12'hcca;
        src41 <= 12'h101;
        src42 <= 12'hb45;
        src43 <= 12'h556;
        src44 <= 12'h7eb;
        src45 <= 12'hf32;
        src46 <= 12'ha9e;
        src47 <= 12'h2e8;
        src48 <= 12'hd14;
        src49 <= 12'h721;
        src50 <= 12'h5f5;
        src51 <= 12'ha58;
        src52 <= 12'h93d;
        src53 <= 12'h51;
        src54 <= 12'h76f;
        src55 <= 12'hd7c;
        src56 <= 12'h56e;
        src57 <= 12'h22c;
        src58 <= 12'h50b;
        src59 <= 12'h52b;
        src60 <= 12'h89b;
        src61 <= 12'ha98;
        src62 <= 12'h6f6;
        src63 <= 12'h3d9;
        src64 <= 12'h8a6;
        src65 <= 12'hda8;
        src66 <= 12'hdfc;
        src67 <= 12'hc2;
        src68 <= 12'hb62;
        src69 <= 12'h77c;
        src70 <= 12'hc4b;
        src71 <= 12'h79a;
        src72 <= 12'h1ce;
        src73 <= 12'h18d;
        src74 <= 12'hdd5;
        src75 <= 12'h20e;
        src76 <= 12'hfd1;
        src77 <= 12'hcb7;
        src78 <= 12'h1b4;
        src79 <= 12'hdca;
        src80 <= 12'h261;
        src81 <= 12'h54e;
        src82 <= 12'h44f;
        src83 <= 12'hc29;
        src84 <= 12'hc32;
        src85 <= 12'hd26;
        src86 <= 12'h91e;
        src87 <= 12'hffc;
        src88 <= 12'h140;
        src89 <= 12'hdd8;
        src90 <= 12'h45c;
        src91 <= 12'hbaf;
        src92 <= 12'hfdf;
        src93 <= 12'hd56;
        src94 <= 12'hf5;
        src95 <= 12'h946;
        src96 <= 12'h547;
        src97 <= 12'h894;
        src98 <= 12'hd6e;
        src99 <= 12'hc11;
        src100 <= 12'h4f;
        src101 <= 12'h859;
        src102 <= 12'ha08;
        src103 <= 12'h94e;
        src104 <= 12'hc6d;
        src105 <= 12'hc73;
        src106 <= 12'hb3a;
        src107 <= 12'h37b;
        src108 <= 12'hc10;
        src109 <= 12'h299;
        src110 <= 12'heac;
        src111 <= 12'h492;
        src112 <= 12'h6af;
        src113 <= 12'h78e;
        src114 <= 12'ha50;
        src115 <= 12'hee0;
        src116 <= 12'ha1d;
        src117 <= 12'h496;
        src118 <= 12'h4cc;
        src119 <= 12'h7e0;
        src120 <= 12'hedc;
        src121 <= 12'hb6b;
        src122 <= 12'h26f;
        src123 <= 12'hbbe;
        src124 <= 12'h741;
        src125 <= 12'hcc0;
        src126 <= 12'h835;
        src127 <= 12'h94c;
        src128 <= 12'h60a;
        src129 <= 12'hf9c;
        src130 <= 12'h8f7;
        src131 <= 12'h665;
        src132 <= 12'h9f6;
        src133 <= 12'h960;
        src134 <= 12'h9f8;
        src135 <= 12'h38d;
        src136 <= 12'hec6;
        src137 <= 12'h482;
        src138 <= 12'h814;
        src139 <= 12'h8b5;
        src140 <= 12'h2fa;
        src141 <= 12'h6f;
        src142 <= 12'h894;
        src143 <= 12'h120;
        src144 <= 12'h2d0;
        src145 <= 12'he9f;
        src146 <= 12'h5cf;
        src147 <= 12'hc37;
        src148 <= 12'h8b7;
        src149 <= 12'h71b;
        src150 <= 12'h9aa;
        src151 <= 12'h297;
        src152 <= 12'hb3e;
        src153 <= 12'h25e;
        src154 <= 12'hba5;
        src155 <= 12'h47;
        src156 <= 12'h3ac;
        src157 <= 12'h870;
        src158 <= 12'h408;
        src159 <= 12'hf9c;
        src160 <= 12'h57;
        src161 <= 12'h195;
        exp <= 20'h50ff2;
        #1
        src0 <= 12'hf6f;
        src1 <= 12'h57b;
        src2 <= 12'hb17;
        src3 <= 12'h5b9;
        src4 <= 12'h1da;
        src5 <= 12'h74f;
        src6 <= 12'hab4;
        src7 <= 12'hc76;
        src8 <= 12'hb43;
        src9 <= 12'h2ad;
        src10 <= 12'hcb4;
        src11 <= 12'h710;
        src12 <= 12'h77;
        src13 <= 12'h9d0;
        src14 <= 12'hbbf;
        src15 <= 12'hd8d;
        src16 <= 12'h7c6;
        src17 <= 12'h1af;
        src18 <= 12'h43e;
        src19 <= 12'hdd;
        src20 <= 12'hefe;
        src21 <= 12'haf6;
        src22 <= 12'h406;
        src23 <= 12'hb8c;
        src24 <= 12'h3c9;
        src25 <= 12'h342;
        src26 <= 12'h865;
        src27 <= 12'h90f;
        src28 <= 12'h634;
        src29 <= 12'h256;
        src30 <= 12'h26b;
        src31 <= 12'ha8a;
        src32 <= 12'h310;
        src33 <= 12'hb1f;
        src34 <= 12'h313;
        src35 <= 12'hc;
        src36 <= 12'h3c4;
        src37 <= 12'hca8;
        src38 <= 12'h520;
        src39 <= 12'hbc7;
        src40 <= 12'hdbd;
        src41 <= 12'h1e5;
        src42 <= 12'hf73;
        src43 <= 12'hb59;
        src44 <= 12'he88;
        src45 <= 12'he7b;
        src46 <= 12'h215;
        src47 <= 12'heae;
        src48 <= 12'h71c;
        src49 <= 12'hee2;
        src50 <= 12'ha2c;
        src51 <= 12'h342;
        src52 <= 12'h44e;
        src53 <= 12'hc36;
        src54 <= 12'hd1b;
        src55 <= 12'h997;
        src56 <= 12'h1cb;
        src57 <= 12'h25c;
        src58 <= 12'h614;
        src59 <= 12'h794;
        src60 <= 12'hb3d;
        src61 <= 12'hc6a;
        src62 <= 12'h643;
        src63 <= 12'h184;
        src64 <= 12'h621;
        src65 <= 12'hf25;
        src66 <= 12'h476;
        src67 <= 12'ha65;
        src68 <= 12'h362;
        src69 <= 12'h55e;
        src70 <= 12'hf01;
        src71 <= 12'h9e6;
        src72 <= 12'h416;
        src73 <= 12'h58d;
        src74 <= 12'h35f;
        src75 <= 12'hea0;
        src76 <= 12'hbd1;
        src77 <= 12'h3d3;
        src78 <= 12'hd0b;
        src79 <= 12'h47;
        src80 <= 12'h7f7;
        src81 <= 12'h7e0;
        src82 <= 12'h9c8;
        src83 <= 12'h687;
        src84 <= 12'hb9f;
        src85 <= 12'h8da;
        src86 <= 12'hce7;
        src87 <= 12'he01;
        src88 <= 12'he64;
        src89 <= 12'h670;
        src90 <= 12'h468;
        src91 <= 12'hb82;
        src92 <= 12'hd76;
        src93 <= 12'h6f;
        src94 <= 12'hab0;
        src95 <= 12'heac;
        src96 <= 12'ha30;
        src97 <= 12'h384;
        src98 <= 12'ha5;
        src99 <= 12'hfdb;
        src100 <= 12'h3c0;
        src101 <= 12'h4ae;
        src102 <= 12'h4f;
        src103 <= 12'hb13;
        src104 <= 12'h864;
        src105 <= 12'h828;
        src106 <= 12'hf33;
        src107 <= 12'hc0a;
        src108 <= 12'h56d;
        src109 <= 12'h85c;
        src110 <= 12'h47d;
        src111 <= 12'h630;
        src112 <= 12'h6cf;
        src113 <= 12'hce2;
        src114 <= 12'h41f;
        src115 <= 12'h6f0;
        src116 <= 12'h8d8;
        src117 <= 12'h702;
        src118 <= 12'h679;
        src119 <= 12'h32;
        src120 <= 12'h777;
        src121 <= 12'h4fc;
        src122 <= 12'hba9;
        src123 <= 12'hdf9;
        src124 <= 12'hb1a;
        src125 <= 12'ha93;
        src126 <= 12'hb08;
        src127 <= 12'h9df;
        src128 <= 12'h66b;
        src129 <= 12'hce3;
        src130 <= 12'hd9b;
        src131 <= 12'h408;
        src132 <= 12'h2cf;
        src133 <= 12'h889;
        src134 <= 12'hc47;
        src135 <= 12'h6b0;
        src136 <= 12'h88c;
        src137 <= 12'hd8c;
        src138 <= 12'h341;
        src139 <= 12'h650;
        src140 <= 12'h990;
        src141 <= 12'hf8a;
        src142 <= 12'h7f8;
        src143 <= 12'he05;
        src144 <= 12'h50d;
        src145 <= 12'h684;
        src146 <= 12'h295;
        src147 <= 12'h1f6;
        src148 <= 12'hed8;
        src149 <= 12'h32d;
        src150 <= 12'h32;
        src151 <= 12'h8d4;
        src152 <= 12'hc47;
        src153 <= 12'h597;
        src154 <= 12'hf95;
        src155 <= 12'h727;
        src156 <= 12'h29a;
        src157 <= 12'he46;
        src158 <= 12'hb8e;
        src159 <= 12'h534;
        src160 <= 12'hb8b;
        src161 <= 12'h2d2;
        exp <= 20'h523f3;
        #1
        src0 <= 12'he85;
        src1 <= 12'hc0d;
        src2 <= 12'h83c;
        src3 <= 12'he9e;
        src4 <= 12'h461;
        src5 <= 12'h98f;
        src6 <= 12'h32d;
        src7 <= 12'h1ee;
        src8 <= 12'hfa;
        src9 <= 12'h12a;
        src10 <= 12'h1c5;
        src11 <= 12'h425;
        src12 <= 12'h98d;
        src13 <= 12'he52;
        src14 <= 12'hf75;
        src15 <= 12'hb5;
        src16 <= 12'hbaa;
        src17 <= 12'hfae;
        src18 <= 12'h20d;
        src19 <= 12'he72;
        src20 <= 12'hde8;
        src21 <= 12'h1f4;
        src22 <= 12'h517;
        src23 <= 12'h3d4;
        src24 <= 12'h9e6;
        src25 <= 12'hb52;
        src26 <= 12'h5c;
        src27 <= 12'h394;
        src28 <= 12'h7b9;
        src29 <= 12'h7b4;
        src30 <= 12'hca5;
        src31 <= 12'he4;
        src32 <= 12'h7a8;
        src33 <= 12'ha1b;
        src34 <= 12'h6b6;
        src35 <= 12'h6b6;
        src36 <= 12'head;
        src37 <= 12'hf34;
        src38 <= 12'hdcc;
        src39 <= 12'hf9d;
        src40 <= 12'h583;
        src41 <= 12'h5ae;
        src42 <= 12'ha7b;
        src43 <= 12'hdc7;
        src44 <= 12'h3aa;
        src45 <= 12'hc1c;
        src46 <= 12'h47e;
        src47 <= 12'h968;
        src48 <= 12'hf65;
        src49 <= 12'hee2;
        src50 <= 12'h574;
        src51 <= 12'hc23;
        src52 <= 12'h372;
        src53 <= 12'hc0d;
        src54 <= 12'h7fa;
        src55 <= 12'hfdc;
        src56 <= 12'he19;
        src57 <= 12'hca9;
        src58 <= 12'h1b3;
        src59 <= 12'hd40;
        src60 <= 12'h3d1;
        src61 <= 12'hafb;
        src62 <= 12'h12b;
        src63 <= 12'h8c;
        src64 <= 12'h9d5;
        src65 <= 12'hcaa;
        src66 <= 12'h48;
        src67 <= 12'hc75;
        src68 <= 12'h712;
        src69 <= 12'h25f;
        src70 <= 12'h1c7;
        src71 <= 12'hf42;
        src72 <= 12'h88f;
        src73 <= 12'h959;
        src74 <= 12'he1a;
        src75 <= 12'hf6b;
        src76 <= 12'h1bf;
        src77 <= 12'h69b;
        src78 <= 12'hf08;
        src79 <= 12'h5f5;
        src80 <= 12'hb7d;
        src81 <= 12'he8a;
        src82 <= 12'h630;
        src83 <= 12'hb03;
        src84 <= 12'hf58;
        src85 <= 12'h8ae;
        src86 <= 12'he20;
        src87 <= 12'h3b4;
        src88 <= 12'hf47;
        src89 <= 12'h712;
        src90 <= 12'h1c9;
        src91 <= 12'h996;
        src92 <= 12'h42f;
        src93 <= 12'h719;
        src94 <= 12'h387;
        src95 <= 12'h969;
        src96 <= 12'hbc1;
        src97 <= 12'hbc1;
        src98 <= 12'hb43;
        src99 <= 12'hf9e;
        src100 <= 12'h369;
        src101 <= 12'hfb8;
        src102 <= 12'h470;
        src103 <= 12'he23;
        src104 <= 12'h218;
        src105 <= 12'h382;
        src106 <= 12'ha9a;
        src107 <= 12'he9;
        src108 <= 12'ha2;
        src109 <= 12'h713;
        src110 <= 12'h706;
        src111 <= 12'hee8;
        src112 <= 12'h8b4;
        src113 <= 12'h285;
        src114 <= 12'h132;
        src115 <= 12'h190;
        src116 <= 12'h152;
        src117 <= 12'h536;
        src118 <= 12'hfff;
        src119 <= 12'h741;
        src120 <= 12'he7f;
        src121 <= 12'h1b5;
        src122 <= 12'he6a;
        src123 <= 12'hf8c;
        src124 <= 12'ha5d;
        src125 <= 12'h5be;
        src126 <= 12'h309;
        src127 <= 12'hc1e;
        src128 <= 12'h3fb;
        src129 <= 12'hd08;
        src130 <= 12'hc12;
        src131 <= 12'h958;
        src132 <= 12'h593;
        src133 <= 12'h74a;
        src134 <= 12'hbb6;
        src135 <= 12'h9d9;
        src136 <= 12'h251;
        src137 <= 12'h219;
        src138 <= 12'h181;
        src139 <= 12'h610;
        src140 <= 12'hf16;
        src141 <= 12'h669;
        src142 <= 12'h3ae;
        src143 <= 12'he;
        src144 <= 12'hf0;
        src145 <= 12'he49;
        src146 <= 12'h663;
        src147 <= 12'h49e;
        src148 <= 12'hc8d;
        src149 <= 12'h87c;
        src150 <= 12'h44b;
        src151 <= 12'hdc9;
        src152 <= 12'h635;
        src153 <= 12'hbb8;
        src154 <= 12'h9b1;
        src155 <= 12'hec7;
        src156 <= 12'h39e;
        src157 <= 12'hf53;
        src158 <= 12'h9d1;
        src159 <= 12'h50d;
        src160 <= 12'h389;
        src161 <= 12'h42e;
        exp <= 20'h53922;
        #1
        src0 <= 12'h3c8;
        src1 <= 12'ha52;
        src2 <= 12'h8b9;
        src3 <= 12'h442;
        src4 <= 12'hf95;
        src5 <= 12'h64b;
        src6 <= 12'h7c0;
        src7 <= 12'h947;
        src8 <= 12'h63e;
        src9 <= 12'hec;
        src10 <= 12'hfdd;
        src11 <= 12'h9c6;
        src12 <= 12'h22;
        src13 <= 12'h4e1;
        src14 <= 12'hdcb;
        src15 <= 12'hdca;
        src16 <= 12'hd76;
        src17 <= 12'h4a2;
        src18 <= 12'hf37;
        src19 <= 12'hce4;
        src20 <= 12'ha02;
        src21 <= 12'h156;
        src22 <= 12'hb6a;
        src23 <= 12'he3f;
        src24 <= 12'hb0b;
        src25 <= 12'hbee;
        src26 <= 12'h749;
        src27 <= 12'hb87;
        src28 <= 12'ha0a;
        src29 <= 12'h4df;
        src30 <= 12'h176;
        src31 <= 12'h395;
        src32 <= 12'h568;
        src33 <= 12'h416;
        src34 <= 12'h4cd;
        src35 <= 12'h4b8;
        src36 <= 12'h6fd;
        src37 <= 12'hf3e;
        src38 <= 12'hecf;
        src39 <= 12'h594;
        src40 <= 12'h30b;
        src41 <= 12'h5a9;
        src42 <= 12'hc04;
        src43 <= 12'h88a;
        src44 <= 12'h52a;
        src45 <= 12'hcbc;
        src46 <= 12'h4fb;
        src47 <= 12'hf62;
        src48 <= 12'hc75;
        src49 <= 12'h5bc;
        src50 <= 12'ha37;
        src51 <= 12'h8e6;
        src52 <= 12'hf17;
        src53 <= 12'h500;
        src54 <= 12'h68e;
        src55 <= 12'hcb;
        src56 <= 12'h8db;
        src57 <= 12'hdfa;
        src58 <= 12'h8d0;
        src59 <= 12'h3a;
        src60 <= 12'hecf;
        src61 <= 12'ha92;
        src62 <= 12'hbd8;
        src63 <= 12'h351;
        src64 <= 12'h7d9;
        src65 <= 12'hc49;
        src66 <= 12'h921;
        src67 <= 12'h47e;
        src68 <= 12'h789;
        src69 <= 12'hec2;
        src70 <= 12'hec;
        src71 <= 12'hbab;
        src72 <= 12'h53f;
        src73 <= 12'hb9f;
        src74 <= 12'hee8;
        src75 <= 12'h12;
        src76 <= 12'h46e;
        src77 <= 12'h82a;
        src78 <= 12'h71a;
        src79 <= 12'h838;
        src80 <= 12'h4de;
        src81 <= 12'h4da;
        src82 <= 12'h946;
        src83 <= 12'h3f6;
        src84 <= 12'hfab;
        src85 <= 12'h5a8;
        src86 <= 12'hc80;
        src87 <= 12'h815;
        src88 <= 12'h22f;
        src89 <= 12'h167;
        src90 <= 12'hc12;
        src91 <= 12'h1a6;
        src92 <= 12'h361;
        src93 <= 12'hbd3;
        src94 <= 12'h770;
        src95 <= 12'h20a;
        src96 <= 12'h8a;
        src97 <= 12'h6ac;
        src98 <= 12'h27;
        src99 <= 12'h73;
        src100 <= 12'ha7d;
        src101 <= 12'h5f8;
        src102 <= 12'h2f1;
        src103 <= 12'h9cc;
        src104 <= 12'h71a;
        src105 <= 12'hf37;
        src106 <= 12'hb35;
        src107 <= 12'ha6f;
        src108 <= 12'h4ef;
        src109 <= 12'hbad;
        src110 <= 12'hd2d;
        src111 <= 12'h5ff;
        src112 <= 12'hd90;
        src113 <= 12'hd80;
        src114 <= 12'h365;
        src115 <= 12'h69b;
        src116 <= 12'h5ae;
        src117 <= 12'ha5;
        src118 <= 12'h521;
        src119 <= 12'hcfe;
        src120 <= 12'h125;
        src121 <= 12'hb1f;
        src122 <= 12'h41f;
        src123 <= 12'h3ca;
        src124 <= 12'h5c7;
        src125 <= 12'hcd1;
        src126 <= 12'he1c;
        src127 <= 12'ha52;
        src128 <= 12'h17d;
        src129 <= 12'h816;
        src130 <= 12'hac5;
        src131 <= 12'hc4f;
        src132 <= 12'h726;
        src133 <= 12'ha84;
        src134 <= 12'hd6a;
        src135 <= 12'h3ea;
        src136 <= 12'hefb;
        src137 <= 12'hf74;
        src138 <= 12'hf81;
        src139 <= 12'h771;
        src140 <= 12'h742;
        src141 <= 12'hf79;
        src142 <= 12'h7ba;
        src143 <= 12'h90e;
        src144 <= 12'h293;
        src145 <= 12'hf4a;
        src146 <= 12'hd84;
        src147 <= 12'hdc8;
        src148 <= 12'h502;
        src149 <= 12'h49b;
        src150 <= 12'hcfa;
        src151 <= 12'he22;
        src152 <= 12'h441;
        src153 <= 12'h397;
        src154 <= 12'haf3;
        src155 <= 12'h38a;
        src156 <= 12'h11e;
        src157 <= 12'hed2;
        src158 <= 12'h953;
        src159 <= 12'h8ae;
        src160 <= 12'hfc0;
        src161 <= 12'h479;
        exp <= 20'h53a3a;
        #1
        src0 <= 12'hc02;
        src1 <= 12'h9f;
        src2 <= 12'he3;
        src3 <= 12'hbe9;
        src4 <= 12'ha2f;
        src5 <= 12'h73f;
        src6 <= 12'hadd;
        src7 <= 12'h9d6;
        src8 <= 12'h796;
        src9 <= 12'h8ba;
        src10 <= 12'ha38;
        src11 <= 12'hace;
        src12 <= 12'h1cd;
        src13 <= 12'h700;
        src14 <= 12'he7;
        src15 <= 12'h3de;
        src16 <= 12'h2ff;
        src17 <= 12'h90b;
        src18 <= 12'h41e;
        src19 <= 12'hfb2;
        src20 <= 12'h40;
        src21 <= 12'hf8;
        src22 <= 12'h71b;
        src23 <= 12'h2c3;
        src24 <= 12'hd72;
        src25 <= 12'h6e0;
        src26 <= 12'h9d;
        src27 <= 12'h89b;
        src28 <= 12'he8;
        src29 <= 12'hf97;
        src30 <= 12'hcec;
        src31 <= 12'h885;
        src32 <= 12'h94;
        src33 <= 12'hb06;
        src34 <= 12'h349;
        src35 <= 12'h936;
        src36 <= 12'h432;
        src37 <= 12'hc1;
        src38 <= 12'h6f9;
        src39 <= 12'h22;
        src40 <= 12'h89b;
        src41 <= 12'h82;
        src42 <= 12'hdfd;
        src43 <= 12'h8b6;
        src44 <= 12'h572;
        src45 <= 12'h382;
        src46 <= 12'h26;
        src47 <= 12'h20f;
        src48 <= 12'h77b;
        src49 <= 12'h39e;
        src50 <= 12'h45f;
        src51 <= 12'hbf;
        src52 <= 12'hb2f;
        src53 <= 12'habe;
        src54 <= 12'he36;
        src55 <= 12'h7b;
        src56 <= 12'h8f4;
        src57 <= 12'h369;
        src58 <= 12'h364;
        src59 <= 12'hd72;
        src60 <= 12'he1;
        src61 <= 12'hf68;
        src62 <= 12'hac9;
        src63 <= 12'h99e;
        src64 <= 12'h271;
        src65 <= 12'h5a0;
        src66 <= 12'h2cf;
        src67 <= 12'hadc;
        src68 <= 12'hbf0;
        src69 <= 12'hb80;
        src70 <= 12'h8f3;
        src71 <= 12'h5a4;
        src72 <= 12'he7a;
        src73 <= 12'hd28;
        src74 <= 12'h4cc;
        src75 <= 12'he6f;
        src76 <= 12'hb04;
        src77 <= 12'h840;
        src78 <= 12'ha2;
        src79 <= 12'h603;
        src80 <= 12'h21e;
        src81 <= 12'hf76;
        src82 <= 12'hd4a;
        src83 <= 12'h2d;
        src84 <= 12'he4;
        src85 <= 12'h7a6;
        src86 <= 12'hbbf;
        src87 <= 12'h55;
        src88 <= 12'h598;
        src89 <= 12'ha7d;
        src90 <= 12'hefc;
        src91 <= 12'h7b4;
        src92 <= 12'h477;
        src93 <= 12'h1b8;
        src94 <= 12'h43c;
        src95 <= 12'h3b2;
        src96 <= 12'he6d;
        src97 <= 12'hd7b;
        src98 <= 12'h9b0;
        src99 <= 12'hff0;
        src100 <= 12'h62;
        src101 <= 12'h5ee;
        src102 <= 12'hf38;
        src103 <= 12'he3e;
        src104 <= 12'h1d2;
        src105 <= 12'h616;
        src106 <= 12'hf7d;
        src107 <= 12'h90f;
        src108 <= 12'h363;
        src109 <= 12'h9ee;
        src110 <= 12'h14d;
        src111 <= 12'h573;
        src112 <= 12'ha29;
        src113 <= 12'h7df;
        src114 <= 12'h665;
        src115 <= 12'h7bb;
        src116 <= 12'hf41;
        src117 <= 12'hc23;
        src118 <= 12'habc;
        src119 <= 12'hca8;
        src120 <= 12'hd7a;
        src121 <= 12'h85d;
        src122 <= 12'h821;
        src123 <= 12'hcd6;
        src124 <= 12'h8b;
        src125 <= 12'hf5c;
        src126 <= 12'he9b;
        src127 <= 12'haf8;
        src128 <= 12'hecd;
        src129 <= 12'hc03;
        src130 <= 12'h6b2;
        src131 <= 12'ha2b;
        src132 <= 12'h92f;
        src133 <= 12'h408;
        src134 <= 12'hdc7;
        src135 <= 12'h475;
        src136 <= 12'h81f;
        src137 <= 12'hd23;
        src138 <= 12'he6c;
        src139 <= 12'hd00;
        src140 <= 12'h5c9;
        src141 <= 12'hcc;
        src142 <= 12'hf86;
        src143 <= 12'ha36;
        src144 <= 12'hb0c;
        src145 <= 12'h9a3;
        src146 <= 12'h7f9;
        src147 <= 12'h573;
        src148 <= 12'h978;
        src149 <= 12'heb7;
        src150 <= 12'h5ac;
        src151 <= 12'hfab;
        src152 <= 12'h515;
        src153 <= 12'h73f;
        src154 <= 12'ha6f;
        src155 <= 12'hc2a;
        src156 <= 12'hb46;
        src157 <= 12'hae9;
        src158 <= 12'he51;
        src159 <= 12'hb5b;
        src160 <= 12'hd3e;
        src161 <= 12'h658;
        exp <= 20'h51af5;
        #1
        src0 <= 12'h54f;
        src1 <= 12'h341;
        src2 <= 12'hef2;
        src3 <= 12'hcfa;
        src4 <= 12'he0a;
        src5 <= 12'h6bd;
        src6 <= 12'hb28;
        src7 <= 12'h513;
        src8 <= 12'h9fa;
        src9 <= 12'h46e;
        src10 <= 12'h8d2;
        src11 <= 12'h903;
        src12 <= 12'h20e;
        src13 <= 12'hde1;
        src14 <= 12'hfb4;
        src15 <= 12'ha3f;
        src16 <= 12'hfe6;
        src17 <= 12'h57;
        src18 <= 12'hf0c;
        src19 <= 12'hc12;
        src20 <= 12'hc84;
        src21 <= 12'hbc1;
        src22 <= 12'hcb3;
        src23 <= 12'h1ad;
        src24 <= 12'h60d;
        src25 <= 12'hbb1;
        src26 <= 12'h90;
        src27 <= 12'hf72;
        src28 <= 12'h6b9;
        src29 <= 12'hac7;
        src30 <= 12'hff7;
        src31 <= 12'h66e;
        src32 <= 12'h201;
        src33 <= 12'hcd4;
        src34 <= 12'h7f1;
        src35 <= 12'hef2;
        src36 <= 12'hc1a;
        src37 <= 12'h991;
        src38 <= 12'h281;
        src39 <= 12'hc20;
        src40 <= 12'hdcd;
        src41 <= 12'hd89;
        src42 <= 12'ha09;
        src43 <= 12'hc0f;
        src44 <= 12'hdd2;
        src45 <= 12'h887;
        src46 <= 12'h119;
        src47 <= 12'hfe3;
        src48 <= 12'h3e8;
        src49 <= 12'h57f;
        src50 <= 12'h2c9;
        src51 <= 12'h9f4;
        src52 <= 12'h2da;
        src53 <= 12'hec;
        src54 <= 12'h81d;
        src55 <= 12'h8f8;
        src56 <= 12'h361;
        src57 <= 12'h6b5;
        src58 <= 12'he71;
        src59 <= 12'h2f0;
        src60 <= 12'heb2;
        src61 <= 12'he68;
        src62 <= 12'h5fb;
        src63 <= 12'h1cb;
        src64 <= 12'hf68;
        src65 <= 12'hc05;
        src66 <= 12'hd34;
        src67 <= 12'h87f;
        src68 <= 12'hd2c;
        src69 <= 12'h6a;
        src70 <= 12'ha06;
        src71 <= 12'h633;
        src72 <= 12'h6ad;
        src73 <= 12'hfd9;
        src74 <= 12'h33b;
        src75 <= 12'h7b7;
        src76 <= 12'h24f;
        src77 <= 12'hcfa;
        src78 <= 12'h208;
        src79 <= 12'h76b;
        src80 <= 12'hc8a;
        src81 <= 12'h612;
        src82 <= 12'he79;
        src83 <= 12'hfe6;
        src84 <= 12'hd9a;
        src85 <= 12'h6b7;
        src86 <= 12'h38d;
        src87 <= 12'h198;
        src88 <= 12'h1a1;
        src89 <= 12'h4f3;
        src90 <= 12'h38a;
        src91 <= 12'h698;
        src92 <= 12'h12d;
        src93 <= 12'h95d;
        src94 <= 12'hfa1;
        src95 <= 12'hbe;
        src96 <= 12'ha6e;
        src97 <= 12'h896;
        src98 <= 12'hc1f;
        src99 <= 12'he4b;
        src100 <= 12'h3a4;
        src101 <= 12'hf39;
        src102 <= 12'h9dd;
        src103 <= 12'hc76;
        src104 <= 12'hfd7;
        src105 <= 12'h1e;
        src106 <= 12'h3a2;
        src107 <= 12'h4ca;
        src108 <= 12'hc8;
        src109 <= 12'h68b;
        src110 <= 12'hb6f;
        src111 <= 12'h897;
        src112 <= 12'hb53;
        src113 <= 12'h844;
        src114 <= 12'h295;
        src115 <= 12'h7b3;
        src116 <= 12'h887;
        src117 <= 12'h995;
        src118 <= 12'hebc;
        src119 <= 12'he2f;
        src120 <= 12'h94f;
        src121 <= 12'h372;
        src122 <= 12'h4df;
        src123 <= 12'h147;
        src124 <= 12'he85;
        src125 <= 12'h83d;
        src126 <= 12'h106;
        src127 <= 12'h8bd;
        src128 <= 12'h851;
        src129 <= 12'h4bd;
        src130 <= 12'h309;
        src131 <= 12'h379;
        src132 <= 12'hdfe;
        src133 <= 12'h10a;
        src134 <= 12'h1b6;
        src135 <= 12'hc49;
        src136 <= 12'h330;
        src137 <= 12'h76;
        src138 <= 12'h32a;
        src139 <= 12'h5d8;
        src140 <= 12'h1cb;
        src141 <= 12'h8c7;
        src142 <= 12'h118;
        src143 <= 12'hf8;
        src144 <= 12'h68b;
        src145 <= 12'h8e4;
        src146 <= 12'h5fc;
        src147 <= 12'h3f6;
        src148 <= 12'h1af;
        src149 <= 12'hdf8;
        src150 <= 12'h823;
        src151 <= 12'h925;
        src152 <= 12'hd0a;
        src153 <= 12'h7e3;
        src154 <= 12'h104;
        src155 <= 12'h76f;
        src156 <= 12'hbde;
        src157 <= 12'h4eb;
        src158 <= 12'h868;
        src159 <= 12'h622;
        src160 <= 12'h94e;
        src161 <= 12'h390;
        exp <= 20'h514fe;
        #1
        src0 <= 12'h272;
        src1 <= 12'h6a3;
        src2 <= 12'haae;
        src3 <= 12'h62e;
        src4 <= 12'h760;
        src5 <= 12'h8a8;
        src6 <= 12'hfc4;
        src7 <= 12'h40;
        src8 <= 12'h77f;
        src9 <= 12'hd28;
        src10 <= 12'hd6b;
        src11 <= 12'hd99;
        src12 <= 12'hb3;
        src13 <= 12'he15;
        src14 <= 12'h6ce;
        src15 <= 12'h30e;
        src16 <= 12'h263;
        src17 <= 12'hccf;
        src18 <= 12'hf31;
        src19 <= 12'h1aa;
        src20 <= 12'h4d0;
        src21 <= 12'h56a;
        src22 <= 12'h51a;
        src23 <= 12'hba;
        src24 <= 12'h5b0;
        src25 <= 12'h7ec;
        src26 <= 12'hd77;
        src27 <= 12'h9aa;
        src28 <= 12'h605;
        src29 <= 12'h75b;
        src30 <= 12'hda2;
        src31 <= 12'hb7a;
        src32 <= 12'h56a;
        src33 <= 12'ha76;
        src34 <= 12'h15e;
        src35 <= 12'ha4f;
        src36 <= 12'h80f;
        src37 <= 12'h31f;
        src38 <= 12'hfc5;
        src39 <= 12'h6b3;
        src40 <= 12'h1d7;
        src41 <= 12'h1cc;
        src42 <= 12'h688;
        src43 <= 12'hc64;
        src44 <= 12'hd2d;
        src45 <= 12'h8fb;
        src46 <= 12'h352;
        src47 <= 12'hb44;
        src48 <= 12'hc88;
        src49 <= 12'hc3c;
        src50 <= 12'hfd6;
        src51 <= 12'h2b3;
        src52 <= 12'hfb0;
        src53 <= 12'ha9;
        src54 <= 12'hc;
        src55 <= 12'h336;
        src56 <= 12'hb83;
        src57 <= 12'hc8d;
        src58 <= 12'ha65;
        src59 <= 12'h56;
        src60 <= 12'h22b;
        src61 <= 12'h816;
        src62 <= 12'hde3;
        src63 <= 12'h56a;
        src64 <= 12'hd8;
        src65 <= 12'h9fb;
        src66 <= 12'h342;
        src67 <= 12'ha6c;
        src68 <= 12'ha19;
        src69 <= 12'h18f;
        src70 <= 12'h23e;
        src71 <= 12'hdcb;
        src72 <= 12'hc0f;
        src73 <= 12'h4d5;
        src74 <= 12'he97;
        src75 <= 12'h862;
        src76 <= 12'h196;
        src77 <= 12'h39b;
        src78 <= 12'h153;
        src79 <= 12'h9e9;
        src80 <= 12'h4c2;
        src81 <= 12'hd98;
        src82 <= 12'hc15;
        src83 <= 12'h305;
        src84 <= 12'hc65;
        src85 <= 12'h8c9;
        src86 <= 12'hcd3;
        src87 <= 12'h814;
        src88 <= 12'h49b;
        src89 <= 12'hf4e;
        src90 <= 12'he25;
        src91 <= 12'hf54;
        src92 <= 12'h850;
        src93 <= 12'hb0e;
        src94 <= 12'he78;
        src95 <= 12'h8e3;
        src96 <= 12'hd24;
        src97 <= 12'hb86;
        src98 <= 12'hd4a;
        src99 <= 12'h7b6;
        src100 <= 12'h9d7;
        src101 <= 12'h455;
        src102 <= 12'h702;
        src103 <= 12'hf73;
        src104 <= 12'h66a;
        src105 <= 12'h1fa;
        src106 <= 12'hce4;
        src107 <= 12'haf9;
        src108 <= 12'h99;
        src109 <= 12'h77a;
        src110 <= 12'he51;
        src111 <= 12'haa8;
        src112 <= 12'hb0a;
        src113 <= 12'h87c;
        src114 <= 12'h593;
        src115 <= 12'hccc;
        src116 <= 12'h4c;
        src117 <= 12'hb65;
        src118 <= 12'h1ce;
        src119 <= 12'h244;
        src120 <= 12'h7fd;
        src121 <= 12'h2d6;
        src122 <= 12'h2c5;
        src123 <= 12'hfb0;
        src124 <= 12'had3;
        src125 <= 12'h30b;
        src126 <= 12'hca6;
        src127 <= 12'h8e8;
        src128 <= 12'h7cf;
        src129 <= 12'h341;
        src130 <= 12'h921;
        src131 <= 12'h626;
        src132 <= 12'h59d;
        src133 <= 12'h9a4;
        src134 <= 12'h5b9;
        src135 <= 12'h2dc;
        src136 <= 12'h56c;
        src137 <= 12'h83f;
        src138 <= 12'h350;
        src139 <= 12'h45f;
        src140 <= 12'h2e8;
        src141 <= 12'h1b7;
        src142 <= 12'h750;
        src143 <= 12'he67;
        src144 <= 12'hdb7;
        src145 <= 12'h169;
        src146 <= 12'ha28;
        src147 <= 12'h2a4;
        src148 <= 12'h616;
        src149 <= 12'hcef;
        src150 <= 12'h266;
        src151 <= 12'hcba;
        src152 <= 12'h136;
        src153 <= 12'h32a;
        src154 <= 12'h9fb;
        src155 <= 12'hcce;
        src156 <= 12'h30e;
        src157 <= 12'h38;
        src158 <= 12'h8bf;
        src159 <= 12'h7c6;
        src160 <= 12'h4f2;
        src161 <= 12'h292;
        exp <= 20'h4e9db;
        #1
        src0 <= 12'h77;
        src1 <= 12'h48a;
        src2 <= 12'hb4d;
        src3 <= 12'hc41;
        src4 <= 12'h1df;
        src5 <= 12'h3df;
        src6 <= 12'he95;
        src7 <= 12'h93e;
        src8 <= 12'h846;
        src9 <= 12'h34c;
        src10 <= 12'h612;
        src11 <= 12'h94c;
        src12 <= 12'h8cf;
        src13 <= 12'ha3a;
        src14 <= 12'h710;
        src15 <= 12'h6da;
        src16 <= 12'h1a6;
        src17 <= 12'ha97;
        src18 <= 12'ha6c;
        src19 <= 12'h4e;
        src20 <= 12'h323;
        src21 <= 12'h4df;
        src22 <= 12'h1c;
        src23 <= 12'h733;
        src24 <= 12'h44a;
        src25 <= 12'h151;
        src26 <= 12'hf54;
        src27 <= 12'h5d7;
        src28 <= 12'ha2f;
        src29 <= 12'h39;
        src30 <= 12'h12b;
        src31 <= 12'h407;
        src32 <= 12'h33e;
        src33 <= 12'h6c2;
        src34 <= 12'hb76;
        src35 <= 12'h79a;
        src36 <= 12'h301;
        src37 <= 12'h101;
        src38 <= 12'hbd2;
        src39 <= 12'hb05;
        src40 <= 12'hff4;
        src41 <= 12'he1c;
        src42 <= 12'h92d;
        src43 <= 12'hef5;
        src44 <= 12'hd82;
        src45 <= 12'hddf;
        src46 <= 12'haab;
        src47 <= 12'h1da;
        src48 <= 12'h3b7;
        src49 <= 12'hd91;
        src50 <= 12'h48e;
        src51 <= 12'hb3b;
        src52 <= 12'h810;
        src53 <= 12'h75d;
        src54 <= 12'h974;
        src55 <= 12'hc94;
        src56 <= 12'h8cb;
        src57 <= 12'hb99;
        src58 <= 12'hc94;
        src59 <= 12'h868;
        src60 <= 12'he79;
        src61 <= 12'h738;
        src62 <= 12'h47c;
        src63 <= 12'h878;
        src64 <= 12'h31b;
        src65 <= 12'hd64;
        src66 <= 12'h42a;
        src67 <= 12'h8ff;
        src68 <= 12'h9b5;
        src69 <= 12'h50c;
        src70 <= 12'h19a;
        src71 <= 12'he23;
        src72 <= 12'h888;
        src73 <= 12'hfc1;
        src74 <= 12'habf;
        src75 <= 12'h770;
        src76 <= 12'h469;
        src77 <= 12'ha47;
        src78 <= 12'h1e;
        src79 <= 12'h213;
        src80 <= 12'h5f1;
        src81 <= 12'h6e9;
        src82 <= 12'h297;
        src83 <= 12'h6f5;
        src84 <= 12'hcfc;
        src85 <= 12'h214;
        src86 <= 12'hfb8;
        src87 <= 12'h321;
        src88 <= 12'hf4c;
        src89 <= 12'h6c6;
        src90 <= 12'hc8a;
        src91 <= 12'h21;
        src92 <= 12'h11;
        src93 <= 12'hc11;
        src94 <= 12'h4e4;
        src95 <= 12'h896;
        src96 <= 12'h526;
        src97 <= 12'he76;
        src98 <= 12'h6f7;
        src99 <= 12'hf93;
        src100 <= 12'h8d5;
        src101 <= 12'he9d;
        src102 <= 12'h7c;
        src103 <= 12'h24d;
        src104 <= 12'hcc2;
        src105 <= 12'hc77;
        src106 <= 12'hbf0;
        src107 <= 12'h3d;
        src108 <= 12'h995;
        src109 <= 12'ha9c;
        src110 <= 12'h440;
        src111 <= 12'h618;
        src112 <= 12'hcb6;
        src113 <= 12'h448;
        src114 <= 12'h2ba;
        src115 <= 12'h393;
        src116 <= 12'hd39;
        src117 <= 12'h152;
        src118 <= 12'h6e8;
        src119 <= 12'h9f0;
        src120 <= 12'hc81;
        src121 <= 12'ha2c;
        src122 <= 12'h991;
        src123 <= 12'h1cf;
        src124 <= 12'hc22;
        src125 <= 12'h1ec;
        src126 <= 12'h3bb;
        src127 <= 12'h76f;
        src128 <= 12'h406;
        src129 <= 12'hffe;
        src130 <= 12'hf71;
        src131 <= 12'hada;
        src132 <= 12'h126;
        src133 <= 12'ha7d;
        src134 <= 12'ha1a;
        src135 <= 12'h4d6;
        src136 <= 12'h8c2;
        src137 <= 12'hf18;
        src138 <= 12'h375;
        src139 <= 12'h311;
        src140 <= 12'h5e6;
        src141 <= 12'hacb;
        src142 <= 12'hfe8;
        src143 <= 12'hfcc;
        src144 <= 12'h358;
        src145 <= 12'hb7;
        src146 <= 12'h70d;
        src147 <= 12'h435;
        src148 <= 12'h2c9;
        src149 <= 12'hfc7;
        src150 <= 12'h2bc;
        src151 <= 12'ha2a;
        src152 <= 12'hf20;
        src153 <= 12'h560;
        src154 <= 12'h596;
        src155 <= 12'h164;
        src156 <= 12'h9d3;
        src157 <= 12'h72f;
        src158 <= 12'h657;
        src159 <= 12'hfba;
        src160 <= 12'ha2;
        src161 <= 12'h273;
        exp <= 20'h4e1b1;
        #1
        src0 <= 12'haaa;
        src1 <= 12'h891;
        src2 <= 12'he9b;
        src3 <= 12'h39c;
        src4 <= 12'h1ca;
        src5 <= 12'h13d;
        src6 <= 12'he87;
        src7 <= 12'h83f;
        src8 <= 12'h1cf;
        src9 <= 12'h21d;
        src10 <= 12'h9b0;
        src11 <= 12'hc03;
        src12 <= 12'hd69;
        src13 <= 12'hb91;
        src14 <= 12'h678;
        src15 <= 12'hd14;
        src16 <= 12'h834;
        src17 <= 12'h43d;
        src18 <= 12'h4ec;
        src19 <= 12'h46;
        src20 <= 12'hbdc;
        src21 <= 12'ha1f;
        src22 <= 12'h6ce;
        src23 <= 12'he1c;
        src24 <= 12'hbce;
        src25 <= 12'h12e;
        src26 <= 12'ha2d;
        src27 <= 12'h4d6;
        src28 <= 12'hc63;
        src29 <= 12'h831;
        src30 <= 12'hb2a;
        src31 <= 12'hfd1;
        src32 <= 12'h5ae;
        src33 <= 12'hed0;
        src34 <= 12'hfae;
        src35 <= 12'ha4f;
        src36 <= 12'h9b1;
        src37 <= 12'he17;
        src38 <= 12'h18a;
        src39 <= 12'h99b;
        src40 <= 12'hc4b;
        src41 <= 12'h246;
        src42 <= 12'hed4;
        src43 <= 12'h1dd;
        src44 <= 12'h39f;
        src45 <= 12'he8f;
        src46 <= 12'h194;
        src47 <= 12'h9f6;
        src48 <= 12'hb5c;
        src49 <= 12'hc13;
        src50 <= 12'h5c5;
        src51 <= 12'h65f;
        src52 <= 12'hf10;
        src53 <= 12'hec7;
        src54 <= 12'hafb;
        src55 <= 12'ha56;
        src56 <= 12'h783;
        src57 <= 12'hdf2;
        src58 <= 12'h867;
        src59 <= 12'hf11;
        src60 <= 12'hfc;
        src61 <= 12'h402;
        src62 <= 12'h50c;
        src63 <= 12'h2c1;
        src64 <= 12'he95;
        src65 <= 12'he15;
        src66 <= 12'h3a7;
        src67 <= 12'h4f4;
        src68 <= 12'h239;
        src69 <= 12'hf11;
        src70 <= 12'h172;
        src71 <= 12'h97;
        src72 <= 12'h873;
        src73 <= 12'h5f3;
        src74 <= 12'h27b;
        src75 <= 12'hd20;
        src76 <= 12'h231;
        src77 <= 12'h615;
        src78 <= 12'h983;
        src79 <= 12'hc81;
        src80 <= 12'he9f;
        src81 <= 12'h3b6;
        src82 <= 12'h896;
        src83 <= 12'ha3b;
        src84 <= 12'h160;
        src85 <= 12'hed9;
        src86 <= 12'h48e;
        src87 <= 12'h278;
        src88 <= 12'h69e;
        src89 <= 12'ha6c;
        src90 <= 12'h244;
        src91 <= 12'hd24;
        src92 <= 12'h8dd;
        src93 <= 12'hfc5;
        src94 <= 12'hffa;
        src95 <= 12'h557;
        src96 <= 12'h9ed;
        src97 <= 12'heff;
        src98 <= 12'h5bd;
        src99 <= 12'hc83;
        src100 <= 12'h253;
        src101 <= 12'hec1;
        src102 <= 12'ha5a;
        src103 <= 12'hf90;
        src104 <= 12'h11b;
        src105 <= 12'hf1e;
        src106 <= 12'h36;
        src107 <= 12'h8fd;
        src108 <= 12'h276;
        src109 <= 12'hc9a;
        src110 <= 12'hafd;
        src111 <= 12'h9;
        src112 <= 12'h7c1;
        src113 <= 12'h284;
        src114 <= 12'h805;
        src115 <= 12'h9fc;
        src116 <= 12'h853;
        src117 <= 12'h88;
        src118 <= 12'h68f;
        src119 <= 12'hc92;
        src120 <= 12'he24;
        src121 <= 12'hc60;
        src122 <= 12'hc6f;
        src123 <= 12'hd2b;
        src124 <= 12'h64e;
        src125 <= 12'h7a8;
        src126 <= 12'hb78;
        src127 <= 12'h418;
        src128 <= 12'hd4a;
        src129 <= 12'haea;
        src130 <= 12'ha8;
        src131 <= 12'hb53;
        src132 <= 12'h5c6;
        src133 <= 12'h7bc;
        src134 <= 12'h884;
        src135 <= 12'h721;
        src136 <= 12'h271;
        src137 <= 12'h369;
        src138 <= 12'hf44;
        src139 <= 12'h2dc;
        src140 <= 12'h44a;
        src141 <= 12'h155;
        src142 <= 12'hdbc;
        src143 <= 12'h752;
        src144 <= 12'h67f;
        src145 <= 12'h702;
        src146 <= 12'he15;
        src147 <= 12'h6f2;
        src148 <= 12'hd36;
        src149 <= 12'h995;
        src150 <= 12'h722;
        src151 <= 12'h655;
        src152 <= 12'h205;
        src153 <= 12'hfa3;
        src154 <= 12'h924;
        src155 <= 12'hdd0;
        src156 <= 12'h3a1;
        src157 <= 12'h1f6;
        src158 <= 12'he56;
        src159 <= 12'h3ed;
        src160 <= 12'h386;
        src161 <= 12'hd30;
        exp <= 20'h54b81;
        #1
        src0 <= 12'h353;
        src1 <= 12'h5d7;
        src2 <= 12'h513;
        src3 <= 12'h150;
        src4 <= 12'h549;
        src5 <= 12'h485;
        src6 <= 12'h89e;
        src7 <= 12'hdd6;
        src8 <= 12'hf43;
        src9 <= 12'hbe1;
        src10 <= 12'h9f;
        src11 <= 12'hb8;
        src12 <= 12'ha78;
        src13 <= 12'h4f1;
        src14 <= 12'hd2;
        src15 <= 12'h2b0;
        src16 <= 12'h524;
        src17 <= 12'h5aa;
        src18 <= 12'h663;
        src19 <= 12'h9d1;
        src20 <= 12'h64e;
        src21 <= 12'hfb7;
        src22 <= 12'hcfe;
        src23 <= 12'hc8c;
        src24 <= 12'h398;
        src25 <= 12'h911;
        src26 <= 12'h3c;
        src27 <= 12'h36c;
        src28 <= 12'hf1f;
        src29 <= 12'hbc;
        src30 <= 12'h4d8;
        src31 <= 12'h3b8;
        src32 <= 12'ha15;
        src33 <= 12'hca8;
        src34 <= 12'hcc5;
        src35 <= 12'h33d;
        src36 <= 12'hb18;
        src37 <= 12'h2ad;
        src38 <= 12'hbd0;
        src39 <= 12'hc4b;
        src40 <= 12'h6d9;
        src41 <= 12'h179;
        src42 <= 12'hed1;
        src43 <= 12'hcf1;
        src44 <= 12'haa0;
        src45 <= 12'h155;
        src46 <= 12'h22c;
        src47 <= 12'h4bc;
        src48 <= 12'h61c;
        src49 <= 12'h38b;
        src50 <= 12'hf2b;
        src51 <= 12'hd30;
        src52 <= 12'h82c;
        src53 <= 12'he29;
        src54 <= 12'h7e7;
        src55 <= 12'ha83;
        src56 <= 12'h9c;
        src57 <= 12'h88;
        src58 <= 12'h18a;
        src59 <= 12'ha44;
        src60 <= 12'hefe;
        src61 <= 12'h656;
        src62 <= 12'h316;
        src63 <= 12'h479;
        src64 <= 12'ha10;
        src65 <= 12'ha51;
        src66 <= 12'h672;
        src67 <= 12'hd75;
        src68 <= 12'hb6e;
        src69 <= 12'h462;
        src70 <= 12'h16f;
        src71 <= 12'h293;
        src72 <= 12'hcb6;
        src73 <= 12'hba;
        src74 <= 12'ha38;
        src75 <= 12'h7c8;
        src76 <= 12'h664;
        src77 <= 12'hc5c;
        src78 <= 12'hafb;
        src79 <= 12'h23c;
        src80 <= 12'h5d5;
        src81 <= 12'h630;
        src82 <= 12'h26e;
        src83 <= 12'haa0;
        src84 <= 12'h15;
        src85 <= 12'ha54;
        src86 <= 12'h11;
        src87 <= 12'hd36;
        src88 <= 12'hb57;
        src89 <= 12'haa8;
        src90 <= 12'h118;
        src91 <= 12'h113;
        src92 <= 12'hbc4;
        src93 <= 12'h8ae;
        src94 <= 12'h50c;
        src95 <= 12'h6de;
        src96 <= 12'hd91;
        src97 <= 12'h2e5;
        src98 <= 12'hd07;
        src99 <= 12'h84d;
        src100 <= 12'hfc6;
        src101 <= 12'h969;
        src102 <= 12'he36;
        src103 <= 12'h64a;
        src104 <= 12'hc0d;
        src105 <= 12'h7cd;
        src106 <= 12'hc66;
        src107 <= 12'h13b;
        src108 <= 12'h148;
        src109 <= 12'h8f0;
        src110 <= 12'h178;
        src111 <= 12'h992;
        src112 <= 12'hf43;
        src113 <= 12'h136;
        src114 <= 12'h5f1;
        src115 <= 12'hf09;
        src116 <= 12'hffa;
        src117 <= 12'h82;
        src118 <= 12'h6ed;
        src119 <= 12'hf9b;
        src120 <= 12'he3d;
        src121 <= 12'he78;
        src122 <= 12'h512;
        src123 <= 12'h5bf;
        src124 <= 12'h1de;
        src125 <= 12'hb81;
        src126 <= 12'h4dc;
        src127 <= 12'h1bb;
        src128 <= 12'h74b;
        src129 <= 12'h4d5;
        src130 <= 12'h906;
        src131 <= 12'h46d;
        src132 <= 12'h377;
        src133 <= 12'hbdd;
        src134 <= 12'h31;
        src135 <= 12'he16;
        src136 <= 12'hd6;
        src137 <= 12'he49;
        src138 <= 12'h29b;
        src139 <= 12'h768;
        src140 <= 12'hf1a;
        src141 <= 12'had8;
        src142 <= 12'hde;
        src143 <= 12'h347;
        src144 <= 12'h99c;
        src145 <= 12'h769;
        src146 <= 12'h924;
        src147 <= 12'h149;
        src148 <= 12'h78e;
        src149 <= 12'hd94;
        src150 <= 12'h9fd;
        src151 <= 12'h925;
        src152 <= 12'h13a;
        src153 <= 12'h469;
        src154 <= 12'hb61;
        src155 <= 12'he11;
        src156 <= 12'hd4f;
        src157 <= 12'h25e;
        src158 <= 12'h92e;
        src159 <= 12'hff6;
        src160 <= 12'h6d8;
        src161 <= 12'h5d0;
        exp <= 20'h4cc46;
        #1
        src0 <= 12'h6d9;
        src1 <= 12'h6ac;
        src2 <= 12'h968;
        src3 <= 12'ha9f;
        src4 <= 12'h820;
        src5 <= 12'h238;
        src6 <= 12'hc44;
        src7 <= 12'h165;
        src8 <= 12'h4c5;
        src9 <= 12'h4bb;
        src10 <= 12'hb14;
        src11 <= 12'h9f6;
        src12 <= 12'h956;
        src13 <= 12'h5bc;
        src14 <= 12'h6f4;
        src15 <= 12'h7c9;
        src16 <= 12'hc5b;
        src17 <= 12'hf1b;
        src18 <= 12'h4cb;
        src19 <= 12'h828;
        src20 <= 12'hb7b;
        src21 <= 12'h749;
        src22 <= 12'h96c;
        src23 <= 12'ha93;
        src24 <= 12'h89a;
        src25 <= 12'hb35;
        src26 <= 12'h60b;
        src27 <= 12'h6c8;
        src28 <= 12'hc8;
        src29 <= 12'h89b;
        src30 <= 12'ha83;
        src31 <= 12'h384;
        src32 <= 12'hac8;
        src33 <= 12'hee9;
        src34 <= 12'h422;
        src35 <= 12'hae9;
        src36 <= 12'h7bf;
        src37 <= 12'hdaf;
        src38 <= 12'hc18;
        src39 <= 12'hb7b;
        src40 <= 12'ha61;
        src41 <= 12'hdde;
        src42 <= 12'h216;
        src43 <= 12'h7a3;
        src44 <= 12'h42a;
        src45 <= 12'h879;
        src46 <= 12'h15e;
        src47 <= 12'h943;
        src48 <= 12'h58d;
        src49 <= 12'h8e9;
        src50 <= 12'h2a6;
        src51 <= 12'h14;
        src52 <= 12'h8d3;
        src53 <= 12'he59;
        src54 <= 12'h2a3;
        src55 <= 12'hde9;
        src56 <= 12'h42d;
        src57 <= 12'h203;
        src58 <= 12'h238;
        src59 <= 12'h294;
        src60 <= 12'h3f5;
        src61 <= 12'hdce;
        src62 <= 12'h40c;
        src63 <= 12'h4b5;
        src64 <= 12'hf77;
        src65 <= 12'hd41;
        src66 <= 12'h22f;
        src67 <= 12'he26;
        src68 <= 12'ha5b;
        src69 <= 12'h204;
        src70 <= 12'hb3d;
        src71 <= 12'hd2d;
        src72 <= 12'he6a;
        src73 <= 12'h2f7;
        src74 <= 12'h9d1;
        src75 <= 12'h48f;
        src76 <= 12'h7df;
        src77 <= 12'h6e1;
        src78 <= 12'h6ed;
        src79 <= 12'he73;
        src80 <= 12'h85b;
        src81 <= 12'h16e;
        src82 <= 12'h9bb;
        src83 <= 12'h328;
        src84 <= 12'h782;
        src85 <= 12'ha04;
        src86 <= 12'h7aa;
        src87 <= 12'h6e1;
        src88 <= 12'h2ac;
        src89 <= 12'hdb6;
        src90 <= 12'h192;
        src91 <= 12'h9ac;
        src92 <= 12'h7be;
        src93 <= 12'h937;
        src94 <= 12'he06;
        src95 <= 12'hfb8;
        src96 <= 12'hd19;
        src97 <= 12'h31;
        src98 <= 12'hc94;
        src99 <= 12'h85e;
        src100 <= 12'h54f;
        src101 <= 12'hc6;
        src102 <= 12'h20a;
        src103 <= 12'h4cd;
        src104 <= 12'h78a;
        src105 <= 12'h5a;
        src106 <= 12'ha5d;
        src107 <= 12'h5a8;
        src108 <= 12'hed1;
        src109 <= 12'h376;
        src110 <= 12'h505;
        src111 <= 12'hc72;
        src112 <= 12'hfe3;
        src113 <= 12'h1e8;
        src114 <= 12'h33;
        src115 <= 12'hfff;
        src116 <= 12'h14;
        src117 <= 12'h1b0;
        src118 <= 12'had9;
        src119 <= 12'h383;
        src120 <= 12'h186;
        src121 <= 12'hb7a;
        src122 <= 12'h93a;
        src123 <= 12'h61d;
        src124 <= 12'h3bf;
        src125 <= 12'h514;
        src126 <= 12'hc5e;
        src127 <= 12'hb1a;
        src128 <= 12'h56c;
        src129 <= 12'h73a;
        src130 <= 12'h935;
        src131 <= 12'hb4a;
        src132 <= 12'hfe3;
        src133 <= 12'h7ae;
        src134 <= 12'h506;
        src135 <= 12'h64a;
        src136 <= 12'h2d5;
        src137 <= 12'h4bb;
        src138 <= 12'h7e3;
        src139 <= 12'hd7f;
        src140 <= 12'hd23;
        src141 <= 12'h436;
        src142 <= 12'h7;
        src143 <= 12'hb20;
        src144 <= 12'h669;
        src145 <= 12'hab1;
        src146 <= 12'hf47;
        src147 <= 12'hfe2;
        src148 <= 12'hc18;
        src149 <= 12'h811;
        src150 <= 12'hd4;
        src151 <= 12'h98b;
        src152 <= 12'hcb;
        src153 <= 12'hf04;
        src154 <= 12'h7ec;
        src155 <= 12'h90b;
        src156 <= 12'h78a;
        src157 <= 12'h2;
        src158 <= 12'hdec;
        src159 <= 12'h4ef;
        src160 <= 12'h7e1;
        src161 <= 12'h5ec;
        exp <= 20'h4f011;
        #1
        src0 <= 12'hcdd;
        src1 <= 12'hb38;
        src2 <= 12'h6fe;
        src3 <= 12'hb6f;
        src4 <= 12'h3a6;
        src5 <= 12'h273;
        src6 <= 12'h774;
        src7 <= 12'hcf3;
        src8 <= 12'hc2d;
        src9 <= 12'h94d;
        src10 <= 12'h835;
        src11 <= 12'hfd6;
        src12 <= 12'h185;
        src13 <= 12'h6de;
        src14 <= 12'hc9c;
        src15 <= 12'h220;
        src16 <= 12'head;
        src17 <= 12'h632;
        src18 <= 12'h937;
        src19 <= 12'hfcb;
        src20 <= 12'hea7;
        src21 <= 12'ha08;
        src22 <= 12'heaa;
        src23 <= 12'h37d;
        src24 <= 12'hbbb;
        src25 <= 12'h916;
        src26 <= 12'h38b;
        src27 <= 12'h168;
        src28 <= 12'hdb3;
        src29 <= 12'h145;
        src30 <= 12'h155;
        src31 <= 12'h701;
        src32 <= 12'hca4;
        src33 <= 12'h23a;
        src34 <= 12'h431;
        src35 <= 12'h169;
        src36 <= 12'hdc1;
        src37 <= 12'ha81;
        src38 <= 12'hd2e;
        src39 <= 12'h663;
        src40 <= 12'h25d;
        src41 <= 12'hc2a;
        src42 <= 12'h559;
        src43 <= 12'h5a0;
        src44 <= 12'hf96;
        src45 <= 12'ha2b;
        src46 <= 12'h320;
        src47 <= 12'h67d;
        src48 <= 12'h79a;
        src49 <= 12'hacf;
        src50 <= 12'h1c0;
        src51 <= 12'hc04;
        src52 <= 12'hbd4;
        src53 <= 12'h965;
        src54 <= 12'h7db;
        src55 <= 12'hbd8;
        src56 <= 12'h90;
        src57 <= 12'ha87;
        src58 <= 12'h273;
        src59 <= 12'hdbf;
        src60 <= 12'h77c;
        src61 <= 12'h30d;
        src62 <= 12'hd0e;
        src63 <= 12'hea1;
        src64 <= 12'h81b;
        src65 <= 12'h44b;
        src66 <= 12'hb66;
        src67 <= 12'hfbb;
        src68 <= 12'h89b;
        src69 <= 12'h1ab;
        src70 <= 12'h879;
        src71 <= 12'hd3b;
        src72 <= 12'h34a;
        src73 <= 12'hbf7;
        src74 <= 12'hfa6;
        src75 <= 12'hc91;
        src76 <= 12'hf88;
        src77 <= 12'h2a2;
        src78 <= 12'h13b;
        src79 <= 12'h1cc;
        src80 <= 12'ha4f;
        src81 <= 12'h376;
        src82 <= 12'hcc7;
        src83 <= 12'h6bb;
        src84 <= 12'ha44;
        src85 <= 12'hd5c;
        src86 <= 12'hddd;
        src87 <= 12'hcff;
        src88 <= 12'hefe;
        src89 <= 12'hdfa;
        src90 <= 12'h25e;
        src91 <= 12'h11a;
        src92 <= 12'h48d;
        src93 <= 12'hbce;
        src94 <= 12'hfa;
        src95 <= 12'h45a;
        src96 <= 12'h200;
        src97 <= 12'he00;
        src98 <= 12'h2bf;
        src99 <= 12'h87e;
        src100 <= 12'haee;
        src101 <= 12'h245;
        src102 <= 12'h189;
        src103 <= 12'h5c2;
        src104 <= 12'h358;
        src105 <= 12'h1db;
        src106 <= 12'h743;
        src107 <= 12'he0e;
        src108 <= 12'he91;
        src109 <= 12'h81b;
        src110 <= 12'hf9;
        src111 <= 12'hffe;
        src112 <= 12'hd67;
        src113 <= 12'h67b;
        src114 <= 12'h96a;
        src115 <= 12'h1f5;
        src116 <= 12'h6a1;
        src117 <= 12'h7c2;
        src118 <= 12'h769;
        src119 <= 12'h1a7;
        src120 <= 12'hd2;
        src121 <= 12'h505;
        src122 <= 12'h2f8;
        src123 <= 12'h8f2;
        src124 <= 12'h6f1;
        src125 <= 12'h8e3;
        src126 <= 12'h185;
        src127 <= 12'h387;
        src128 <= 12'h5de;
        src129 <= 12'hfc5;
        src130 <= 12'he0b;
        src131 <= 12'h3f2;
        src132 <= 12'h7e1;
        src133 <= 12'h97c;
        src134 <= 12'h999;
        src135 <= 12'h84e;
        src136 <= 12'h80b;
        src137 <= 12'h11e;
        src138 <= 12'h48c;
        src139 <= 12'h751;
        src140 <= 12'h4bd;
        src141 <= 12'hbc7;
        src142 <= 12'h1f1;
        src143 <= 12'h2f4;
        src144 <= 12'hce6;
        src145 <= 12'ha09;
        src146 <= 12'h279;
        src147 <= 12'h20d;
        src148 <= 12'h75f;
        src149 <= 12'hd5b;
        src150 <= 12'h13;
        src151 <= 12'h6c0;
        src152 <= 12'h2ea;
        src153 <= 12'hcf5;
        src154 <= 12'h6ef;
        src155 <= 12'hfcf;
        src156 <= 12'he73;
        src157 <= 12'h5b0;
        src158 <= 12'h74e;
        src159 <= 12'h14d;
        src160 <= 12'h793;
        src161 <= 12'h3c9;
        exp <= 20'h4f781;
        #1
        src0 <= 12'h306;
        src1 <= 12'h596;
        src2 <= 12'hef2;
        src3 <= 12'h110;
        src4 <= 12'h849;
        src5 <= 12'h7f7;
        src6 <= 12'h399;
        src7 <= 12'h103;
        src8 <= 12'h5f5;
        src9 <= 12'hba0;
        src10 <= 12'h538;
        src11 <= 12'h676;
        src12 <= 12'h787;
        src13 <= 12'h2e7;
        src14 <= 12'ha10;
        src15 <= 12'hbe7;
        src16 <= 12'h8bd;
        src17 <= 12'h9a;
        src18 <= 12'h52d;
        src19 <= 12'h12;
        src20 <= 12'h7c6;
        src21 <= 12'h7ad;
        src22 <= 12'h87e;
        src23 <= 12'h574;
        src24 <= 12'h6e9;
        src25 <= 12'h62e;
        src26 <= 12'h25c;
        src27 <= 12'h5d7;
        src28 <= 12'h26a;
        src29 <= 12'he31;
        src30 <= 12'h447;
        src31 <= 12'h87e;
        src32 <= 12'h98b;
        src33 <= 12'hbe;
        src34 <= 12'h1d0;
        src35 <= 12'hc82;
        src36 <= 12'h7bb;
        src37 <= 12'hb2a;
        src38 <= 12'hd24;
        src39 <= 12'hba7;
        src40 <= 12'h629;
        src41 <= 12'he16;
        src42 <= 12'hb7;
        src43 <= 12'h6bf;
        src44 <= 12'h9cd;
        src45 <= 12'hcab;
        src46 <= 12'h539;
        src47 <= 12'hb9d;
        src48 <= 12'h20d;
        src49 <= 12'hb69;
        src50 <= 12'hd0c;
        src51 <= 12'hc64;
        src52 <= 12'hed8;
        src53 <= 12'hddd;
        src54 <= 12'h296;
        src55 <= 12'h258;
        src56 <= 12'h1dc;
        src57 <= 12'h3ce;
        src58 <= 12'h1bd;
        src59 <= 12'h681;
        src60 <= 12'h904;
        src61 <= 12'hae;
        src62 <= 12'hb1b;
        src63 <= 12'h81b;
        src64 <= 12'he96;
        src65 <= 12'hbcb;
        src66 <= 12'h432;
        src67 <= 12'hd9a;
        src68 <= 12'h2b1;
        src69 <= 12'h79d;
        src70 <= 12'h68e;
        src71 <= 12'h2e6;
        src72 <= 12'h548;
        src73 <= 12'hadd;
        src74 <= 12'hb65;
        src75 <= 12'ha73;
        src76 <= 12'h696;
        src77 <= 12'hed3;
        src78 <= 12'h131;
        src79 <= 12'hbd5;
        src80 <= 12'haa7;
        src81 <= 12'h14;
        src82 <= 12'h6c2;
        src83 <= 12'h644;
        src84 <= 12'he73;
        src85 <= 12'h512;
        src86 <= 12'h7cb;
        src87 <= 12'h57;
        src88 <= 12'h48;
        src89 <= 12'h5f6;
        src90 <= 12'h781;
        src91 <= 12'h821;
        src92 <= 12'h6d4;
        src93 <= 12'h6be;
        src94 <= 12'h462;
        src95 <= 12'h1c9;
        src96 <= 12'hcdf;
        src97 <= 12'h26c;
        src98 <= 12'h59c;
        src99 <= 12'hb67;
        src100 <= 12'h4b0;
        src101 <= 12'hc49;
        src102 <= 12'h234;
        src103 <= 12'h4ef;
        src104 <= 12'hf93;
        src105 <= 12'h4ae;
        src106 <= 12'ha4c;
        src107 <= 12'h7be;
        src108 <= 12'h78d;
        src109 <= 12'h778;
        src110 <= 12'h2d1;
        src111 <= 12'h6ba;
        src112 <= 12'he0;
        src113 <= 12'hd70;
        src114 <= 12'hc78;
        src115 <= 12'h3bd;
        src116 <= 12'h3da;
        src117 <= 12'h3dc;
        src118 <= 12'hd1d;
        src119 <= 12'h19f;
        src120 <= 12'hd33;
        src121 <= 12'h68e;
        src122 <= 12'h1a6;
        src123 <= 12'h97;
        src124 <= 12'h74d;
        src125 <= 12'heb;
        src126 <= 12'hcb5;
        src127 <= 12'he7c;
        src128 <= 12'hbbb;
        src129 <= 12'hb57;
        src130 <= 12'h68d;
        src131 <= 12'hb30;
        src132 <= 12'h5ed;
        src133 <= 12'hab4;
        src134 <= 12'hdc1;
        src135 <= 12'ha70;
        src136 <= 12'h1eb;
        src137 <= 12'h6e6;
        src138 <= 12'h13b;
        src139 <= 12'h132;
        src140 <= 12'hf95;
        src141 <= 12'h96c;
        src142 <= 12'ha34;
        src143 <= 12'hebe;
        src144 <= 12'ha07;
        src145 <= 12'haf5;
        src146 <= 12'h39f;
        src147 <= 12'hd05;
        src148 <= 12'hf00;
        src149 <= 12'h6f5;
        src150 <= 12'h865;
        src151 <= 12'h546;
        src152 <= 12'h15c;
        src153 <= 12'he8e;
        src154 <= 12'h556;
        src155 <= 12'he43;
        src156 <= 12'ha16;
        src157 <= 12'h700;
        src158 <= 12'h1d0;
        src159 <= 12'h20c;
        src160 <= 12'h3a4;
        src161 <= 12'hfac;
        exp <= 20'h4b348;
        #1
        src0 <= 12'h696;
        src1 <= 12'h25a;
        src2 <= 12'hbf;
        src3 <= 12'h527;
        src4 <= 12'he02;
        src5 <= 12'hab3;
        src6 <= 12'hfe2;
        src7 <= 12'h7;
        src8 <= 12'hc51;
        src9 <= 12'h77b;
        src10 <= 12'h5ed;
        src11 <= 12'h456;
        src12 <= 12'hb91;
        src13 <= 12'hbd0;
        src14 <= 12'h238;
        src15 <= 12'h63;
        src16 <= 12'h6bb;
        src17 <= 12'h87d;
        src18 <= 12'h6ca;
        src19 <= 12'hbfa;
        src20 <= 12'h277;
        src21 <= 12'hbdf;
        src22 <= 12'h81c;
        src23 <= 12'hff6;
        src24 <= 12'h5aa;
        src25 <= 12'h532;
        src26 <= 12'h368;
        src27 <= 12'hfd9;
        src28 <= 12'h90d;
        src29 <= 12'hd59;
        src30 <= 12'h669;
        src31 <= 12'h983;
        src32 <= 12'h7d;
        src33 <= 12'h282;
        src34 <= 12'hb9a;
        src35 <= 12'h2ef;
        src36 <= 12'hecb;
        src37 <= 12'h795;
        src38 <= 12'h1df;
        src39 <= 12'h5bc;
        src40 <= 12'h25f;
        src41 <= 12'h1cf;
        src42 <= 12'hb88;
        src43 <= 12'h57b;
        src44 <= 12'h85d;
        src45 <= 12'h9bb;
        src46 <= 12'h262;
        src47 <= 12'h9ed;
        src48 <= 12'h509;
        src49 <= 12'hbb3;
        src50 <= 12'he1f;
        src51 <= 12'h353;
        src52 <= 12'h5f3;
        src53 <= 12'h999;
        src54 <= 12'h7c2;
        src55 <= 12'hcd1;
        src56 <= 12'h3d5;
        src57 <= 12'h7e2;
        src58 <= 12'hdd4;
        src59 <= 12'hfde;
        src60 <= 12'h5e7;
        src61 <= 12'h966;
        src62 <= 12'hd86;
        src63 <= 12'h94a;
        src64 <= 12'hce5;
        src65 <= 12'hf3e;
        src66 <= 12'ha0f;
        src67 <= 12'h776;
        src68 <= 12'h58;
        src69 <= 12'h933;
        src70 <= 12'h216;
        src71 <= 12'h677;
        src72 <= 12'hea3;
        src73 <= 12'h627;
        src74 <= 12'haf5;
        src75 <= 12'h25;
        src76 <= 12'h8c5;
        src77 <= 12'hfad;
        src78 <= 12'h11b;
        src79 <= 12'h4f1;
        src80 <= 12'hb44;
        src81 <= 12'hdf6;
        src82 <= 12'h992;
        src83 <= 12'h944;
        src84 <= 12'h84c;
        src85 <= 12'ha2e;
        src86 <= 12'hd9b;
        src87 <= 12'hd2e;
        src88 <= 12'h915;
        src89 <= 12'h52d;
        src90 <= 12'h914;
        src91 <= 12'h7d1;
        src92 <= 12'he6c;
        src93 <= 12'h963;
        src94 <= 12'hfb7;
        src95 <= 12'hb27;
        src96 <= 12'hfcd;
        src97 <= 12'hc6a;
        src98 <= 12'hd4b;
        src99 <= 12'h1b7;
        src100 <= 12'h54;
        src101 <= 12'h99d;
        src102 <= 12'hf57;
        src103 <= 12'hb37;
        src104 <= 12'h24b;
        src105 <= 12'hc5;
        src106 <= 12'h2f0;
        src107 <= 12'hd03;
        src108 <= 12'h245;
        src109 <= 12'h358;
        src110 <= 12'h6eb;
        src111 <= 12'hd45;
        src112 <= 12'h7c9;
        src113 <= 12'h786;
        src114 <= 12'h82b;
        src115 <= 12'he4e;
        src116 <= 12'h33f;
        src117 <= 12'h99f;
        src118 <= 12'h4f2;
        src119 <= 12'h320;
        src120 <= 12'h916;
        src121 <= 12'hdbb;
        src122 <= 12'h5cd;
        src123 <= 12'h671;
        src124 <= 12'h4d3;
        src125 <= 12'h9f8;
        src126 <= 12'h9b5;
        src127 <= 12'h7a3;
        src128 <= 12'h3c0;
        src129 <= 12'h3db;
        src130 <= 12'h11e;
        src131 <= 12'h9d2;
        src132 <= 12'he07;
        src133 <= 12'hbf3;
        src134 <= 12'hf24;
        src135 <= 12'h73c;
        src136 <= 12'h94a;
        src137 <= 12'he51;
        src138 <= 12'h916;
        src139 <= 12'h525;
        src140 <= 12'he40;
        src141 <= 12'h89b;
        src142 <= 12'h54b;
        src143 <= 12'hdc9;
        src144 <= 12'h4df;
        src145 <= 12'h4a2;
        src146 <= 12'h6d1;
        src147 <= 12'he2c;
        src148 <= 12'haac;
        src149 <= 12'h20a;
        src150 <= 12'hf9f;
        src151 <= 12'h88a;
        src152 <= 12'h464;
        src153 <= 12'hbe5;
        src154 <= 12'h536;
        src155 <= 12'hd3e;
        src156 <= 12'h6e4;
        src157 <= 12'hacc;
        src158 <= 12'h59;
        src159 <= 12'h38b;
        src160 <= 12'hb4;
        src161 <= 12'h73d;
        exp <= 20'h52f44;
        #1
        src0 <= 12'h12a;
        src1 <= 12'he00;
        src2 <= 12'h2f5;
        src3 <= 12'hdf6;
        src4 <= 12'he10;
        src5 <= 12'h908;
        src6 <= 12'h83d;
        src7 <= 12'h599;
        src8 <= 12'hd05;
        src9 <= 12'h93c;
        src10 <= 12'h610;
        src11 <= 12'h14;
        src12 <= 12'h2a5;
        src13 <= 12'hee7;
        src14 <= 12'hdb1;
        src15 <= 12'hd46;
        src16 <= 12'h768;
        src17 <= 12'he26;
        src18 <= 12'h171;
        src19 <= 12'h1bb;
        src20 <= 12'h9fe;
        src21 <= 12'h4a3;
        src22 <= 12'hc42;
        src23 <= 12'hb15;
        src24 <= 12'h6a5;
        src25 <= 12'h8ef;
        src26 <= 12'hfc;
        src27 <= 12'h737;
        src28 <= 12'hc35;
        src29 <= 12'hc8c;
        src30 <= 12'hf38;
        src31 <= 12'h570;
        src32 <= 12'hfc4;
        src33 <= 12'h7f7;
        src34 <= 12'h109;
        src35 <= 12'hcc0;
        src36 <= 12'h671;
        src37 <= 12'hd2;
        src38 <= 12'h324;
        src39 <= 12'hbfd;
        src40 <= 12'hd81;
        src41 <= 12'h7f5;
        src42 <= 12'h83c;
        src43 <= 12'h6ac;
        src44 <= 12'h8ad;
        src45 <= 12'h2d7;
        src46 <= 12'h4b5;
        src47 <= 12'h391;
        src48 <= 12'hbc5;
        src49 <= 12'h12d;
        src50 <= 12'h9f7;
        src51 <= 12'hfb5;
        src52 <= 12'h565;
        src53 <= 12'h118;
        src54 <= 12'hb0;
        src55 <= 12'h7fd;
        src56 <= 12'hd24;
        src57 <= 12'h9db;
        src58 <= 12'h607;
        src59 <= 12'hd3e;
        src60 <= 12'h14;
        src61 <= 12'h46c;
        src62 <= 12'h191;
        src63 <= 12'he9f;
        src64 <= 12'h630;
        src65 <= 12'hf44;
        src66 <= 12'h8bc;
        src67 <= 12'hc6;
        src68 <= 12'h754;
        src69 <= 12'h472;
        src70 <= 12'h311;
        src71 <= 12'h24f;
        src72 <= 12'h408;
        src73 <= 12'h34f;
        src74 <= 12'h939;
        src75 <= 12'hf4d;
        src76 <= 12'h6f3;
        src77 <= 12'hb97;
        src78 <= 12'h67;
        src79 <= 12'h14b;
        src80 <= 12'hca0;
        src81 <= 12'h940;
        src82 <= 12'he2a;
        src83 <= 12'hcf6;
        src84 <= 12'h446;
        src85 <= 12'h999;
        src86 <= 12'h638;
        src87 <= 12'hcab;
        src88 <= 12'hee5;
        src89 <= 12'h877;
        src90 <= 12'hf50;
        src91 <= 12'ha0e;
        src92 <= 12'hd38;
        src93 <= 12'h69b;
        src94 <= 12'ha7c;
        src95 <= 12'hf96;
        src96 <= 12'h5f8;
        src97 <= 12'h3ec;
        src98 <= 12'h95d;
        src99 <= 12'h6bc;
        src100 <= 12'hd17;
        src101 <= 12'h310;
        src102 <= 12'hb05;
        src103 <= 12'h56f;
        src104 <= 12'h231;
        src105 <= 12'h61b;
        src106 <= 12'h277;
        src107 <= 12'h4eb;
        src108 <= 12'ha88;
        src109 <= 12'hc15;
        src110 <= 12'hb3d;
        src111 <= 12'hd3e;
        src112 <= 12'ha90;
        src113 <= 12'h2c1;
        src114 <= 12'hede;
        src115 <= 12'he6c;
        src116 <= 12'h81;
        src117 <= 12'h91c;
        src118 <= 12'h850;
        src119 <= 12'h162;
        src120 <= 12'h2d2;
        src121 <= 12'ha3f;
        src122 <= 12'hc42;
        src123 <= 12'h921;
        src124 <= 12'h7ba;
        src125 <= 12'h6f5;
        src126 <= 12'hddc;
        src127 <= 12'h3cd;
        src128 <= 12'hf09;
        src129 <= 12'h998;
        src130 <= 12'hfc1;
        src131 <= 12'h749;
        src132 <= 12'h6b0;
        src133 <= 12'h70;
        src134 <= 12'h4a0;
        src135 <= 12'hbcc;
        src136 <= 12'h580;
        src137 <= 12'hcab;
        src138 <= 12'h580;
        src139 <= 12'h7a2;
        src140 <= 12'h65f;
        src141 <= 12'ha79;
        src142 <= 12'hba9;
        src143 <= 12'h75c;
        src144 <= 12'h50d;
        src145 <= 12'h44e;
        src146 <= 12'h164;
        src147 <= 12'hbba;
        src148 <= 12'h175;
        src149 <= 12'h3f7;
        src150 <= 12'h8f9;
        src151 <= 12'h4e4;
        src152 <= 12'h70;
        src153 <= 12'h60d;
        src154 <= 12'h8ef;
        src155 <= 12'hf34;
        src156 <= 12'h745;
        src157 <= 12'hb2a;
        src158 <= 12'h3d5;
        src159 <= 12'h392;
        src160 <= 12'h86a;
        src161 <= 12'hef8;
        exp <= 20'h50d3e;
        #1
        src0 <= 12'h71e;
        src1 <= 12'heb;
        src2 <= 12'h1b3;
        src3 <= 12'hbc8;
        src4 <= 12'hb49;
        src5 <= 12'hd60;
        src6 <= 12'h81f;
        src7 <= 12'h489;
        src8 <= 12'h32e;
        src9 <= 12'h4ad;
        src10 <= 12'h86b;
        src11 <= 12'hf40;
        src12 <= 12'h4a6;
        src13 <= 12'h2ed;
        src14 <= 12'he53;
        src15 <= 12'hf49;
        src16 <= 12'h756;
        src17 <= 12'h17d;
        src18 <= 12'hddc;
        src19 <= 12'h5aa;
        src20 <= 12'h675;
        src21 <= 12'h342;
        src22 <= 12'hc2a;
        src23 <= 12'hb93;
        src24 <= 12'h4e1;
        src25 <= 12'h530;
        src26 <= 12'h671;
        src27 <= 12'h78f;
        src28 <= 12'h765;
        src29 <= 12'hc2;
        src30 <= 12'h100;
        src31 <= 12'hf2;
        src32 <= 12'h24b;
        src33 <= 12'h712;
        src34 <= 12'h31b;
        src35 <= 12'h76f;
        src36 <= 12'hde1;
        src37 <= 12'h5fa;
        src38 <= 12'h918;
        src39 <= 12'hcb3;
        src40 <= 12'h6d6;
        src41 <= 12'ha32;
        src42 <= 12'h23e;
        src43 <= 12'ha91;
        src44 <= 12'h585;
        src45 <= 12'h21d;
        src46 <= 12'ha1;
        src47 <= 12'hbbe;
        src48 <= 12'he71;
        src49 <= 12'ha7a;
        src50 <= 12'hb82;
        src51 <= 12'he73;
        src52 <= 12'h8ab;
        src53 <= 12'h114;
        src54 <= 12'h14;
        src55 <= 12'h626;
        src56 <= 12'h2d9;
        src57 <= 12'h44f;
        src58 <= 12'h425;
        src59 <= 12'h3d1;
        src60 <= 12'h18b;
        src61 <= 12'hb63;
        src62 <= 12'h305;
        src63 <= 12'hd3f;
        src64 <= 12'hc58;
        src65 <= 12'h30d;
        src66 <= 12'h8e9;
        src67 <= 12'hf22;
        src68 <= 12'he6d;
        src69 <= 12'h50a;
        src70 <= 12'hf47;
        src71 <= 12'he13;
        src72 <= 12'h615;
        src73 <= 12'h1d5;
        src74 <= 12'ha65;
        src75 <= 12'he24;
        src76 <= 12'h2e7;
        src77 <= 12'hb18;
        src78 <= 12'hd5;
        src79 <= 12'hd02;
        src80 <= 12'hb6;
        src81 <= 12'h2b;
        src82 <= 12'h30d;
        src83 <= 12'hc5c;
        src84 <= 12'hcb4;
        src85 <= 12'ha9;
        src86 <= 12'h123;
        src87 <= 12'h9a0;
        src88 <= 12'h85c;
        src89 <= 12'hc32;
        src90 <= 12'hc32;
        src91 <= 12'h1b5;
        src92 <= 12'hd69;
        src93 <= 12'ha9;
        src94 <= 12'h872;
        src95 <= 12'ha2f;
        src96 <= 12'h769;
        src97 <= 12'h965;
        src98 <= 12'h53;
        src99 <= 12'h25e;
        src100 <= 12'h7c1;
        src101 <= 12'hb0c;
        src102 <= 12'hd87;
        src103 <= 12'hf05;
        src104 <= 12'h1e5;
        src105 <= 12'hb7b;
        src106 <= 12'h7aa;
        src107 <= 12'h489;
        src108 <= 12'hb23;
        src109 <= 12'hb82;
        src110 <= 12'h4c5;
        src111 <= 12'hfe1;
        src112 <= 12'hf18;
        src113 <= 12'hd48;
        src114 <= 12'h164;
        src115 <= 12'h852;
        src116 <= 12'h8a4;
        src117 <= 12'haba;
        src118 <= 12'hc4b;
        src119 <= 12'h993;
        src120 <= 12'h14e;
        src121 <= 12'h76b;
        src122 <= 12'h42b;
        src123 <= 12'h510;
        src124 <= 12'hda1;
        src125 <= 12'h3be;
        src126 <= 12'hfaf;
        src127 <= 12'hb40;
        src128 <= 12'h6e4;
        src129 <= 12'h849;
        src130 <= 12'h12b;
        src131 <= 12'ha2c;
        src132 <= 12'h15b;
        src133 <= 12'h53b;
        src134 <= 12'hfb9;
        src135 <= 12'hc61;
        src136 <= 12'h7b7;
        src137 <= 12'h730;
        src138 <= 12'hbcf;
        src139 <= 12'he2;
        src140 <= 12'hbe8;
        src141 <= 12'h627;
        src142 <= 12'h3da;
        src143 <= 12'hbd4;
        src144 <= 12'h19b;
        src145 <= 12'h9ca;
        src146 <= 12'hb4b;
        src147 <= 12'h16e;
        src148 <= 12'h997;
        src149 <= 12'ha4c;
        src150 <= 12'h601;
        src151 <= 12'h1bf;
        src152 <= 12'hbc1;
        src153 <= 12'h49b;
        src154 <= 12'h8da;
        src155 <= 12'hea2;
        src156 <= 12'hf39;
        src157 <= 12'h8ad;
        src158 <= 12'h25f;
        src159 <= 12'hc50;
        src160 <= 12'h6d7;
        src161 <= 12'h5b9;
        exp <= 20'h4dcbc;
        #1
        src0 <= 12'h60;
        src1 <= 12'hc0a;
        src2 <= 12'h898;
        src3 <= 12'hea7;
        src4 <= 12'hbfb;
        src5 <= 12'h23f;
        src6 <= 12'h1fc;
        src7 <= 12'h65;
        src8 <= 12'ha23;
        src9 <= 12'h9e0;
        src10 <= 12'h7c6;
        src11 <= 12'hefe;
        src12 <= 12'h2b6;
        src13 <= 12'hd7;
        src14 <= 12'h799;
        src15 <= 12'h61f;
        src16 <= 12'h8e3;
        src17 <= 12'h7d;
        src18 <= 12'h47c;
        src19 <= 12'h639;
        src20 <= 12'hbdf;
        src21 <= 12'hb43;
        src22 <= 12'hd8c;
        src23 <= 12'h3e0;
        src24 <= 12'h8bc;
        src25 <= 12'hfaa;
        src26 <= 12'h84d;
        src27 <= 12'h98f;
        src28 <= 12'ha18;
        src29 <= 12'h1d9;
        src30 <= 12'h16f;
        src31 <= 12'hcc0;
        src32 <= 12'h315;
        src33 <= 12'hf7e;
        src34 <= 12'h6b1;
        src35 <= 12'h87f;
        src36 <= 12'h17e;
        src37 <= 12'h2d7;
        src38 <= 12'h1cf;
        src39 <= 12'h580;
        src40 <= 12'hfe1;
        src41 <= 12'had2;
        src42 <= 12'h945;
        src43 <= 12'h75a;
        src44 <= 12'h32d;
        src45 <= 12'h438;
        src46 <= 12'h69c;
        src47 <= 12'hce7;
        src48 <= 12'h3b4;
        src49 <= 12'hee7;
        src50 <= 12'hb1d;
        src51 <= 12'h785;
        src52 <= 12'h5b0;
        src53 <= 12'h2db;
        src54 <= 12'h5f8;
        src55 <= 12'h518;
        src56 <= 12'h26a;
        src57 <= 12'h6f3;
        src58 <= 12'h8de;
        src59 <= 12'hce1;
        src60 <= 12'h5ea;
        src61 <= 12'h847;
        src62 <= 12'h24d;
        src63 <= 12'ha61;
        src64 <= 12'ha93;
        src65 <= 12'hfb4;
        src66 <= 12'h72e;
        src67 <= 12'hede;
        src68 <= 12'h17d;
        src69 <= 12'h28c;
        src70 <= 12'h53d;
        src71 <= 12'h7ae;
        src72 <= 12'h4b8;
        src73 <= 12'hd9;
        src74 <= 12'heb5;
        src75 <= 12'hb24;
        src76 <= 12'haa0;
        src77 <= 12'h4bb;
        src78 <= 12'h227;
        src79 <= 12'hc84;
        src80 <= 12'ha98;
        src81 <= 12'h7b;
        src82 <= 12'h8d3;
        src83 <= 12'h661;
        src84 <= 12'h1d7;
        src85 <= 12'h9a3;
        src86 <= 12'h407;
        src87 <= 12'h1c7;
        src88 <= 12'h1d7;
        src89 <= 12'hfce;
        src90 <= 12'h962;
        src91 <= 12'h9b6;
        src92 <= 12'h6c9;
        src93 <= 12'h13f;
        src94 <= 12'hf9d;
        src95 <= 12'h642;
        src96 <= 12'h820;
        src97 <= 12'hb48;
        src98 <= 12'h9fe;
        src99 <= 12'h7ae;
        src100 <= 12'h90f;
        src101 <= 12'h3c4;
        src102 <= 12'h7ce;
        src103 <= 12'ha51;
        src104 <= 12'h235;
        src105 <= 12'hd64;
        src106 <= 12'h7e3;
        src107 <= 12'ha1a;
        src108 <= 12'h403;
        src109 <= 12'h4e1;
        src110 <= 12'hb35;
        src111 <= 12'ha60;
        src112 <= 12'hf5c;
        src113 <= 12'hbd5;
        src114 <= 12'h765;
        src115 <= 12'h46a;
        src116 <= 12'h1d;
        src117 <= 12'hccf;
        src118 <= 12'h359;
        src119 <= 12'h43b;
        src120 <= 12'hec3;
        src121 <= 12'h37a;
        src122 <= 12'h209;
        src123 <= 12'hadd;
        src124 <= 12'h73c;
        src125 <= 12'hb78;
        src126 <= 12'h458;
        src127 <= 12'hff7;
        src128 <= 12'hff7;
        src129 <= 12'h276;
        src130 <= 12'heeb;
        src131 <= 12'hcd;
        src132 <= 12'hdf4;
        src133 <= 12'hac;
        src134 <= 12'hb8;
        src135 <= 12'hd3e;
        src136 <= 12'hca9;
        src137 <= 12'h4a9;
        src138 <= 12'h6ed;
        src139 <= 12'he8d;
        src140 <= 12'h811;
        src141 <= 12'h5ab;
        src142 <= 12'hbf6;
        src143 <= 12'hcd6;
        src144 <= 12'hbb5;
        src145 <= 12'h2c3;
        src146 <= 12'he13;
        src147 <= 12'hf64;
        src148 <= 12'hb8e;
        src149 <= 12'h75d;
        src150 <= 12'hd5a;
        src151 <= 12'hb07;
        src152 <= 12'hb30;
        src153 <= 12'h10d;
        src154 <= 12'h281;
        src155 <= 12'hdc1;
        src156 <= 12'h9d0;
        src157 <= 12'he57;
        src158 <= 12'hef9;
        src159 <= 12'h52a;
        src160 <= 12'hf4c;
        src161 <= 12'h28;
        exp <= 20'h505f5;
        #1
        src0 <= 12'h944;
        src1 <= 12'hc02;
        src2 <= 12'h8;
        src3 <= 12'h583;
        src4 <= 12'hd57;
        src5 <= 12'hc17;
        src6 <= 12'h342;
        src7 <= 12'hc74;
        src8 <= 12'h30f;
        src9 <= 12'he99;
        src10 <= 12'h186;
        src11 <= 12'he52;
        src12 <= 12'h829;
        src13 <= 12'h889;
        src14 <= 12'h8b1;
        src15 <= 12'hdf5;
        src16 <= 12'hc46;
        src17 <= 12'hec2;
        src18 <= 12'hf61;
        src19 <= 12'h40d;
        src20 <= 12'hdf3;
        src21 <= 12'hd60;
        src22 <= 12'hcb1;
        src23 <= 12'hda0;
        src24 <= 12'h470;
        src25 <= 12'h635;
        src26 <= 12'hb8f;
        src27 <= 12'h8e8;
        src28 <= 12'hd47;
        src29 <= 12'hf6e;
        src30 <= 12'h30b;
        src31 <= 12'hee2;
        src32 <= 12'h2c7;
        src33 <= 12'hc32;
        src34 <= 12'h504;
        src35 <= 12'hebc;
        src36 <= 12'h8b4;
        src37 <= 12'h3fb;
        src38 <= 12'h3c9;
        src39 <= 12'hcd;
        src40 <= 12'ha86;
        src41 <= 12'h99a;
        src42 <= 12'h53b;
        src43 <= 12'h565;
        src44 <= 12'h33a;
        src45 <= 12'hc12;
        src46 <= 12'h4b6;
        src47 <= 12'heb4;
        src48 <= 12'h3bc;
        src49 <= 12'h7f8;
        src50 <= 12'hb3d;
        src51 <= 12'h1ca;
        src52 <= 12'hbcc;
        src53 <= 12'h2b;
        src54 <= 12'h7ee;
        src55 <= 12'h222;
        src56 <= 12'h559;
        src57 <= 12'h8bb;
        src58 <= 12'h28;
        src59 <= 12'h6e8;
        src60 <= 12'hccf;
        src61 <= 12'h51;
        src62 <= 12'hef8;
        src63 <= 12'h31f;
        src64 <= 12'h6c1;
        src65 <= 12'h217;
        src66 <= 12'h8ae;
        src67 <= 12'hb0f;
        src68 <= 12'h346;
        src69 <= 12'hffd;
        src70 <= 12'h154;
        src71 <= 12'h1c4;
        src72 <= 12'h40b;
        src73 <= 12'h993;
        src74 <= 12'hc1a;
        src75 <= 12'h50a;
        src76 <= 12'h677;
        src77 <= 12'hb21;
        src78 <= 12'h2e7;
        src79 <= 12'h2c3;
        src80 <= 12'hd4e;
        src81 <= 12'h7db;
        src82 <= 12'h46c;
        src83 <= 12'h64b;
        src84 <= 12'h783;
        src85 <= 12'hd8f;
        src86 <= 12'h9bc;
        src87 <= 12'h4a9;
        src88 <= 12'hd7d;
        src89 <= 12'h494;
        src90 <= 12'h3e9;
        src91 <= 12'he7e;
        src92 <= 12'hb36;
        src93 <= 12'h756;
        src94 <= 12'hf4;
        src95 <= 12'hd60;
        src96 <= 12'h939;
        src97 <= 12'h69e;
        src98 <= 12'hd20;
        src99 <= 12'h39a;
        src100 <= 12'h4e1;
        src101 <= 12'hce7;
        src102 <= 12'ha64;
        src103 <= 12'h993;
        src104 <= 12'h7d2;
        src105 <= 12'h346;
        src106 <= 12'hffc;
        src107 <= 12'h279;
        src108 <= 12'h398;
        src109 <= 12'h81b;
        src110 <= 12'hdfc;
        src111 <= 12'hf60;
        src112 <= 12'h9a8;
        src113 <= 12'h6e5;
        src114 <= 12'hb45;
        src115 <= 12'h404;
        src116 <= 12'h55a;
        src117 <= 12'h476;
        src118 <= 12'h343;
        src119 <= 12'h7d;
        src120 <= 12'h879;
        src121 <= 12'h618;
        src122 <= 12'he96;
        src123 <= 12'he78;
        src124 <= 12'h4f7;
        src125 <= 12'h3c0;
        src126 <= 12'h954;
        src127 <= 12'hbd0;
        src128 <= 12'h829;
        src129 <= 12'h28;
        src130 <= 12'h952;
        src131 <= 12'h9d2;
        src132 <= 12'hb65;
        src133 <= 12'haa7;
        src134 <= 12'h6de;
        src135 <= 12'h956;
        src136 <= 12'hc4d;
        src137 <= 12'h83e;
        src138 <= 12'h2d1;
        src139 <= 12'had7;
        src140 <= 12'hdd7;
        src141 <= 12'h227;
        src142 <= 12'h834;
        src143 <= 12'h920;
        src144 <= 12'h8e9;
        src145 <= 12'h25c;
        src146 <= 12'ha75;
        src147 <= 12'h59a;
        src148 <= 12'h3d7;
        src149 <= 12'hca9;
        src150 <= 12'h982;
        src151 <= 12'h5bc;
        src152 <= 12'h31f;
        src153 <= 12'h53d;
        src154 <= 12'h4b4;
        src155 <= 12'habe;
        src156 <= 12'ha03;
        src157 <= 12'ha9c;
        src158 <= 12'hd8b;
        src159 <= 12'h82;
        src160 <= 12'hca1;
        src161 <= 12'h317;
        exp <= 20'h51723;
        #1
        src0 <= 12'h6b9;
        src1 <= 12'h4d8;
        src2 <= 12'h8a8;
        src3 <= 12'hb5d;
        src4 <= 12'h1b1;
        src5 <= 12'hd78;
        src6 <= 12'h516;
        src7 <= 12'h285;
        src8 <= 12'hdac;
        src9 <= 12'hd9b;
        src10 <= 12'ha66;
        src11 <= 12'hd35;
        src12 <= 12'h90a;
        src13 <= 12'h99e;
        src14 <= 12'h263;
        src15 <= 12'h680;
        src16 <= 12'hea0;
        src17 <= 12'hc3d;
        src18 <= 12'hc59;
        src19 <= 12'he76;
        src20 <= 12'h26e;
        src21 <= 12'h86f;
        src22 <= 12'h3fc;
        src23 <= 12'h9fb;
        src24 <= 12'h7db;
        src25 <= 12'h266;
        src26 <= 12'h5c7;
        src27 <= 12'h7cf;
        src28 <= 12'h228;
        src29 <= 12'h423;
        src30 <= 12'hfbc;
        src31 <= 12'h4a8;
        src32 <= 12'h1e8;
        src33 <= 12'h2ff;
        src34 <= 12'ha58;
        src35 <= 12'h960;
        src36 <= 12'h649;
        src37 <= 12'h662;
        src38 <= 12'heaa;
        src39 <= 12'h935;
        src40 <= 12'hf90;
        src41 <= 12'he8b;
        src42 <= 12'h2ff;
        src43 <= 12'haa;
        src44 <= 12'h158;
        src45 <= 12'h80c;
        src46 <= 12'hb4c;
        src47 <= 12'h233;
        src48 <= 12'h9c7;
        src49 <= 12'h342;
        src50 <= 12'hbd1;
        src51 <= 12'hc55;
        src52 <= 12'he86;
        src53 <= 12'h4fc;
        src54 <= 12'h705;
        src55 <= 12'h1b2;
        src56 <= 12'hf87;
        src57 <= 12'h785;
        src58 <= 12'h873;
        src59 <= 12'h324;
        src60 <= 12'hfc3;
        src61 <= 12'h6f2;
        src62 <= 12'h6bb;
        src63 <= 12'h59d;
        src64 <= 12'h84;
        src65 <= 12'h486;
        src66 <= 12'h1f6;
        src67 <= 12'h37e;
        src68 <= 12'hdf0;
        src69 <= 12'he4a;
        src70 <= 12'he27;
        src71 <= 12'haf5;
        src72 <= 12'hb4d;
        src73 <= 12'hc59;
        src74 <= 12'h75b;
        src75 <= 12'h847;
        src76 <= 12'h520;
        src77 <= 12'he20;
        src78 <= 12'h8fb;
        src79 <= 12'hee0;
        src80 <= 12'h92e;
        src81 <= 12'h99f;
        src82 <= 12'ha23;
        src83 <= 12'hecb;
        src84 <= 12'h947;
        src85 <= 12'h8;
        src86 <= 12'h422;
        src87 <= 12'h937;
        src88 <= 12'h2cd;
        src89 <= 12'hb07;
        src90 <= 12'h457;
        src91 <= 12'h5cc;
        src92 <= 12'h41e;
        src93 <= 12'h111;
        src94 <= 12'h953;
        src95 <= 12'h80e;
        src96 <= 12'hcd9;
        src97 <= 12'hd2d;
        src98 <= 12'h1e6;
        src99 <= 12'he8d;
        src100 <= 12'ha6d;
        src101 <= 12'hf0b;
        src102 <= 12'h76d;
        src103 <= 12'hcfb;
        src104 <= 12'hb98;
        src105 <= 12'h2d0;
        src106 <= 12'h8d4;
        src107 <= 12'h6b0;
        src108 <= 12'hbaa;
        src109 <= 12'h1f1;
        src110 <= 12'hf05;
        src111 <= 12'h6a2;
        src112 <= 12'hfcc;
        src113 <= 12'h180;
        src114 <= 12'h85e;
        src115 <= 12'h7f1;
        src116 <= 12'h281;
        src117 <= 12'hfd0;
        src118 <= 12'h5c2;
        src119 <= 12'ha7;
        src120 <= 12'h72d;
        src121 <= 12'h698;
        src122 <= 12'h517;
        src123 <= 12'h9d0;
        src124 <= 12'h122;
        src125 <= 12'h34c;
        src126 <= 12'h2ad;
        src127 <= 12'h5f2;
        src128 <= 12'h392;
        src129 <= 12'haa9;
        src130 <= 12'he70;
        src131 <= 12'h57c;
        src132 <= 12'h1b5;
        src133 <= 12'h90e;
        src134 <= 12'hbd0;
        src135 <= 12'hb93;
        src136 <= 12'h328;
        src137 <= 12'h832;
        src138 <= 12'h17a;
        src139 <= 12'h4f0;
        src140 <= 12'h555;
        src141 <= 12'h7f1;
        src142 <= 12'hb70;
        src143 <= 12'h264;
        src144 <= 12'hc4e;
        src145 <= 12'he15;
        src146 <= 12'hbfc;
        src147 <= 12'hbbd;
        src148 <= 12'he14;
        src149 <= 12'ha8e;
        src150 <= 12'ha3c;
        src151 <= 12'h11d;
        src152 <= 12'h565;
        src153 <= 12'h276;
        src154 <= 12'h5a1;
        src155 <= 12'h570;
        src156 <= 12'h864;
        src157 <= 12'h37d;
        src158 <= 12'h9aa;
        src159 <= 12'hb05;
        src160 <= 12'hdc7;
        src161 <= 12'h4bc;
        exp <= 20'h510ac;
        #1
        src0 <= 12'h384;
        src1 <= 12'h4d6;
        src2 <= 12'h5ae;
        src3 <= 12'h881;
        src4 <= 12'h9c3;
        src5 <= 12'h53b;
        src6 <= 12'hf40;
        src7 <= 12'h3f5;
        src8 <= 12'hce1;
        src9 <= 12'hb1c;
        src10 <= 12'h26e;
        src11 <= 12'h6f4;
        src12 <= 12'h964;
        src13 <= 12'h526;
        src14 <= 12'h855;
        src15 <= 12'h167;
        src16 <= 12'h57b;
        src17 <= 12'h558;
        src18 <= 12'hd50;
        src19 <= 12'ha65;
        src20 <= 12'hfd8;
        src21 <= 12'h983;
        src22 <= 12'h266;
        src23 <= 12'h538;
        src24 <= 12'h61a;
        src25 <= 12'h9d2;
        src26 <= 12'h5a3;
        src27 <= 12'h409;
        src28 <= 12'h5ec;
        src29 <= 12'h13a;
        src30 <= 12'h246;
        src31 <= 12'h42c;
        src32 <= 12'h5f0;
        src33 <= 12'hb7a;
        src34 <= 12'ha58;
        src35 <= 12'h166;
        src36 <= 12'h1e0;
        src37 <= 12'h9d0;
        src38 <= 12'h2a7;
        src39 <= 12'h46a;
        src40 <= 12'h36c;
        src41 <= 12'h154;
        src42 <= 12'h31;
        src43 <= 12'h4d2;
        src44 <= 12'h3ea;
        src45 <= 12'h989;
        src46 <= 12'hf87;
        src47 <= 12'hb4;
        src48 <= 12'h541;
        src49 <= 12'h6e3;
        src50 <= 12'h91;
        src51 <= 12'h35d;
        src52 <= 12'h541;
        src53 <= 12'ha65;
        src54 <= 12'hd48;
        src55 <= 12'h280;
        src56 <= 12'h8a8;
        src57 <= 12'hcb7;
        src58 <= 12'h5b5;
        src59 <= 12'ha9c;
        src60 <= 12'h1fe;
        src61 <= 12'hcfc;
        src62 <= 12'hbd7;
        src63 <= 12'h86f;
        src64 <= 12'ha16;
        src65 <= 12'h697;
        src66 <= 12'hf12;
        src67 <= 12'h62f;
        src68 <= 12'h195;
        src69 <= 12'hbc0;
        src70 <= 12'h5b8;
        src71 <= 12'h476;
        src72 <= 12'h1cf;
        src73 <= 12'h377;
        src74 <= 12'h415;
        src75 <= 12'h8b1;
        src76 <= 12'hf51;
        src77 <= 12'h516;
        src78 <= 12'h312;
        src79 <= 12'h613;
        src80 <= 12'h761;
        src81 <= 12'hd5b;
        src82 <= 12'h9cc;
        src83 <= 12'h4f7;
        src84 <= 12'hf39;
        src85 <= 12'h2ae;
        src86 <= 12'h13;
        src87 <= 12'h205;
        src88 <= 12'h923;
        src89 <= 12'h5b2;
        src90 <= 12'h1df;
        src91 <= 12'hfaf;
        src92 <= 12'h6d2;
        src93 <= 12'h560;
        src94 <= 12'hf44;
        src95 <= 12'h565;
        src96 <= 12'h26;
        src97 <= 12'hd0f;
        src98 <= 12'h457;
        src99 <= 12'h783;
        src100 <= 12'hedd;
        src101 <= 12'hd6e;
        src102 <= 12'hbb7;
        src103 <= 12'h4bf;
        src104 <= 12'h3a5;
        src105 <= 12'h15;
        src106 <= 12'h881;
        src107 <= 12'h622;
        src108 <= 12'h74c;
        src109 <= 12'hd68;
        src110 <= 12'hd84;
        src111 <= 12'h6a8;
        src112 <= 12'h344;
        src113 <= 12'heed;
        src114 <= 12'he54;
        src115 <= 12'hbd3;
        src116 <= 12'hbab;
        src117 <= 12'h471;
        src118 <= 12'hc6d;
        src119 <= 12'h701;
        src120 <= 12'hd15;
        src121 <= 12'h22f;
        src122 <= 12'ha19;
        src123 <= 12'h1eb;
        src124 <= 12'h76e;
        src125 <= 12'hb05;
        src126 <= 12'hcef;
        src127 <= 12'ha69;
        src128 <= 12'h5fe;
        src129 <= 12'h8bb;
        src130 <= 12'hbf5;
        src131 <= 12'hb53;
        src132 <= 12'h7aa;
        src133 <= 12'hc56;
        src134 <= 12'ha45;
        src135 <= 12'h207;
        src136 <= 12'hff5;
        src137 <= 12'hc74;
        src138 <= 12'h5d3;
        src139 <= 12'h82c;
        src140 <= 12'ha14;
        src141 <= 12'h2d;
        src142 <= 12'h92c;
        src143 <= 12'hf2d;
        src144 <= 12'h313;
        src145 <= 12'hddc;
        src146 <= 12'h9cc;
        src147 <= 12'h5d;
        src148 <= 12'ha8a;
        src149 <= 12'h86e;
        src150 <= 12'h165;
        src151 <= 12'hb15;
        src152 <= 12'h2f2;
        src153 <= 12'h1d5;
        src154 <= 12'h69e;
        src155 <= 12'h66e;
        src156 <= 12'h518;
        src157 <= 12'h105;
        src158 <= 12'hcdd;
        src159 <= 12'hf1b;
        src160 <= 12'h663;
        src161 <= 12'hd89;
        exp <= 20'h4be50;
        #1
        src0 <= 12'h583;
        src1 <= 12'hda2;
        src2 <= 12'he5;
        src3 <= 12'hc23;
        src4 <= 12'h72b;
        src5 <= 12'h7d3;
        src6 <= 12'h5e;
        src7 <= 12'h336;
        src8 <= 12'hfe6;
        src9 <= 12'h5ce;
        src10 <= 12'h2e4;
        src11 <= 12'h58c;
        src12 <= 12'hc0c;
        src13 <= 12'h92b;
        src14 <= 12'h2e4;
        src15 <= 12'hb4e;
        src16 <= 12'h4c1;
        src17 <= 12'ha3c;
        src18 <= 12'h7fc;
        src19 <= 12'hacc;
        src20 <= 12'h5b0;
        src21 <= 12'h8f9;
        src22 <= 12'h717;
        src23 <= 12'h4e4;
        src24 <= 12'h299;
        src25 <= 12'hd16;
        src26 <= 12'h721;
        src27 <= 12'h5ac;
        src28 <= 12'hb21;
        src29 <= 12'h7ae;
        src30 <= 12'h75d;
        src31 <= 12'h239;
        src32 <= 12'hfc7;
        src33 <= 12'h165;
        src34 <= 12'hd73;
        src35 <= 12'hc4e;
        src36 <= 12'h11d;
        src37 <= 12'h2c1;
        src38 <= 12'h802;
        src39 <= 12'h33e;
        src40 <= 12'h8fa;
        src41 <= 12'h754;
        src42 <= 12'hb78;
        src43 <= 12'h8d0;
        src44 <= 12'hd21;
        src45 <= 12'h482;
        src46 <= 12'haaf;
        src47 <= 12'h837;
        src48 <= 12'h54c;
        src49 <= 12'hcb7;
        src50 <= 12'hb47;
        src51 <= 12'ha17;
        src52 <= 12'h351;
        src53 <= 12'hefb;
        src54 <= 12'h1bc;
        src55 <= 12'hd3;
        src56 <= 12'h1d8;
        src57 <= 12'h589;
        src58 <= 12'h591;
        src59 <= 12'ha21;
        src60 <= 12'h27f;
        src61 <= 12'h8f3;
        src62 <= 12'hacc;
        src63 <= 12'h5b;
        src64 <= 12'hd1a;
        src65 <= 12'h295;
        src66 <= 12'hba9;
        src67 <= 12'h5e1;
        src68 <= 12'hca7;
        src69 <= 12'h979;
        src70 <= 12'he83;
        src71 <= 12'hb10;
        src72 <= 12'h432;
        src73 <= 12'h6b6;
        src74 <= 12'h2ab;
        src75 <= 12'h473;
        src76 <= 12'h607;
        src77 <= 12'hffb;
        src78 <= 12'hc8e;
        src79 <= 12'hbd2;
        src80 <= 12'hf6c;
        src81 <= 12'h313;
        src82 <= 12'h8d;
        src83 <= 12'hc7b;
        src84 <= 12'hd1a;
        src85 <= 12'h82f;
        src86 <= 12'h386;
        src87 <= 12'h38a;
        src88 <= 12'h92f;
        src89 <= 12'hc1;
        src90 <= 12'h665;
        src91 <= 12'heea;
        src92 <= 12'hd0f;
        src93 <= 12'he54;
        src94 <= 12'h45f;
        src95 <= 12'hf11;
        src96 <= 12'h46c;
        src97 <= 12'h129;
        src98 <= 12'h879;
        src99 <= 12'h5c3;
        src100 <= 12'hfb2;
        src101 <= 12'hb84;
        src102 <= 12'hc54;
        src103 <= 12'h4ee;
        src104 <= 12'h3c3;
        src105 <= 12'h214;
        src106 <= 12'hc36;
        src107 <= 12'h89b;
        src108 <= 12'hb2a;
        src109 <= 12'he73;
        src110 <= 12'hf3f;
        src111 <= 12'h2d1;
        src112 <= 12'h3d1;
        src113 <= 12'h13;
        src114 <= 12'h8ec;
        src115 <= 12'hca2;
        src116 <= 12'hc17;
        src117 <= 12'hb16;
        src118 <= 12'h22a;
        src119 <= 12'he40;
        src120 <= 12'h484;
        src121 <= 12'hdb3;
        src122 <= 12'h329;
        src123 <= 12'h419;
        src124 <= 12'hcc4;
        src125 <= 12'hc9c;
        src126 <= 12'hf29;
        src127 <= 12'ha79;
        src128 <= 12'h7ec;
        src129 <= 12'h61b;
        src130 <= 12'h20f;
        src131 <= 12'h9e6;
        src132 <= 12'h19b;
        src133 <= 12'h323;
        src134 <= 12'h9cb;
        src135 <= 12'h75b;
        src136 <= 12'h462;
        src137 <= 12'hc26;
        src138 <= 12'heb6;
        src139 <= 12'hef4;
        src140 <= 12'hca4;
        src141 <= 12'h228;
        src142 <= 12'h9b2;
        src143 <= 12'he30;
        src144 <= 12'h653;
        src145 <= 12'he23;
        src146 <= 12'h8e8;
        src147 <= 12'h970;
        src148 <= 12'h48a;
        src149 <= 12'h622;
        src150 <= 12'h459;
        src151 <= 12'h18;
        src152 <= 12'h97;
        src153 <= 12'h283;
        src154 <= 12'hc72;
        src155 <= 12'h3d7;
        src156 <= 12'h43e;
        src157 <= 12'hb60;
        src158 <= 12'he43;
        src159 <= 12'h56e;
        src160 <= 12'h531;
        src161 <= 12'hff5;
        exp <= 20'h50c93;
        #1
        src0 <= 12'hb58;
        src1 <= 12'hb28;
        src2 <= 12'h9af;
        src3 <= 12'hd4c;
        src4 <= 12'h9f;
        src5 <= 12'hadc;
        src6 <= 12'h2ff;
        src7 <= 12'hc73;
        src8 <= 12'hcbe;
        src9 <= 12'h27d;
        src10 <= 12'h8fc;
        src11 <= 12'h383;
        src12 <= 12'hcc3;
        src13 <= 12'h5cd;
        src14 <= 12'h170;
        src15 <= 12'h350;
        src16 <= 12'ha7e;
        src17 <= 12'hafb;
        src18 <= 12'h785;
        src19 <= 12'h6b6;
        src20 <= 12'h1ff;
        src21 <= 12'h9c9;
        src22 <= 12'hb02;
        src23 <= 12'h14d;
        src24 <= 12'h5d8;
        src25 <= 12'he03;
        src26 <= 12'hf72;
        src27 <= 12'h883;
        src28 <= 12'hea;
        src29 <= 12'h112;
        src30 <= 12'h4c2;
        src31 <= 12'h3a1;
        src32 <= 12'h0;
        src33 <= 12'h5b4;
        src34 <= 12'h90d;
        src35 <= 12'h38c;
        src36 <= 12'h4c9;
        src37 <= 12'hc5b;
        src38 <= 12'h296;
        src39 <= 12'hca8;
        src40 <= 12'hc0d;
        src41 <= 12'h62;
        src42 <= 12'he60;
        src43 <= 12'h64c;
        src44 <= 12'h4ec;
        src45 <= 12'hfdc;
        src46 <= 12'hc77;
        src47 <= 12'h46f;
        src48 <= 12'h8fe;
        src49 <= 12'hb34;
        src50 <= 12'ha1;
        src51 <= 12'h63;
        src52 <= 12'ha21;
        src53 <= 12'h540;
        src54 <= 12'h2a0;
        src55 <= 12'hd98;
        src56 <= 12'he49;
        src57 <= 12'hd27;
        src58 <= 12'h884;
        src59 <= 12'hc51;
        src60 <= 12'h4cb;
        src61 <= 12'h697;
        src62 <= 12'h633;
        src63 <= 12'h14b;
        src64 <= 12'hfd5;
        src65 <= 12'hefa;
        src66 <= 12'h9bc;
        src67 <= 12'h90f;
        src68 <= 12'h670;
        src69 <= 12'hb2e;
        src70 <= 12'h769;
        src71 <= 12'h396;
        src72 <= 12'h40b;
        src73 <= 12'h70b;
        src74 <= 12'haff;
        src75 <= 12'h956;
        src76 <= 12'h899;
        src77 <= 12'h1c;
        src78 <= 12'h11;
        src79 <= 12'hba8;
        src80 <= 12'hae1;
        src81 <= 12'hf34;
        src82 <= 12'h76b;
        src83 <= 12'hf08;
        src84 <= 12'hb18;
        src85 <= 12'heb9;
        src86 <= 12'hc3;
        src87 <= 12'h579;
        src88 <= 12'hafe;
        src89 <= 12'h669;
        src90 <= 12'h974;
        src91 <= 12'h1a;
        src92 <= 12'h18e;
        src93 <= 12'hcca;
        src94 <= 12'h520;
        src95 <= 12'hf67;
        src96 <= 12'h66;
        src97 <= 12'h2c;
        src98 <= 12'h4b;
        src99 <= 12'h248;
        src100 <= 12'h5d2;
        src101 <= 12'hcb8;
        src102 <= 12'h7f;
        src103 <= 12'h848;
        src104 <= 12'h2eb;
        src105 <= 12'h58d;
        src106 <= 12'hbbe;
        src107 <= 12'h58b;
        src108 <= 12'h3a3;
        src109 <= 12'h8af;
        src110 <= 12'h300;
        src111 <= 12'he5d;
        src112 <= 12'h857;
        src113 <= 12'hfb6;
        src114 <= 12'hd48;
        src115 <= 12'hf1f;
        src116 <= 12'h21c;
        src117 <= 12'hb2d;
        src118 <= 12'he89;
        src119 <= 12'hea7;
        src120 <= 12'hae3;
        src121 <= 12'hc4b;
        src122 <= 12'hda2;
        src123 <= 12'hee;
        src124 <= 12'h9a8;
        src125 <= 12'h8ca;
        src126 <= 12'he93;
        src127 <= 12'h26d;
        src128 <= 12'hbb1;
        src129 <= 12'h8b4;
        src130 <= 12'h708;
        src131 <= 12'h3cb;
        src132 <= 12'h4c3;
        src133 <= 12'h878;
        src134 <= 12'hdb2;
        src135 <= 12'h956;
        src136 <= 12'h4a6;
        src137 <= 12'ha1b;
        src138 <= 12'hff6;
        src139 <= 12'h634;
        src140 <= 12'hbaf;
        src141 <= 12'had;
        src142 <= 12'hf15;
        src143 <= 12'h24b;
        src144 <= 12'heb;
        src145 <= 12'h673;
        src146 <= 12'hae3;
        src147 <= 12'h385;
        src148 <= 12'hd57;
        src149 <= 12'h950;
        src150 <= 12'h246;
        src151 <= 12'h6e8;
        src152 <= 12'h798;
        src153 <= 12'h964;
        src154 <= 12'h57;
        src155 <= 12'h985;
        src156 <= 12'h9ab;
        src157 <= 12'h849;
        src158 <= 12'h100;
        src159 <= 12'hd90;
        src160 <= 12'h905;
        src161 <= 12'hfed;
        exp <= 20'h4fd5f;
        #1
        src0 <= 12'h865;
        src1 <= 12'h9d;
        src2 <= 12'hd6e;
        src3 <= 12'h204;
        src4 <= 12'hf5b;
        src5 <= 12'h43d;
        src6 <= 12'h949;
        src7 <= 12'ha5d;
        src8 <= 12'h4c7;
        src9 <= 12'h99d;
        src10 <= 12'h79c;
        src11 <= 12'h4df;
        src12 <= 12'hec3;
        src13 <= 12'hf1;
        src14 <= 12'h460;
        src15 <= 12'hbb9;
        src16 <= 12'h778;
        src17 <= 12'hb47;
        src18 <= 12'h52;
        src19 <= 12'h7c5;
        src20 <= 12'h426;
        src21 <= 12'h96f;
        src22 <= 12'h235;
        src23 <= 12'hb8c;
        src24 <= 12'heaa;
        src25 <= 12'ha1a;
        src26 <= 12'h19f;
        src27 <= 12'h639;
        src28 <= 12'hb2b;
        src29 <= 12'h9bc;
        src30 <= 12'h30a;
        src31 <= 12'h1ab;
        src32 <= 12'h2ed;
        src33 <= 12'hd57;
        src34 <= 12'hf9f;
        src35 <= 12'hf62;
        src36 <= 12'hf4b;
        src37 <= 12'h98c;
        src38 <= 12'hf33;
        src39 <= 12'hbc8;
        src40 <= 12'h6ef;
        src41 <= 12'h713;
        src42 <= 12'h10e;
        src43 <= 12'h71e;
        src44 <= 12'he49;
        src45 <= 12'h38d;
        src46 <= 12'hdf0;
        src47 <= 12'hc9b;
        src48 <= 12'hbc9;
        src49 <= 12'hefa;
        src50 <= 12'h927;
        src51 <= 12'hc24;
        src52 <= 12'h89a;
        src53 <= 12'hc0f;
        src54 <= 12'hd3d;
        src55 <= 12'hb0e;
        src56 <= 12'hc80;
        src57 <= 12'ha69;
        src58 <= 12'h6d2;
        src59 <= 12'h61;
        src60 <= 12'h76d;
        src61 <= 12'he2c;
        src62 <= 12'h8e0;
        src63 <= 12'hba9;
        src64 <= 12'h385;
        src65 <= 12'habd;
        src66 <= 12'hba6;
        src67 <= 12'h9cf;
        src68 <= 12'ha4e;
        src69 <= 12'hec4;
        src70 <= 12'hffb;
        src71 <= 12'hf76;
        src72 <= 12'h7eb;
        src73 <= 12'hee8;
        src74 <= 12'ha81;
        src75 <= 12'ha15;
        src76 <= 12'h4da;
        src77 <= 12'h810;
        src78 <= 12'ha88;
        src79 <= 12'h2b5;
        src80 <= 12'h5a3;
        src81 <= 12'h5b3;
        src82 <= 12'hc7d;
        src83 <= 12'hfc3;
        src84 <= 12'h6ac;
        src85 <= 12'h572;
        src86 <= 12'h11d;
        src87 <= 12'h364;
        src88 <= 12'h33e;
        src89 <= 12'h21e;
        src90 <= 12'hc04;
        src91 <= 12'hf79;
        src92 <= 12'h26b;
        src93 <= 12'heda;
        src94 <= 12'hc0a;
        src95 <= 12'hcb6;
        src96 <= 12'h47f;
        src97 <= 12'h710;
        src98 <= 12'h921;
        src99 <= 12'hfdd;
        src100 <= 12'hc89;
        src101 <= 12'hd61;
        src102 <= 12'h483;
        src103 <= 12'hc3b;
        src104 <= 12'h956;
        src105 <= 12'hce7;
        src106 <= 12'h301;
        src107 <= 12'h8bf;
        src108 <= 12'he0;
        src109 <= 12'heb3;
        src110 <= 12'h6b6;
        src111 <= 12'h4cc;
        src112 <= 12'hb6;
        src113 <= 12'he20;
        src114 <= 12'h1af;
        src115 <= 12'haa4;
        src116 <= 12'h1ce;
        src117 <= 12'h4d;
        src118 <= 12'ha89;
        src119 <= 12'hb7f;
        src120 <= 12'h2e5;
        src121 <= 12'hbc9;
        src122 <= 12'hb2d;
        src123 <= 12'h4b0;
        src124 <= 12'h2dd;
        src125 <= 12'hb9a;
        src126 <= 12'h322;
        src127 <= 12'hc1;
        src128 <= 12'hc89;
        src129 <= 12'hc4c;
        src130 <= 12'h11;
        src131 <= 12'h2c8;
        src132 <= 12'he71;
        src133 <= 12'h878;
        src134 <= 12'hd50;
        src135 <= 12'hd16;
        src136 <= 12'hf53;
        src137 <= 12'hbf7;
        src138 <= 12'h9c2;
        src139 <= 12'hfca;
        src140 <= 12'hc0e;
        src141 <= 12'h7e9;
        src142 <= 12'h9f7;
        src143 <= 12'h59b;
        src144 <= 12'h460;
        src145 <= 12'h193;
        src146 <= 12'h9e6;
        src147 <= 12'h986;
        src148 <= 12'h996;
        src149 <= 12'h7ce;
        src150 <= 12'h641;
        src151 <= 12'he5;
        src152 <= 12'hc2c;
        src153 <= 12'h8e;
        src154 <= 12'hda;
        src155 <= 12'h263;
        src156 <= 12'h1c9;
        src157 <= 12'hbf7;
        src158 <= 12'h4fc;
        src159 <= 12'h76f;
        src160 <= 12'h576;
        src161 <= 12'h2e5;
        exp <= 20'h554bf;
        #1
        src0 <= 12'h519;
        src1 <= 12'h390;
        src2 <= 12'hadf;
        src3 <= 12'hdd;
        src4 <= 12'h613;
        src5 <= 12'h911;
        src6 <= 12'h348;
        src7 <= 12'h386;
        src8 <= 12'h9a5;
        src9 <= 12'h52f;
        src10 <= 12'h255;
        src11 <= 12'h4e;
        src12 <= 12'h89f;
        src13 <= 12'h3e5;
        src14 <= 12'h38f;
        src15 <= 12'h6b3;
        src16 <= 12'h416;
        src17 <= 12'hdb2;
        src18 <= 12'h8f6;
        src19 <= 12'h6f7;
        src20 <= 12'h465;
        src21 <= 12'ha65;
        src22 <= 12'h62;
        src23 <= 12'h454;
        src24 <= 12'hcf3;
        src25 <= 12'hd4e;
        src26 <= 12'hec1;
        src27 <= 12'h19a;
        src28 <= 12'h159;
        src29 <= 12'h22f;
        src30 <= 12'h40a;
        src31 <= 12'h6a2;
        src32 <= 12'h9af;
        src33 <= 12'h12b;
        src34 <= 12'hf9e;
        src35 <= 12'hf1e;
        src36 <= 12'hafb;
        src37 <= 12'hc96;
        src38 <= 12'hca3;
        src39 <= 12'h152;
        src40 <= 12'h9e1;
        src41 <= 12'hf41;
        src42 <= 12'h64e;
        src43 <= 12'h617;
        src44 <= 12'hcc2;
        src45 <= 12'h5ff;
        src46 <= 12'h1;
        src47 <= 12'h866;
        src48 <= 12'h66b;
        src49 <= 12'h6a;
        src50 <= 12'h25b;
        src51 <= 12'he1;
        src52 <= 12'hcff;
        src53 <= 12'h861;
        src54 <= 12'hece;
        src55 <= 12'h453;
        src56 <= 12'hf14;
        src57 <= 12'h466;
        src58 <= 12'h91b;
        src59 <= 12'hc5b;
        src60 <= 12'hf05;
        src61 <= 12'h6a;
        src62 <= 12'hf24;
        src63 <= 12'h3d3;
        src64 <= 12'h10;
        src65 <= 12'h2e5;
        src66 <= 12'hae;
        src67 <= 12'h1ae;
        src68 <= 12'h97b;
        src69 <= 12'ha90;
        src70 <= 12'h5dc;
        src71 <= 12'h803;
        src72 <= 12'he9f;
        src73 <= 12'h815;
        src74 <= 12'h64c;
        src75 <= 12'h64c;
        src76 <= 12'h2b1;
        src77 <= 12'hda2;
        src78 <= 12'h5d2;
        src79 <= 12'h69b;
        src80 <= 12'hc4a;
        src81 <= 12'hf61;
        src82 <= 12'he4c;
        src83 <= 12'h6af;
        src84 <= 12'hca1;
        src85 <= 12'ha01;
        src86 <= 12'ha46;
        src87 <= 12'hdd8;
        src88 <= 12'h74e;
        src89 <= 12'h29d;
        src90 <= 12'hc9f;
        src91 <= 12'h598;
        src92 <= 12'hfbf;
        src93 <= 12'hba2;
        src94 <= 12'h4ee;
        src95 <= 12'h698;
        src96 <= 12'hd31;
        src97 <= 12'h841;
        src98 <= 12'hdeb;
        src99 <= 12'h8d6;
        src100 <= 12'hdbf;
        src101 <= 12'h8ff;
        src102 <= 12'h584;
        src103 <= 12'hf08;
        src104 <= 12'h1bf;
        src105 <= 12'h453;
        src106 <= 12'h985;
        src107 <= 12'h9e7;
        src108 <= 12'hb7d;
        src109 <= 12'h752;
        src110 <= 12'he1a;
        src111 <= 12'h2a5;
        src112 <= 12'h28;
        src113 <= 12'h881;
        src114 <= 12'hb43;
        src115 <= 12'h432;
        src116 <= 12'h935;
        src117 <= 12'hb31;
        src118 <= 12'he95;
        src119 <= 12'h399;
        src120 <= 12'h668;
        src121 <= 12'h531;
        src122 <= 12'h76b;
        src123 <= 12'h2ce;
        src124 <= 12'h39b;
        src125 <= 12'h6f5;
        src126 <= 12'haeb;
        src127 <= 12'hbe1;
        src128 <= 12'he6d;
        src129 <= 12'he1c;
        src130 <= 12'h4ef;
        src131 <= 12'hfc8;
        src132 <= 12'hd7;
        src133 <= 12'h8cf;
        src134 <= 12'h77f;
        src135 <= 12'h191;
        src136 <= 12'h98e;
        src137 <= 12'ha71;
        src138 <= 12'h8f;
        src139 <= 12'hb94;
        src140 <= 12'hc2c;
        src141 <= 12'haf5;
        src142 <= 12'h1fd;
        src143 <= 12'h141;
        src144 <= 12'hb2c;
        src145 <= 12'h2d3;
        src146 <= 12'h31e;
        src147 <= 12'h328;
        src148 <= 12'h9d9;
        src149 <= 12'h826;
        src150 <= 12'hda3;
        src151 <= 12'ha04;
        src152 <= 12'he8d;
        src153 <= 12'hfe7;
        src154 <= 12'h87b;
        src155 <= 12'hc53;
        src156 <= 12'hc35;
        src157 <= 12'hf7d;
        src158 <= 12'hc82;
        src159 <= 12'h554;
        src160 <= 12'hb8d;
        src161 <= 12'h663;
        exp <= 20'h51187;
        #1
        src0 <= 12'h8c2;
        src1 <= 12'hc1f;
        src2 <= 12'hfc0;
        src3 <= 12'h1c5;
        src4 <= 12'h393;
        src5 <= 12'he35;
        src6 <= 12'hd4d;
        src7 <= 12'h75f;
        src8 <= 12'h49d;
        src9 <= 12'h9ae;
        src10 <= 12'h6f6;
        src11 <= 12'heaf;
        src12 <= 12'h270;
        src13 <= 12'h293;
        src14 <= 12'h2d7;
        src15 <= 12'h481;
        src16 <= 12'hb8c;
        src17 <= 12'h5a4;
        src18 <= 12'hf4;
        src19 <= 12'h8b3;
        src20 <= 12'h91e;
        src21 <= 12'h184;
        src22 <= 12'hf8f;
        src23 <= 12'h33e;
        src24 <= 12'h97c;
        src25 <= 12'hde5;
        src26 <= 12'hee3;
        src27 <= 12'h27a;
        src28 <= 12'h5cd;
        src29 <= 12'h17f;
        src30 <= 12'hfeb;
        src31 <= 12'h684;
        src32 <= 12'he46;
        src33 <= 12'h35c;
        src34 <= 12'h8d4;
        src35 <= 12'h5ce;
        src36 <= 12'hfaa;
        src37 <= 12'hae7;
        src38 <= 12'h6a5;
        src39 <= 12'h2da;
        src40 <= 12'hb72;
        src41 <= 12'h273;
        src42 <= 12'h733;
        src43 <= 12'h877;
        src44 <= 12'h9b8;
        src45 <= 12'hff6;
        src46 <= 12'h7b6;
        src47 <= 12'h538;
        src48 <= 12'h7bb;
        src49 <= 12'h9f3;
        src50 <= 12'h8ac;
        src51 <= 12'h188;
        src52 <= 12'h767;
        src53 <= 12'h104;
        src54 <= 12'hac6;
        src55 <= 12'ha2b;
        src56 <= 12'he8;
        src57 <= 12'ha0e;
        src58 <= 12'h182;
        src59 <= 12'h1ca;
        src60 <= 12'h204;
        src61 <= 12'h352;
        src62 <= 12'ha98;
        src63 <= 12'h7ff;
        src64 <= 12'h1f8;
        src65 <= 12'h609;
        src66 <= 12'h311;
        src67 <= 12'h58c;
        src68 <= 12'h8b1;
        src69 <= 12'h375;
        src70 <= 12'hc35;
        src71 <= 12'h392;
        src72 <= 12'h3cc;
        src73 <= 12'h380;
        src74 <= 12'h20e;
        src75 <= 12'hebc;
        src76 <= 12'h3e2;
        src77 <= 12'hc4;
        src78 <= 12'h61;
        src79 <= 12'hfac;
        src80 <= 12'he3b;
        src81 <= 12'h95f;
        src82 <= 12'h62;
        src83 <= 12'h8ca;
        src84 <= 12'h6dc;
        src85 <= 12'he24;
        src86 <= 12'h377;
        src87 <= 12'h46c;
        src88 <= 12'hd13;
        src89 <= 12'h4c0;
        src90 <= 12'hfc;
        src91 <= 12'ha7a;
        src92 <= 12'hb1d;
        src93 <= 12'h4ce;
        src94 <= 12'h351;
        src95 <= 12'hf6f;
        src96 <= 12'h57f;
        src97 <= 12'hd74;
        src98 <= 12'h5bd;
        src99 <= 12'h429;
        src100 <= 12'h18c;
        src101 <= 12'hed2;
        src102 <= 12'hbc0;
        src103 <= 12'h260;
        src104 <= 12'h237;
        src105 <= 12'h61c;
        src106 <= 12'h6b6;
        src107 <= 12'h188;
        src108 <= 12'ha55;
        src109 <= 12'h61c;
        src110 <= 12'hf6f;
        src111 <= 12'hc46;
        src112 <= 12'h5e3;
        src113 <= 12'h1ae;
        src114 <= 12'h610;
        src115 <= 12'h20a;
        src116 <= 12'hc1d;
        src117 <= 12'h91;
        src118 <= 12'h1a7;
        src119 <= 12'h149;
        src120 <= 12'hfb5;
        src121 <= 12'h282;
        src122 <= 12'h434;
        src123 <= 12'h40d;
        src124 <= 12'he69;
        src125 <= 12'hccf;
        src126 <= 12'h657;
        src127 <= 12'h620;
        src128 <= 12'h45d;
        src129 <= 12'h2d0;
        src130 <= 12'hfd5;
        src131 <= 12'hd77;
        src132 <= 12'h97d;
        src133 <= 12'h5b6;
        src134 <= 12'h192;
        src135 <= 12'h1d1;
        src136 <= 12'he38;
        src137 <= 12'h9f6;
        src138 <= 12'h5c0;
        src139 <= 12'hae9;
        src140 <= 12'h837;
        src141 <= 12'hbc7;
        src142 <= 12'h76d;
        src143 <= 12'hcce;
        src144 <= 12'h428;
        src145 <= 12'h4d2;
        src146 <= 12'h350;
        src147 <= 12'h2f6;
        src148 <= 12'h30b;
        src149 <= 12'h47e;
        src150 <= 12'hdc1;
        src151 <= 12'hea;
        src152 <= 12'hcd8;
        src153 <= 12'h93b;
        src154 <= 12'h454;
        src155 <= 12'ha1e;
        src156 <= 12'h7e9;
        src157 <= 12'hb68;
        src158 <= 12'h496;
        src159 <= 12'h3b1;
        src160 <= 12'he09;
        src161 <= 12'h280;
        exp <= 20'h49278;
        #1
        src0 <= 12'h882;
        src1 <= 12'h2ab;
        src2 <= 12'h7ae;
        src3 <= 12'hbb5;
        src4 <= 12'h56a;
        src5 <= 12'h111;
        src6 <= 12'h94e;
        src7 <= 12'h691;
        src8 <= 12'heb;
        src9 <= 12'hd33;
        src10 <= 12'he1;
        src11 <= 12'hd55;
        src12 <= 12'hfaf;
        src13 <= 12'h4be;
        src14 <= 12'h326;
        src15 <= 12'hf00;
        src16 <= 12'h9c5;
        src17 <= 12'h54a;
        src18 <= 12'hbad;
        src19 <= 12'h630;
        src20 <= 12'hc22;
        src21 <= 12'hdb2;
        src22 <= 12'h186;
        src23 <= 12'h86d;
        src24 <= 12'h9ee;
        src25 <= 12'h358;
        src26 <= 12'hf5f;
        src27 <= 12'h4d3;
        src28 <= 12'hda3;
        src29 <= 12'hda2;
        src30 <= 12'h86a;
        src31 <= 12'h6e;
        src32 <= 12'h9b9;
        src33 <= 12'h355;
        src34 <= 12'h8bf;
        src35 <= 12'h548;
        src36 <= 12'h4a8;
        src37 <= 12'h8d4;
        src38 <= 12'h7db;
        src39 <= 12'haee;
        src40 <= 12'hab4;
        src41 <= 12'hd1a;
        src42 <= 12'h2d9;
        src43 <= 12'hfc6;
        src44 <= 12'h45c;
        src45 <= 12'hf9e;
        src46 <= 12'h596;
        src47 <= 12'he38;
        src48 <= 12'hd45;
        src49 <= 12'hcf8;
        src50 <= 12'hc9d;
        src51 <= 12'hc8d;
        src52 <= 12'h35;
        src53 <= 12'h55;
        src54 <= 12'h4d2;
        src55 <= 12'h17a;
        src56 <= 12'h898;
        src57 <= 12'ha4c;
        src58 <= 12'h2e;
        src59 <= 12'h44;
        src60 <= 12'hc47;
        src61 <= 12'h519;
        src62 <= 12'hfa;
        src63 <= 12'hb93;
        src64 <= 12'h2ad;
        src65 <= 12'hcc7;
        src66 <= 12'h716;
        src67 <= 12'h8cb;
        src68 <= 12'hfad;
        src69 <= 12'h10a;
        src70 <= 12'h846;
        src71 <= 12'h18a;
        src72 <= 12'h864;
        src73 <= 12'hab4;
        src74 <= 12'h5e7;
        src75 <= 12'h74f;
        src76 <= 12'h557;
        src77 <= 12'h102;
        src78 <= 12'hbd;
        src79 <= 12'ha5b;
        src80 <= 12'hc0e;
        src81 <= 12'h24d;
        src82 <= 12'h181;
        src83 <= 12'h852;
        src84 <= 12'h560;
        src85 <= 12'h5cf;
        src86 <= 12'h35d;
        src87 <= 12'hc35;
        src88 <= 12'h43e;
        src89 <= 12'h86d;
        src90 <= 12'h222;
        src91 <= 12'h885;
        src92 <= 12'h187;
        src93 <= 12'h60e;
        src94 <= 12'h1da;
        src95 <= 12'h43b;
        src96 <= 12'hb7d;
        src97 <= 12'hfc8;
        src98 <= 12'h2cd;
        src99 <= 12'hc37;
        src100 <= 12'h653;
        src101 <= 12'h592;
        src102 <= 12'hf9f;
        src103 <= 12'he78;
        src104 <= 12'hccd;
        src105 <= 12'h668;
        src106 <= 12'h661;
        src107 <= 12'h8cb;
        src108 <= 12'h19f;
        src109 <= 12'h2d;
        src110 <= 12'hf1e;
        src111 <= 12'h171;
        src112 <= 12'h643;
        src113 <= 12'ha1c;
        src114 <= 12'hd3d;
        src115 <= 12'hd43;
        src116 <= 12'h6e7;
        src117 <= 12'hafe;
        src118 <= 12'hedb;
        src119 <= 12'h167;
        src120 <= 12'h46;
        src121 <= 12'h9e2;
        src122 <= 12'he3;
        src123 <= 12'h17f;
        src124 <= 12'h11a;
        src125 <= 12'h7be;
        src126 <= 12'h92e;
        src127 <= 12'hdf3;
        src128 <= 12'hb1e;
        src129 <= 12'h85e;
        src130 <= 12'hed6;
        src131 <= 12'hed2;
        src132 <= 12'h260;
        src133 <= 12'hcdc;
        src134 <= 12'h403;
        src135 <= 12'h868;
        src136 <= 12'hfdd;
        src137 <= 12'hbe2;
        src138 <= 12'h57e;
        src139 <= 12'ha0f;
        src140 <= 12'hff7;
        src141 <= 12'h97b;
        src142 <= 12'ha02;
        src143 <= 12'h55b;
        src144 <= 12'hb10;
        src145 <= 12'hd89;
        src146 <= 12'hb2d;
        src147 <= 12'h668;
        src148 <= 12'h90e;
        src149 <= 12'h251;
        src150 <= 12'h7e5;
        src151 <= 12'hdf4;
        src152 <= 12'h8fe;
        src153 <= 12'he53;
        src154 <= 12'h2e2;
        src155 <= 12'h25c;
        src156 <= 12'hece;
        src157 <= 12'hdf5;
        src158 <= 12'h4e0;
        src159 <= 12'hf6a;
        src160 <= 12'h804;
        src161 <= 12'h60f;
        exp <= 20'h50933;
        #1
        src0 <= 12'h27e;
        src1 <= 12'hfe7;
        src2 <= 12'h48f;
        src3 <= 12'hf78;
        src4 <= 12'h129;
        src5 <= 12'h2a8;
        src6 <= 12'hca0;
        src7 <= 12'h97b;
        src8 <= 12'h8bc;
        src9 <= 12'h884;
        src10 <= 12'h456;
        src11 <= 12'h8e8;
        src12 <= 12'h1f1;
        src13 <= 12'h19e;
        src14 <= 12'hc42;
        src15 <= 12'h37f;
        src16 <= 12'hef9;
        src17 <= 12'hc35;
        src18 <= 12'hbc4;
        src19 <= 12'hfca;
        src20 <= 12'hb6e;
        src21 <= 12'h530;
        src22 <= 12'h7f1;
        src23 <= 12'h20e;
        src24 <= 12'hf9e;
        src25 <= 12'hc60;
        src26 <= 12'h9f7;
        src27 <= 12'h97c;
        src28 <= 12'h524;
        src29 <= 12'h408;
        src30 <= 12'h2e6;
        src31 <= 12'hcf;
        src32 <= 12'ha8b;
        src33 <= 12'h483;
        src34 <= 12'h91;
        src35 <= 12'hbbb;
        src36 <= 12'heb1;
        src37 <= 12'h8c2;
        src38 <= 12'h72;
        src39 <= 12'h40c;
        src40 <= 12'ha3a;
        src41 <= 12'had2;
        src42 <= 12'hba3;
        src43 <= 12'h755;
        src44 <= 12'h47e;
        src45 <= 12'h72d;
        src46 <= 12'h2c4;
        src47 <= 12'h6da;
        src48 <= 12'h214;
        src49 <= 12'hfb1;
        src50 <= 12'hbad;
        src51 <= 12'h404;
        src52 <= 12'he5c;
        src53 <= 12'h1bc;
        src54 <= 12'hd3e;
        src55 <= 12'h68f;
        src56 <= 12'h776;
        src57 <= 12'he43;
        src58 <= 12'hc03;
        src59 <= 12'hf6f;
        src60 <= 12'hedf;
        src61 <= 12'hfb2;
        src62 <= 12'hc44;
        src63 <= 12'h984;
        src64 <= 12'h125;
        src65 <= 12'h1f0;
        src66 <= 12'h2de;
        src67 <= 12'ha0;
        src68 <= 12'h55;
        src69 <= 12'hce8;
        src70 <= 12'hf78;
        src71 <= 12'h48b;
        src72 <= 12'he76;
        src73 <= 12'hf2f;
        src74 <= 12'h65a;
        src75 <= 12'h24e;
        src76 <= 12'hc04;
        src77 <= 12'hd5e;
        src78 <= 12'h17a;
        src79 <= 12'ha05;
        src80 <= 12'h39e;
        src81 <= 12'h493;
        src82 <= 12'h601;
        src83 <= 12'h6b4;
        src84 <= 12'hc4f;
        src85 <= 12'h19;
        src86 <= 12'h3a1;
        src87 <= 12'h77f;
        src88 <= 12'h50b;
        src89 <= 12'h56d;
        src90 <= 12'h341;
        src91 <= 12'h567;
        src92 <= 12'hf4;
        src93 <= 12'h90e;
        src94 <= 12'h451;
        src95 <= 12'hc03;
        src96 <= 12'h5ed;
        src97 <= 12'hc3e;
        src98 <= 12'h7bb;
        src99 <= 12'h6cd;
        src100 <= 12'hd98;
        src101 <= 12'h435;
        src102 <= 12'h4f1;
        src103 <= 12'h66f;
        src104 <= 12'hf90;
        src105 <= 12'h789;
        src106 <= 12'hf1a;
        src107 <= 12'h9a0;
        src108 <= 12'hc03;
        src109 <= 12'h3a7;
        src110 <= 12'h6e7;
        src111 <= 12'h152;
        src112 <= 12'hb13;
        src113 <= 12'h653;
        src114 <= 12'h4eb;
        src115 <= 12'he32;
        src116 <= 12'h7a7;
        src117 <= 12'h331;
        src118 <= 12'hd9;
        src119 <= 12'h56a;
        src120 <= 12'h1;
        src121 <= 12'h3e3;
        src122 <= 12'hd8e;
        src123 <= 12'hf00;
        src124 <= 12'hb5d;
        src125 <= 12'h3d0;
        src126 <= 12'haf0;
        src127 <= 12'h6cd;
        src128 <= 12'he31;
        src129 <= 12'h5fa;
        src130 <= 12'h712;
        src131 <= 12'hdb4;
        src132 <= 12'h917;
        src133 <= 12'h3e1;
        src134 <= 12'h13c;
        src135 <= 12'h2a1;
        src136 <= 12'hb44;
        src137 <= 12'h84c;
        src138 <= 12'h136;
        src139 <= 12'hf61;
        src140 <= 12'hdde;
        src141 <= 12'heaf;
        src142 <= 12'h2f9;
        src143 <= 12'h363;
        src144 <= 12'h951;
        src145 <= 12'h1b6;
        src146 <= 12'hdd3;
        src147 <= 12'h82;
        src148 <= 12'h5dc;
        src149 <= 12'h6e9;
        src150 <= 12'h7a1;
        src151 <= 12'h149;
        src152 <= 12'h329;
        src153 <= 12'h538;
        src154 <= 12'h66;
        src155 <= 12'h88e;
        src156 <= 12'h914;
        src157 <= 12'h314;
        src158 <= 12'h7e6;
        src159 <= 12'hba4;
        src160 <= 12'hd5f;
        src161 <= 12'hf5f;
        exp <= 20'h4e663;
        #1
        src0 <= 12'h6d0;
        src1 <= 12'h389;
        src2 <= 12'h79a;
        src3 <= 12'h763;
        src4 <= 12'h10f;
        src5 <= 12'h218;
        src6 <= 12'h616;
        src7 <= 12'h904;
        src8 <= 12'he20;
        src9 <= 12'h109;
        src10 <= 12'h97b;
        src11 <= 12'hdd2;
        src12 <= 12'h668;
        src13 <= 12'h250;
        src14 <= 12'hf83;
        src15 <= 12'haf0;
        src16 <= 12'hcdd;
        src17 <= 12'h999;
        src18 <= 12'hc0d;
        src19 <= 12'hff;
        src20 <= 12'h5d8;
        src21 <= 12'h856;
        src22 <= 12'hb5b;
        src23 <= 12'h701;
        src24 <= 12'h559;
        src25 <= 12'h308;
        src26 <= 12'h1ed;
        src27 <= 12'h842;
        src28 <= 12'h9e;
        src29 <= 12'he7c;
        src30 <= 12'hc51;
        src31 <= 12'hab8;
        src32 <= 12'hb87;
        src33 <= 12'h4da;
        src34 <= 12'h5a8;
        src35 <= 12'h370;
        src36 <= 12'h118;
        src37 <= 12'h441;
        src38 <= 12'h39f;
        src39 <= 12'hd73;
        src40 <= 12'hd62;
        src41 <= 12'hcae;
        src42 <= 12'h3c0;
        src43 <= 12'ha63;
        src44 <= 12'h21a;
        src45 <= 12'h223;
        src46 <= 12'hc2b;
        src47 <= 12'he82;
        src48 <= 12'h8ff;
        src49 <= 12'h633;
        src50 <= 12'haff;
        src51 <= 12'h462;
        src52 <= 12'hb5a;
        src53 <= 12'h256;
        src54 <= 12'h2e2;
        src55 <= 12'h74a;
        src56 <= 12'hdeb;
        src57 <= 12'h45;
        src58 <= 12'h836;
        src59 <= 12'h4c4;
        src60 <= 12'h814;
        src61 <= 12'hbee;
        src62 <= 12'hf0e;
        src63 <= 12'hbb5;
        src64 <= 12'he8f;
        src65 <= 12'h5b2;
        src66 <= 12'he34;
        src67 <= 12'h722;
        src68 <= 12'h4bf;
        src69 <= 12'hb53;
        src70 <= 12'h9aa;
        src71 <= 12'hb80;
        src72 <= 12'h89;
        src73 <= 12'h80d;
        src74 <= 12'h76c;
        src75 <= 12'h114;
        src76 <= 12'h1be;
        src77 <= 12'h7d;
        src78 <= 12'h124;
        src79 <= 12'hab9;
        src80 <= 12'h9f2;
        src81 <= 12'h2f1;
        src82 <= 12'hdf5;
        src83 <= 12'h424;
        src84 <= 12'hbbe;
        src85 <= 12'h88d;
        src86 <= 12'hcdb;
        src87 <= 12'hf3e;
        src88 <= 12'hcc4;
        src89 <= 12'h63f;
        src90 <= 12'h19d;
        src91 <= 12'h876;
        src92 <= 12'h872;
        src93 <= 12'h787;
        src94 <= 12'h7b7;
        src95 <= 12'hdf1;
        src96 <= 12'h89b;
        src97 <= 12'h177;
        src98 <= 12'h3a0;
        src99 <= 12'h3b7;
        src100 <= 12'h764;
        src101 <= 12'h68c;
        src102 <= 12'ha4c;
        src103 <= 12'h215;
        src104 <= 12'h13b;
        src105 <= 12'h500;
        src106 <= 12'h448;
        src107 <= 12'h9d9;
        src108 <= 12'h21b;
        src109 <= 12'h6f4;
        src110 <= 12'h632;
        src111 <= 12'hb4b;
        src112 <= 12'hb71;
        src113 <= 12'h4ca;
        src114 <= 12'h46a;
        src115 <= 12'h6bf;
        src116 <= 12'h5a4;
        src117 <= 12'h3f5;
        src118 <= 12'h8dd;
        src119 <= 12'he0e;
        src120 <= 12'h474;
        src121 <= 12'h777;
        src122 <= 12'h608;
        src123 <= 12'hf54;
        src124 <= 12'hd23;
        src125 <= 12'hc8b;
        src126 <= 12'hae5;
        src127 <= 12'hecb;
        src128 <= 12'h9e9;
        src129 <= 12'hca4;
        src130 <= 12'h1a2;
        src131 <= 12'h291;
        src132 <= 12'h97e;
        src133 <= 12'hca6;
        src134 <= 12'h129;
        src135 <= 12'hd12;
        src136 <= 12'h65d;
        src137 <= 12'hec9;
        src138 <= 12'hc5c;
        src139 <= 12'h9c8;
        src140 <= 12'h1dc;
        src141 <= 12'h4cb;
        src142 <= 12'hb8f;
        src143 <= 12'hd1f;
        src144 <= 12'h95d;
        src145 <= 12'h204;
        src146 <= 12'h615;
        src147 <= 12'h7a2;
        src148 <= 12'h882;
        src149 <= 12'h80;
        src150 <= 12'h169;
        src151 <= 12'h86c;
        src152 <= 12'h45b;
        src153 <= 12'h9f2;
        src154 <= 12'h647;
        src155 <= 12'hb68;
        src156 <= 12'hb3e;
        src157 <= 12'h8f0;
        src158 <= 12'ha09;
        src159 <= 12'h52b;
        src160 <= 12'he22;
        src161 <= 12'h48f;
        exp <= 20'h4e059;
        #1
        src0 <= 12'hee5;
        src1 <= 12'h6b;
        src2 <= 12'hac7;
        src3 <= 12'h388;
        src4 <= 12'hb29;
        src5 <= 12'hbb7;
        src6 <= 12'h3ee;
        src7 <= 12'h7ce;
        src8 <= 12'h36;
        src9 <= 12'h769;
        src10 <= 12'hed5;
        src11 <= 12'hc86;
        src12 <= 12'h8c6;
        src13 <= 12'h421;
        src14 <= 12'h906;
        src15 <= 12'h8dc;
        src16 <= 12'hf67;
        src17 <= 12'ha71;
        src18 <= 12'ha51;
        src19 <= 12'hd8a;
        src20 <= 12'h6be;
        src21 <= 12'h3f6;
        src22 <= 12'h10b;
        src23 <= 12'h3ec;
        src24 <= 12'hc5f;
        src25 <= 12'h6be;
        src26 <= 12'h190;
        src27 <= 12'he98;
        src28 <= 12'h6d3;
        src29 <= 12'hd9b;
        src30 <= 12'h6fc;
        src31 <= 12'hd9a;
        src32 <= 12'h426;
        src33 <= 12'hf7;
        src34 <= 12'hdef;
        src35 <= 12'hd1e;
        src36 <= 12'h3e6;
        src37 <= 12'hd3;
        src38 <= 12'h2;
        src39 <= 12'ha07;
        src40 <= 12'h32a;
        src41 <= 12'h9ae;
        src42 <= 12'h31;
        src43 <= 12'h161;
        src44 <= 12'h28a;
        src45 <= 12'h2e8;
        src46 <= 12'h692;
        src47 <= 12'h49;
        src48 <= 12'hf68;
        src49 <= 12'h7e9;
        src50 <= 12'h77a;
        src51 <= 12'h21a;
        src52 <= 12'h181;
        src53 <= 12'haef;
        src54 <= 12'h58a;
        src55 <= 12'hc53;
        src56 <= 12'hbb;
        src57 <= 12'hede;
        src58 <= 12'h521;
        src59 <= 12'h7d;
        src60 <= 12'h781;
        src61 <= 12'he1a;
        src62 <= 12'h76e;
        src63 <= 12'hac7;
        src64 <= 12'hd45;
        src65 <= 12'h9e4;
        src66 <= 12'h6a9;
        src67 <= 12'h310;
        src68 <= 12'hd27;
        src69 <= 12'h3aa;
        src70 <= 12'hdbb;
        src71 <= 12'hbbe;
        src72 <= 12'h4c4;
        src73 <= 12'h77e;
        src74 <= 12'ha91;
        src75 <= 12'h86c;
        src76 <= 12'h90f;
        src77 <= 12'hc9d;
        src78 <= 12'h1d7;
        src79 <= 12'hbaa;
        src80 <= 12'ha25;
        src81 <= 12'hba3;
        src82 <= 12'h309;
        src83 <= 12'hece;
        src84 <= 12'h5d3;
        src85 <= 12'h947;
        src86 <= 12'hb8a;
        src87 <= 12'h509;
        src88 <= 12'h93a;
        src89 <= 12'h2fa;
        src90 <= 12'hd1d;
        src91 <= 12'hf13;
        src92 <= 12'ha52;
        src93 <= 12'hf0a;
        src94 <= 12'hdd4;
        src95 <= 12'hf24;
        src96 <= 12'hbf4;
        src97 <= 12'hc21;
        src98 <= 12'h159;
        src99 <= 12'h440;
        src100 <= 12'h2b;
        src101 <= 12'hf5b;
        src102 <= 12'h79f;
        src103 <= 12'h72c;
        src104 <= 12'h792;
        src105 <= 12'hd01;
        src106 <= 12'hb57;
        src107 <= 12'h3ec;
        src108 <= 12'h7d1;
        src109 <= 12'he83;
        src110 <= 12'h9ac;
        src111 <= 12'hc00;
        src112 <= 12'ha7e;
        src113 <= 12'h3ba;
        src114 <= 12'h513;
        src115 <= 12'h7b7;
        src116 <= 12'ha66;
        src117 <= 12'h37c;
        src118 <= 12'h9e0;
        src119 <= 12'h795;
        src120 <= 12'hde7;
        src121 <= 12'h57f;
        src122 <= 12'hb2b;
        src123 <= 12'h2d6;
        src124 <= 12'h4be;
        src125 <= 12'h394;
        src126 <= 12'h2ab;
        src127 <= 12'h31a;
        src128 <= 12'h93a;
        src129 <= 12'hc7;
        src130 <= 12'h44a;
        src131 <= 12'hcee;
        src132 <= 12'h7a4;
        src133 <= 12'hfab;
        src134 <= 12'ha61;
        src135 <= 12'h179;
        src136 <= 12'h905;
        src137 <= 12'he3b;
        src138 <= 12'hc6f;
        src139 <= 12'h4cd;
        src140 <= 12'h465;
        src141 <= 12'h5ca;
        src142 <= 12'hff2;
        src143 <= 12'hc2c;
        src144 <= 12'hdf1;
        src145 <= 12'h3ca;
        src146 <= 12'h289;
        src147 <= 12'hbd3;
        src148 <= 12'hb57;
        src149 <= 12'h80f;
        src150 <= 12'h480;
        src151 <= 12'hf00;
        src152 <= 12'h34c;
        src153 <= 12'he0c;
        src154 <= 12'he02;
        src155 <= 12'hcad;
        src156 <= 12'h51f;
        src157 <= 12'ha9d;
        src158 <= 12'hff0;
        src159 <= 12'h633;
        src160 <= 12'h758;
        src161 <= 12'hfe;
        exp <= 20'h52d2d;
        #1
        src0 <= 12'h9e0;
        src1 <= 12'hd88;
        src2 <= 12'hea5;
        src3 <= 12'hb10;
        src4 <= 12'h5cf;
        src5 <= 12'h4e3;
        src6 <= 12'h568;
        src7 <= 12'h9d8;
        src8 <= 12'h370;
        src9 <= 12'h208;
        src10 <= 12'hec9;
        src11 <= 12'hb70;
        src12 <= 12'h3a0;
        src13 <= 12'h7b5;
        src14 <= 12'he5f;
        src15 <= 12'ha;
        src16 <= 12'hfa3;
        src17 <= 12'he95;
        src18 <= 12'h97b;
        src19 <= 12'hca3;
        src20 <= 12'h308;
        src21 <= 12'h828;
        src22 <= 12'h198;
        src23 <= 12'hd83;
        src24 <= 12'h829;
        src25 <= 12'h96d;
        src26 <= 12'h61a;
        src27 <= 12'hd13;
        src28 <= 12'h708;
        src29 <= 12'h1ce;
        src30 <= 12'hb31;
        src31 <= 12'hea0;
        src32 <= 12'hd4b;
        src33 <= 12'h753;
        src34 <= 12'h113;
        src35 <= 12'h6df;
        src36 <= 12'h59d;
        src37 <= 12'h54b;
        src38 <= 12'hbfe;
        src39 <= 12'h7a9;
        src40 <= 12'h72;
        src41 <= 12'hc78;
        src42 <= 12'hd0f;
        src43 <= 12'hab;
        src44 <= 12'h750;
        src45 <= 12'hc2d;
        src46 <= 12'hcae;
        src47 <= 12'h372;
        src48 <= 12'hf63;
        src49 <= 12'hcf5;
        src50 <= 12'h876;
        src51 <= 12'hdad;
        src52 <= 12'hf7b;
        src53 <= 12'h23b;
        src54 <= 12'ha5f;
        src55 <= 12'h55a;
        src56 <= 12'h6a4;
        src57 <= 12'h330;
        src58 <= 12'hd4f;
        src59 <= 12'hfca;
        src60 <= 12'h1f3;
        src61 <= 12'h4ed;
        src62 <= 12'h72;
        src63 <= 12'h85f;
        src64 <= 12'h666;
        src65 <= 12'h116;
        src66 <= 12'h5ed;
        src67 <= 12'h50f;
        src68 <= 12'hf8c;
        src69 <= 12'h5ee;
        src70 <= 12'h998;
        src71 <= 12'hcb7;
        src72 <= 12'h532;
        src73 <= 12'hf7b;
        src74 <= 12'hb6b;
        src75 <= 12'h9ee;
        src76 <= 12'hc77;
        src77 <= 12'he8b;
        src78 <= 12'haef;
        src79 <= 12'hf8b;
        src80 <= 12'h96d;
        src81 <= 12'ha95;
        src82 <= 12'h9a2;
        src83 <= 12'h29d;
        src84 <= 12'h753;
        src85 <= 12'hb33;
        src86 <= 12'hcc1;
        src87 <= 12'hbb7;
        src88 <= 12'h506;
        src89 <= 12'he53;
        src90 <= 12'h861;
        src91 <= 12'h6eb;
        src92 <= 12'h898;
        src93 <= 12'h8da;
        src94 <= 12'hf04;
        src95 <= 12'hffd;
        src96 <= 12'h32f;
        src97 <= 12'haf4;
        src98 <= 12'hf5e;
        src99 <= 12'ha80;
        src100 <= 12'h357;
        src101 <= 12'ha0f;
        src102 <= 12'hab4;
        src103 <= 12'heb;
        src104 <= 12'had9;
        src105 <= 12'he00;
        src106 <= 12'h8ac;
        src107 <= 12'h606;
        src108 <= 12'ha2f;
        src109 <= 12'h86e;
        src110 <= 12'he47;
        src111 <= 12'h141;
        src112 <= 12'hc1d;
        src113 <= 12'h6b2;
        src114 <= 12'hf81;
        src115 <= 12'h384;
        src116 <= 12'hbc1;
        src117 <= 12'h850;
        src118 <= 12'h333;
        src119 <= 12'hc36;
        src120 <= 12'ha1a;
        src121 <= 12'h6de;
        src122 <= 12'h5fd;
        src123 <= 12'h568;
        src124 <= 12'he2a;
        src125 <= 12'hddf;
        src126 <= 12'hf9f;
        src127 <= 12'h52;
        src128 <= 12'h713;
        src129 <= 12'h2a7;
        src130 <= 12'hc35;
        src131 <= 12'h2be;
        src132 <= 12'h507;
        src133 <= 12'h524;
        src134 <= 12'h635;
        src135 <= 12'h8d6;
        src136 <= 12'hcca;
        src137 <= 12'h846;
        src138 <= 12'h1f1;
        src139 <= 12'h679;
        src140 <= 12'h596;
        src141 <= 12'ha07;
        src142 <= 12'h3a;
        src143 <= 12'h68e;
        src144 <= 12'ha60;
        src145 <= 12'h73b;
        src146 <= 12'h7d1;
        src147 <= 12'hb02;
        src148 <= 12'h1c;
        src149 <= 12'h4c5;
        src150 <= 12'h17b;
        src151 <= 12'h28a;
        src152 <= 12'hf22;
        src153 <= 12'h104;
        src154 <= 12'h2cf;
        src155 <= 12'h6f5;
        src156 <= 12'h713;
        src157 <= 12'hd40;
        src158 <= 12'hd98;
        src159 <= 12'h69d;
        src160 <= 12'h30d;
        src161 <= 12'h18a;
        exp <= 20'h55105;
        #1
        src0 <= 12'hdb2;
        src1 <= 12'hbd9;
        src2 <= 12'h7f8;
        src3 <= 12'h388;
        src4 <= 12'hb32;
        src5 <= 12'hc3e;
        src6 <= 12'h126;
        src7 <= 12'h679;
        src8 <= 12'h3ff;
        src9 <= 12'h265;
        src10 <= 12'hd46;
        src11 <= 12'h59f;
        src12 <= 12'h31d;
        src13 <= 12'hefa;
        src14 <= 12'h151;
        src15 <= 12'he18;
        src16 <= 12'hbdd;
        src17 <= 12'h552;
        src18 <= 12'h2e5;
        src19 <= 12'h5dc;
        src20 <= 12'hd10;
        src21 <= 12'hd93;
        src22 <= 12'haf6;
        src23 <= 12'hbf;
        src24 <= 12'h5b6;
        src25 <= 12'h82c;
        src26 <= 12'h353;
        src27 <= 12'ha40;
        src28 <= 12'h743;
        src29 <= 12'hec6;
        src30 <= 12'h3d3;
        src31 <= 12'h4cc;
        src32 <= 12'h69b;
        src33 <= 12'h9a0;
        src34 <= 12'h802;
        src35 <= 12'h692;
        src36 <= 12'he44;
        src37 <= 12'hb8a;
        src38 <= 12'h5a9;
        src39 <= 12'hb22;
        src40 <= 12'hafd;
        src41 <= 12'hae0;
        src42 <= 12'h659;
        src43 <= 12'ha06;
        src44 <= 12'ha41;
        src45 <= 12'h22f;
        src46 <= 12'h2a4;
        src47 <= 12'hd0a;
        src48 <= 12'hf83;
        src49 <= 12'h530;
        src50 <= 12'hb79;
        src51 <= 12'h424;
        src52 <= 12'h4d1;
        src53 <= 12'hc18;
        src54 <= 12'h883;
        src55 <= 12'hbf1;
        src56 <= 12'h7f3;
        src57 <= 12'h789;
        src58 <= 12'h50b;
        src59 <= 12'hb24;
        src60 <= 12'h98c;
        src61 <= 12'h427;
        src62 <= 12'h872;
        src63 <= 12'hf3a;
        src64 <= 12'h7f6;
        src65 <= 12'h45a;
        src66 <= 12'h170;
        src67 <= 12'hd49;
        src68 <= 12'h3ee;
        src69 <= 12'h6c5;
        src70 <= 12'h136;
        src71 <= 12'hb49;
        src72 <= 12'ha7c;
        src73 <= 12'hc3a;
        src74 <= 12'h65f;
        src75 <= 12'hfa0;
        src76 <= 12'h389;
        src77 <= 12'h5a4;
        src78 <= 12'he8a;
        src79 <= 12'h77a;
        src80 <= 12'h6a0;
        src81 <= 12'h9e9;
        src82 <= 12'hfdd;
        src83 <= 12'h931;
        src84 <= 12'hf91;
        src85 <= 12'h92c;
        src86 <= 12'hc37;
        src87 <= 12'he33;
        src88 <= 12'h1f3;
        src89 <= 12'hcb8;
        src90 <= 12'h41c;
        src91 <= 12'h53d;
        src92 <= 12'h323;
        src93 <= 12'h561;
        src94 <= 12'hf25;
        src95 <= 12'h39e;
        src96 <= 12'h543;
        src97 <= 12'hae;
        src98 <= 12'hcfe;
        src99 <= 12'h36;
        src100 <= 12'hd5a;
        src101 <= 12'h658;
        src102 <= 12'hd76;
        src103 <= 12'h695;
        src104 <= 12'h683;
        src105 <= 12'h2c8;
        src106 <= 12'h922;
        src107 <= 12'hca8;
        src108 <= 12'h8a5;
        src109 <= 12'h14e;
        src110 <= 12'hb7e;
        src111 <= 12'h974;
        src112 <= 12'h6e6;
        src113 <= 12'h2a;
        src114 <= 12'h53b;
        src115 <= 12'h6ff;
        src116 <= 12'h414;
        src117 <= 12'h69f;
        src118 <= 12'h7f8;
        src119 <= 12'hb7b;
        src120 <= 12'ha1c;
        src121 <= 12'h837;
        src122 <= 12'h3e5;
        src123 <= 12'h9cc;
        src124 <= 12'hf78;
        src125 <= 12'h1eb;
        src126 <= 12'h146;
        src127 <= 12'h799;
        src128 <= 12'h39d;
        src129 <= 12'h1a3;
        src130 <= 12'h281;
        src131 <= 12'h252;
        src132 <= 12'haba;
        src133 <= 12'hb54;
        src134 <= 12'hb02;
        src135 <= 12'h88;
        src136 <= 12'h5ed;
        src137 <= 12'h152;
        src138 <= 12'h345;
        src139 <= 12'h3eb;
        src140 <= 12'h69a;
        src141 <= 12'h906;
        src142 <= 12'h35;
        src143 <= 12'he9b;
        src144 <= 12'h8dc;
        src145 <= 12'h5d9;
        src146 <= 12'hebf;
        src147 <= 12'ha2c;
        src148 <= 12'ha4;
        src149 <= 12'hca6;
        src150 <= 12'ha68;
        src151 <= 12'h771;
        src152 <= 12'h6ac;
        src153 <= 12'hb9;
        src154 <= 12'hb78;
        src155 <= 12'hd49;
        src156 <= 12'hd1e;
        src157 <= 12'hfb2;
        src158 <= 12'h62a;
        src159 <= 12'h87e;
        src160 <= 12'h33;
        src161 <= 12'h12e;
        exp <= 20'h4f2c9;
        #1
        src0 <= 12'ha0a;
        src1 <= 12'h7e6;
        src2 <= 12'h7d1;
        src3 <= 12'h427;
        src4 <= 12'hd0e;
        src5 <= 12'hb1a;
        src6 <= 12'h5ca;
        src7 <= 12'h2a6;
        src8 <= 12'he18;
        src9 <= 12'hba6;
        src10 <= 12'h6a6;
        src11 <= 12'h555;
        src12 <= 12'hf77;
        src13 <= 12'h9c3;
        src14 <= 12'h3b1;
        src15 <= 12'hc34;
        src16 <= 12'hec9;
        src17 <= 12'h923;
        src18 <= 12'h652;
        src19 <= 12'h8f4;
        src20 <= 12'hcd3;
        src21 <= 12'he9a;
        src22 <= 12'h808;
        src23 <= 12'h5b5;
        src24 <= 12'hd29;
        src25 <= 12'hf4b;
        src26 <= 12'h708;
        src27 <= 12'h565;
        src28 <= 12'h270;
        src29 <= 12'h318;
        src30 <= 12'h301;
        src31 <= 12'h47c;
        src32 <= 12'hb60;
        src33 <= 12'h1cf;
        src34 <= 12'hc10;
        src35 <= 12'hcf5;
        src36 <= 12'h21c;
        src37 <= 12'h51c;
        src38 <= 12'h910;
        src39 <= 12'he1f;
        src40 <= 12'h14;
        src41 <= 12'h5ad;
        src42 <= 12'h2a6;
        src43 <= 12'h259;
        src44 <= 12'he;
        src45 <= 12'h83;
        src46 <= 12'hd32;
        src47 <= 12'h670;
        src48 <= 12'h757;
        src49 <= 12'h2fe;
        src50 <= 12'hc0d;
        src51 <= 12'hbe1;
        src52 <= 12'h3bf;
        src53 <= 12'hd43;
        src54 <= 12'ha5;
        src55 <= 12'h43f;
        src56 <= 12'hec8;
        src57 <= 12'h5bb;
        src58 <= 12'h8c;
        src59 <= 12'h246;
        src60 <= 12'h838;
        src61 <= 12'hfc0;
        src62 <= 12'hf22;
        src63 <= 12'hc35;
        src64 <= 12'hd2e;
        src65 <= 12'h7be;
        src66 <= 12'h991;
        src67 <= 12'h4a5;
        src68 <= 12'he2b;
        src69 <= 12'h69a;
        src70 <= 12'ha3;
        src71 <= 12'hfbb;
        src72 <= 12'hdf9;
        src73 <= 12'h258;
        src74 <= 12'hf2e;
        src75 <= 12'h1a1;
        src76 <= 12'h4dc;
        src77 <= 12'ha9d;
        src78 <= 12'h346;
        src79 <= 12'h627;
        src80 <= 12'h4ba;
        src81 <= 12'hd86;
        src82 <= 12'hcfc;
        src83 <= 12'h853;
        src84 <= 12'ha10;
        src85 <= 12'h793;
        src86 <= 12'hf73;
        src87 <= 12'h17e;
        src88 <= 12'ha6e;
        src89 <= 12'hacb;
        src90 <= 12'h45e;
        src91 <= 12'h277;
        src92 <= 12'hade;
        src93 <= 12'hae3;
        src94 <= 12'hf87;
        src95 <= 12'h8c9;
        src96 <= 12'hb51;
        src97 <= 12'hecc;
        src98 <= 12'h34;
        src99 <= 12'hddc;
        src100 <= 12'h45c;
        src101 <= 12'h394;
        src102 <= 12'h765;
        src103 <= 12'hd33;
        src104 <= 12'hb13;
        src105 <= 12'h55b;
        src106 <= 12'hf45;
        src107 <= 12'hf4f;
        src108 <= 12'h8c2;
        src109 <= 12'hf0b;
        src110 <= 12'h914;
        src111 <= 12'h8e7;
        src112 <= 12'h260;
        src113 <= 12'h56c;
        src114 <= 12'h6e1;
        src115 <= 12'h4f;
        src116 <= 12'h5a3;
        src117 <= 12'ha45;
        src118 <= 12'hf26;
        src119 <= 12'h21d;
        src120 <= 12'hdb5;
        src121 <= 12'h2e;
        src122 <= 12'h3df;
        src123 <= 12'h39b;
        src124 <= 12'ha75;
        src125 <= 12'h7ed;
        src126 <= 12'h93;
        src127 <= 12'h8d5;
        src128 <= 12'hb1f;
        src129 <= 12'h918;
        src130 <= 12'hce4;
        src131 <= 12'h775;
        src132 <= 12'h4dd;
        src133 <= 12'h22f;
        src134 <= 12'he7;
        src135 <= 12'h4bb;
        src136 <= 12'h62c;
        src137 <= 12'hbaa;
        src138 <= 12'h75f;
        src139 <= 12'h3d6;
        src140 <= 12'h23a;
        src141 <= 12'h6ab;
        src142 <= 12'hc14;
        src143 <= 12'ha43;
        src144 <= 12'h7bf;
        src145 <= 12'hd61;
        src146 <= 12'h999;
        src147 <= 12'h3b7;
        src148 <= 12'hab5;
        src149 <= 12'heb0;
        src150 <= 12'h17e;
        src151 <= 12'h555;
        src152 <= 12'had9;
        src153 <= 12'h108;
        src154 <= 12'hfa2;
        src155 <= 12'hdb0;
        src156 <= 12'hee;
        src157 <= 12'h133;
        src158 <= 12'h73b;
        src159 <= 12'h7d2;
        src160 <= 12'hda;
        src161 <= 12'hdf0;
        exp <= 20'h50ca7;
        #1
        src0 <= 12'h64b;
        src1 <= 12'h169;
        src2 <= 12'hf3d;
        src3 <= 12'h7bd;
        src4 <= 12'ha26;
        src5 <= 12'hd7a;
        src6 <= 12'h564;
        src7 <= 12'h1df;
        src8 <= 12'hb61;
        src9 <= 12'hb08;
        src10 <= 12'he24;
        src11 <= 12'hc1e;
        src12 <= 12'ha59;
        src13 <= 12'h16f;
        src14 <= 12'hd20;
        src15 <= 12'h540;
        src16 <= 12'h49e;
        src17 <= 12'h71a;
        src18 <= 12'h98e;
        src19 <= 12'hc43;
        src20 <= 12'hfe2;
        src21 <= 12'he58;
        src22 <= 12'h871;
        src23 <= 12'h8d1;
        src24 <= 12'hd46;
        src25 <= 12'he38;
        src26 <= 12'hb88;
        src27 <= 12'hba;
        src28 <= 12'h447;
        src29 <= 12'h898;
        src30 <= 12'hf87;
        src31 <= 12'h467;
        src32 <= 12'hf96;
        src33 <= 12'h79b;
        src34 <= 12'h9a;
        src35 <= 12'hef2;
        src36 <= 12'h48e;
        src37 <= 12'h222;
        src38 <= 12'h52b;
        src39 <= 12'h795;
        src40 <= 12'hc2e;
        src41 <= 12'h5b2;
        src42 <= 12'h100;
        src43 <= 12'h756;
        src44 <= 12'h120;
        src45 <= 12'hbf0;
        src46 <= 12'hb54;
        src47 <= 12'h9b0;
        src48 <= 12'h102;
        src49 <= 12'hc76;
        src50 <= 12'h42a;
        src51 <= 12'hef3;
        src52 <= 12'h365;
        src53 <= 12'h7a5;
        src54 <= 12'h84b;
        src55 <= 12'h84;
        src56 <= 12'h325;
        src57 <= 12'h1cf;
        src58 <= 12'h69c;
        src59 <= 12'h151;
        src60 <= 12'h93c;
        src61 <= 12'ha56;
        src62 <= 12'ha2e;
        src63 <= 12'h400;
        src64 <= 12'h739;
        src65 <= 12'had9;
        src66 <= 12'hcc7;
        src67 <= 12'hd79;
        src68 <= 12'h3dd;
        src69 <= 12'ha5a;
        src70 <= 12'ha96;
        src71 <= 12'h2f2;
        src72 <= 12'h7df;
        src73 <= 12'hf53;
        src74 <= 12'hf6b;
        src75 <= 12'h162;
        src76 <= 12'hcf1;
        src77 <= 12'hd66;
        src78 <= 12'hb4f;
        src79 <= 12'h452;
        src80 <= 12'h257;
        src81 <= 12'h2d5;
        src82 <= 12'hb9d;
        src83 <= 12'h7e8;
        src84 <= 12'h2c7;
        src85 <= 12'hb66;
        src86 <= 12'h184;
        src87 <= 12'h9a5;
        src88 <= 12'he83;
        src89 <= 12'h29d;
        src90 <= 12'hd0c;
        src91 <= 12'h7ec;
        src92 <= 12'ha55;
        src93 <= 12'hc8b;
        src94 <= 12'h74f;
        src95 <= 12'h9dd;
        src96 <= 12'hb72;
        src97 <= 12'h1ab;
        src98 <= 12'h4e5;
        src99 <= 12'h258;
        src100 <= 12'h990;
        src101 <= 12'h269;
        src102 <= 12'h4fa;
        src103 <= 12'h1d1;
        src104 <= 12'h669;
        src105 <= 12'h2d9;
        src106 <= 12'hc1b;
        src107 <= 12'h585;
        src108 <= 12'h80;
        src109 <= 12'h695;
        src110 <= 12'h94;
        src111 <= 12'h547;
        src112 <= 12'h7f7;
        src113 <= 12'h889;
        src114 <= 12'haef;
        src115 <= 12'hc6c;
        src116 <= 12'hcbf;
        src117 <= 12'hf71;
        src118 <= 12'h5e7;
        src119 <= 12'hfd5;
        src120 <= 12'hb30;
        src121 <= 12'hf98;
        src122 <= 12'h9ba;
        src123 <= 12'hd0;
        src124 <= 12'hc27;
        src125 <= 12'h984;
        src126 <= 12'hdb3;
        src127 <= 12'hf3b;
        src128 <= 12'hf41;
        src129 <= 12'h3c5;
        src130 <= 12'h262;
        src131 <= 12'hc7f;
        src132 <= 12'hff5;
        src133 <= 12'h945;
        src134 <= 12'h70a;
        src135 <= 12'h6b8;
        src136 <= 12'h240;
        src137 <= 12'h906;
        src138 <= 12'haa7;
        src139 <= 12'hed1;
        src140 <= 12'h351;
        src141 <= 12'h31a;
        src142 <= 12'h82e;
        src143 <= 12'hf96;
        src144 <= 12'h99a;
        src145 <= 12'h9d3;
        src146 <= 12'h7eb;
        src147 <= 12'hdb4;
        src148 <= 12'ha8;
        src149 <= 12'hb35;
        src150 <= 12'hd63;
        src151 <= 12'h27b;
        src152 <= 12'h604;
        src153 <= 12'h182;
        src154 <= 12'h7ba;
        src155 <= 12'h73d;
        src156 <= 12'hcb1;
        src157 <= 12'hd82;
        src158 <= 12'h8;
        src159 <= 12'hba5;
        src160 <= 12'he7;
        src161 <= 12'h6c7;
        exp <= 20'h52ef3;
        #1
        src0 <= 12'hd80;
        src1 <= 12'hf22;
        src2 <= 12'h6b9;
        src3 <= 12'h9f6;
        src4 <= 12'h335;
        src5 <= 12'hdf7;
        src6 <= 12'h2e7;
        src7 <= 12'h742;
        src8 <= 12'h3be;
        src9 <= 12'hbb8;
        src10 <= 12'h2b7;
        src11 <= 12'hde4;
        src12 <= 12'h7e5;
        src13 <= 12'hf48;
        src14 <= 12'hcb9;
        src15 <= 12'hb15;
        src16 <= 12'hbc8;
        src17 <= 12'hf82;
        src18 <= 12'hf32;
        src19 <= 12'h6f9;
        src20 <= 12'h3eb;
        src21 <= 12'hb3b;
        src22 <= 12'h119;
        src23 <= 12'h86d;
        src24 <= 12'h28c;
        src25 <= 12'hd0;
        src26 <= 12'h405;
        src27 <= 12'hf5a;
        src28 <= 12'hf37;
        src29 <= 12'h641;
        src30 <= 12'ha51;
        src31 <= 12'h5fe;
        src32 <= 12'h839;
        src33 <= 12'h7b6;
        src34 <= 12'hbee;
        src35 <= 12'h7a8;
        src36 <= 12'hf52;
        src37 <= 12'hda4;
        src38 <= 12'ha91;
        src39 <= 12'hc5a;
        src40 <= 12'he27;
        src41 <= 12'hbae;
        src42 <= 12'h97a;
        src43 <= 12'h4f3;
        src44 <= 12'hd48;
        src45 <= 12'h63b;
        src46 <= 12'h280;
        src47 <= 12'h558;
        src48 <= 12'h96e;
        src49 <= 12'ha9;
        src50 <= 12'heab;
        src51 <= 12'h524;
        src52 <= 12'haea;
        src53 <= 12'h27;
        src54 <= 12'h77b;
        src55 <= 12'h88d;
        src56 <= 12'h9b6;
        src57 <= 12'h6da;
        src58 <= 12'h266;
        src59 <= 12'h723;
        src60 <= 12'h3d0;
        src61 <= 12'ha15;
        src62 <= 12'h616;
        src63 <= 12'hcab;
        src64 <= 12'haa7;
        src65 <= 12'hdf9;
        src66 <= 12'h9ca;
        src67 <= 12'h71c;
        src68 <= 12'h1fe;
        src69 <= 12'h99e;
        src70 <= 12'h15b;
        src71 <= 12'h6ac;
        src72 <= 12'hd26;
        src73 <= 12'h455;
        src74 <= 12'hc9e;
        src75 <= 12'hf64;
        src76 <= 12'h43a;
        src77 <= 12'h349;
        src78 <= 12'h852;
        src79 <= 12'hefc;
        src80 <= 12'h45c;
        src81 <= 12'ha70;
        src82 <= 12'h668;
        src83 <= 12'hd0c;
        src84 <= 12'h1cb;
        src85 <= 12'h902;
        src86 <= 12'h999;
        src87 <= 12'h1a2;
        src88 <= 12'h3f9;
        src89 <= 12'h50d;
        src90 <= 12'h848;
        src91 <= 12'hdb;
        src92 <= 12'h9e0;
        src93 <= 12'h86c;
        src94 <= 12'hfc4;
        src95 <= 12'h370;
        src96 <= 12'h192;
        src97 <= 12'h509;
        src98 <= 12'hbf5;
        src99 <= 12'h265;
        src100 <= 12'h8dc;
        src101 <= 12'h127;
        src102 <= 12'h3a1;
        src103 <= 12'hddb;
        src104 <= 12'hdf5;
        src105 <= 12'h438;
        src106 <= 12'h81e;
        src107 <= 12'h9ee;
        src108 <= 12'hc83;
        src109 <= 12'hb3e;
        src110 <= 12'h5d8;
        src111 <= 12'h444;
        src112 <= 12'haec;
        src113 <= 12'hbc5;
        src114 <= 12'hb06;
        src115 <= 12'h144;
        src116 <= 12'h9e2;
        src117 <= 12'hf39;
        src118 <= 12'h110;
        src119 <= 12'h67d;
        src120 <= 12'h584;
        src121 <= 12'h760;
        src122 <= 12'hede;
        src123 <= 12'h8ae;
        src124 <= 12'he2;
        src125 <= 12'hf8;
        src126 <= 12'h733;
        src127 <= 12'ha6f;
        src128 <= 12'h2b4;
        src129 <= 12'ha91;
        src130 <= 12'h848;
        src131 <= 12'h585;
        src132 <= 12'h8f5;
        src133 <= 12'hf8e;
        src134 <= 12'hef6;
        src135 <= 12'hf91;
        src136 <= 12'he84;
        src137 <= 12'h7a7;
        src138 <= 12'hd58;
        src139 <= 12'h961;
        src140 <= 12'hef3;
        src141 <= 12'h5d3;
        src142 <= 12'h64c;
        src143 <= 12'hd4;
        src144 <= 12'h72f;
        src145 <= 12'h72b;
        src146 <= 12'h476;
        src147 <= 12'ha82;
        src148 <= 12'h8a2;
        src149 <= 12'hca8;
        src150 <= 12'h533;
        src151 <= 12'hcac;
        src152 <= 12'h6cc;
        src153 <= 12'h14c;
        src154 <= 12'h243;
        src155 <= 12'h979;
        src156 <= 12'h9f0;
        src157 <= 12'hb73;
        src158 <= 12'h21e;
        src159 <= 12'h7c6;
        src160 <= 12'h7b8;
        src161 <= 12'ha40;
        exp <= 20'h53d0b;
        #1
        src0 <= 12'h3c7;
        src1 <= 12'hc58;
        src2 <= 12'hba7;
        src3 <= 12'h39d;
        src4 <= 12'h367;
        src5 <= 12'h3ab;
        src6 <= 12'h565;
        src7 <= 12'hae6;
        src8 <= 12'h859;
        src9 <= 12'h824;
        src10 <= 12'h17f;
        src11 <= 12'hd99;
        src12 <= 12'hb7c;
        src13 <= 12'h46c;
        src14 <= 12'hb3b;
        src15 <= 12'h188;
        src16 <= 12'h311;
        src17 <= 12'hc77;
        src18 <= 12'hd49;
        src19 <= 12'hc1a;
        src20 <= 12'h4a;
        src21 <= 12'h23b;
        src22 <= 12'h1bd;
        src23 <= 12'h492;
        src24 <= 12'h5f9;
        src25 <= 12'hd6f;
        src26 <= 12'h53f;
        src27 <= 12'he54;
        src28 <= 12'h4cb;
        src29 <= 12'h188;
        src30 <= 12'hb43;
        src31 <= 12'h4b5;
        src32 <= 12'h13e;
        src33 <= 12'h9c4;
        src34 <= 12'hb9f;
        src35 <= 12'ha61;
        src36 <= 12'h7b2;
        src37 <= 12'he;
        src38 <= 12'h3d6;
        src39 <= 12'h5d4;
        src40 <= 12'h5ab;
        src41 <= 12'h341;
        src42 <= 12'hb9e;
        src43 <= 12'h4d2;
        src44 <= 12'h9c8;
        src45 <= 12'h529;
        src46 <= 12'h191;
        src47 <= 12'h209;
        src48 <= 12'h54d;
        src49 <= 12'hf3a;
        src50 <= 12'hf43;
        src51 <= 12'hb62;
        src52 <= 12'hbb2;
        src53 <= 12'hd7d;
        src54 <= 12'h71a;
        src55 <= 12'hcfb;
        src56 <= 12'he5;
        src57 <= 12'ha8e;
        src58 <= 12'ha23;
        src59 <= 12'h543;
        src60 <= 12'hc87;
        src61 <= 12'h8dd;
        src62 <= 12'hc50;
        src63 <= 12'ha2a;
        src64 <= 12'hc73;
        src65 <= 12'hdae;
        src66 <= 12'h37f;
        src67 <= 12'h141;
        src68 <= 12'h3e1;
        src69 <= 12'h6f4;
        src70 <= 12'h68f;
        src71 <= 12'h7c5;
        src72 <= 12'he35;
        src73 <= 12'h5cb;
        src74 <= 12'h7c4;
        src75 <= 12'ha3f;
        src76 <= 12'ha9c;
        src77 <= 12'h7af;
        src78 <= 12'hc45;
        src79 <= 12'h951;
        src80 <= 12'h348;
        src81 <= 12'hffe;
        src82 <= 12'hdb;
        src83 <= 12'h7b1;
        src84 <= 12'h209;
        src85 <= 12'ha6d;
        src86 <= 12'h6fc;
        src87 <= 12'h58a;
        src88 <= 12'h428;
        src89 <= 12'h9f0;
        src90 <= 12'h670;
        src91 <= 12'h16f;
        src92 <= 12'h2c4;
        src93 <= 12'h97f;
        src94 <= 12'hbf0;
        src95 <= 12'h60e;
        src96 <= 12'he88;
        src97 <= 12'hf28;
        src98 <= 12'ha00;
        src99 <= 12'h128;
        src100 <= 12'h5d1;
        src101 <= 12'h36f;
        src102 <= 12'h7bc;
        src103 <= 12'hde7;
        src104 <= 12'he1b;
        src105 <= 12'he48;
        src106 <= 12'h288;
        src107 <= 12'haad;
        src108 <= 12'h281;
        src109 <= 12'h620;
        src110 <= 12'hadd;
        src111 <= 12'hfd;
        src112 <= 12'h111;
        src113 <= 12'h3bf;
        src114 <= 12'hc6f;
        src115 <= 12'h537;
        src116 <= 12'h3b8;
        src117 <= 12'hb89;
        src118 <= 12'ha60;
        src119 <= 12'h369;
        src120 <= 12'h49c;
        src121 <= 12'h172;
        src122 <= 12'h311;
        src123 <= 12'h185;
        src124 <= 12'h1bd;
        src125 <= 12'hb80;
        src126 <= 12'hcdd;
        src127 <= 12'h3cd;
        src128 <= 12'h39a;
        src129 <= 12'hfd7;
        src130 <= 12'h617;
        src131 <= 12'h4f0;
        src132 <= 12'hc51;
        src133 <= 12'ha5;
        src134 <= 12'h444;
        src135 <= 12'h371;
        src136 <= 12'h12c;
        src137 <= 12'hb56;
        src138 <= 12'h38a;
        src139 <= 12'h4b4;
        src140 <= 12'h861;
        src141 <= 12'h4ca;
        src142 <= 12'h665;
        src143 <= 12'hb58;
        src144 <= 12'hf50;
        src145 <= 12'hefc;
        src146 <= 12'he76;
        src147 <= 12'ha3d;
        src148 <= 12'h553;
        src149 <= 12'hcbf;
        src150 <= 12'h780;
        src151 <= 12'hb24;
        src152 <= 12'h417;
        src153 <= 12'he9e;
        src154 <= 12'hade;
        src155 <= 12'h9ff;
        src156 <= 12'ha91;
        src157 <= 12'hd4;
        src158 <= 12'hdaf;
        src159 <= 12'h775;
        src160 <= 12'h8a0;
        src161 <= 12'h96a;
        exp <= 20'h4d0f1;
        #1
        src0 <= 12'h50f;
        src1 <= 12'h384;
        src2 <= 12'hf81;
        src3 <= 12'h2c2;
        src4 <= 12'h6c2;
        src5 <= 12'h581;
        src6 <= 12'hdc4;
        src7 <= 12'h465;
        src8 <= 12'hedd;
        src9 <= 12'h880;
        src10 <= 12'h61;
        src11 <= 12'hea6;
        src12 <= 12'h1e6;
        src13 <= 12'hb34;
        src14 <= 12'h955;
        src15 <= 12'h2b3;
        src16 <= 12'h1bf;
        src17 <= 12'h2d4;
        src18 <= 12'h48b;
        src19 <= 12'h7f0;
        src20 <= 12'he2b;
        src21 <= 12'h331;
        src22 <= 12'hb82;
        src23 <= 12'hb26;
        src24 <= 12'h39f;
        src25 <= 12'h7d4;
        src26 <= 12'h802;
        src27 <= 12'h703;
        src28 <= 12'hf8b;
        src29 <= 12'h385;
        src30 <= 12'h6c;
        src31 <= 12'hd06;
        src32 <= 12'h134;
        src33 <= 12'h270;
        src34 <= 12'h3f5;
        src35 <= 12'hebf;
        src36 <= 12'h56c;
        src37 <= 12'h81a;
        src38 <= 12'hed5;
        src39 <= 12'he16;
        src40 <= 12'h22;
        src41 <= 12'h3d4;
        src42 <= 12'h4da;
        src43 <= 12'h3a7;
        src44 <= 12'h3a3;
        src45 <= 12'h726;
        src46 <= 12'heb0;
        src47 <= 12'h33f;
        src48 <= 12'hd4e;
        src49 <= 12'ha6c;
        src50 <= 12'h484;
        src51 <= 12'h1b;
        src52 <= 12'h6e;
        src53 <= 12'hb21;
        src54 <= 12'hae1;
        src55 <= 12'h56b;
        src56 <= 12'h382;
        src57 <= 12'h539;
        src58 <= 12'h6dc;
        src59 <= 12'h2fc;
        src60 <= 12'h4c4;
        src61 <= 12'h887;
        src62 <= 12'hcc7;
        src63 <= 12'h621;
        src64 <= 12'h686;
        src65 <= 12'h5ac;
        src66 <= 12'h9f9;
        src67 <= 12'h458;
        src68 <= 12'h26c;
        src69 <= 12'h8a;
        src70 <= 12'h909;
        src71 <= 12'h12f;
        src72 <= 12'hb1c;
        src73 <= 12'h138;
        src74 <= 12'h518;
        src75 <= 12'h70;
        src76 <= 12'h825;
        src77 <= 12'h525;
        src78 <= 12'hb9b;
        src79 <= 12'h736;
        src80 <= 12'h693;
        src81 <= 12'h249;
        src82 <= 12'had0;
        src83 <= 12'hd8d;
        src84 <= 12'hbc0;
        src85 <= 12'h90b;
        src86 <= 12'he6b;
        src87 <= 12'hca9;
        src88 <= 12'h9f0;
        src89 <= 12'h6ed;
        src90 <= 12'hf4a;
        src91 <= 12'h4e4;
        src92 <= 12'h78;
        src93 <= 12'h1f9;
        src94 <= 12'h9b3;
        src95 <= 12'h8d4;
        src96 <= 12'h793;
        src97 <= 12'h8b8;
        src98 <= 12'hb84;
        src99 <= 12'h7f8;
        src100 <= 12'h7c6;
        src101 <= 12'hc4c;
        src102 <= 12'hd64;
        src103 <= 12'h42;
        src104 <= 12'h740;
        src105 <= 12'ha3b;
        src106 <= 12'h861;
        src107 <= 12'h61c;
        src108 <= 12'h91e;
        src109 <= 12'h9fc;
        src110 <= 12'hccd;
        src111 <= 12'h790;
        src112 <= 12'hd9d;
        src113 <= 12'h888;
        src114 <= 12'hadc;
        src115 <= 12'h242;
        src116 <= 12'h6d;
        src117 <= 12'h7b3;
        src118 <= 12'he3f;
        src119 <= 12'h325;
        src120 <= 12'h6ee;
        src121 <= 12'hce4;
        src122 <= 12'h7d3;
        src123 <= 12'h1b1;
        src124 <= 12'h7a8;
        src125 <= 12'hdde;
        src126 <= 12'hbb9;
        src127 <= 12'h296;
        src128 <= 12'h4f;
        src129 <= 12'h27c;
        src130 <= 12'h94;
        src131 <= 12'h2cf;
        src132 <= 12'hc0d;
        src133 <= 12'h1ee;
        src134 <= 12'h325;
        src135 <= 12'h938;
        src136 <= 12'h1e4;
        src137 <= 12'h461;
        src138 <= 12'h1f6;
        src139 <= 12'h9fb;
        src140 <= 12'hfb3;
        src141 <= 12'h6c9;
        src142 <= 12'hd07;
        src143 <= 12'h8cf;
        src144 <= 12'hb4d;
        src145 <= 12'h90;
        src146 <= 12'h25a;
        src147 <= 12'h625;
        src148 <= 12'hc4f;
        src149 <= 12'hedf;
        src150 <= 12'he8e;
        src151 <= 12'h1d1;
        src152 <= 12'he48;
        src153 <= 12'h450;
        src154 <= 12'ha0a;
        src155 <= 12'hcbb;
        src156 <= 12'he03;
        src157 <= 12'h831;
        src158 <= 12'h1b1;
        src159 <= 12'hc04;
        src160 <= 12'hded;
        src161 <= 12'hfb3;
        exp <= 20'h4bb46;
        #1
        src0 <= 12'h7d5;
        src1 <= 12'hbb0;
        src2 <= 12'h3f7;
        src3 <= 12'h63b;
        src4 <= 12'h41d;
        src5 <= 12'h9d5;
        src6 <= 12'hf4f;
        src7 <= 12'h16f;
        src8 <= 12'h775;
        src9 <= 12'h961;
        src10 <= 12'h45a;
        src11 <= 12'h529;
        src12 <= 12'had2;
        src13 <= 12'hf79;
        src14 <= 12'h2dc;
        src15 <= 12'hf5f;
        src16 <= 12'h6d6;
        src17 <= 12'h8df;
        src18 <= 12'hba1;
        src19 <= 12'h8f6;
        src20 <= 12'hc42;
        src21 <= 12'h31e;
        src22 <= 12'h44a;
        src23 <= 12'h719;
        src24 <= 12'ha0c;
        src25 <= 12'h63a;
        src26 <= 12'h352;
        src27 <= 12'ha93;
        src28 <= 12'hc3a;
        src29 <= 12'h54;
        src30 <= 12'h9bb;
        src31 <= 12'h2b8;
        src32 <= 12'hef7;
        src33 <= 12'h968;
        src34 <= 12'h562;
        src35 <= 12'h86a;
        src36 <= 12'h41b;
        src37 <= 12'h9d9;
        src38 <= 12'h465;
        src39 <= 12'ha3f;
        src40 <= 12'h785;
        src41 <= 12'h146;
        src42 <= 12'h2e3;
        src43 <= 12'hf8f;
        src44 <= 12'h1f1;
        src45 <= 12'h7d7;
        src46 <= 12'h9e3;
        src47 <= 12'ha04;
        src48 <= 12'h7a7;
        src49 <= 12'h8b8;
        src50 <= 12'hddb;
        src51 <= 12'h2a;
        src52 <= 12'h9b1;
        src53 <= 12'hb24;
        src54 <= 12'h451;
        src55 <= 12'h1a;
        src56 <= 12'h2d4;
        src57 <= 12'hb7f;
        src58 <= 12'h1c9;
        src59 <= 12'h57e;
        src60 <= 12'h139;
        src61 <= 12'hb71;
        src62 <= 12'h171;
        src63 <= 12'h1ff;
        src64 <= 12'hc00;
        src65 <= 12'h84b;
        src66 <= 12'h309;
        src67 <= 12'h181;
        src68 <= 12'h5dd;
        src69 <= 12'hae1;
        src70 <= 12'hae3;
        src71 <= 12'h5bc;
        src72 <= 12'hba4;
        src73 <= 12'hdf1;
        src74 <= 12'h870;
        src75 <= 12'h17d;
        src76 <= 12'hcf9;
        src77 <= 12'h741;
        src78 <= 12'hdf6;
        src79 <= 12'h673;
        src80 <= 12'hee9;
        src81 <= 12'h90c;
        src82 <= 12'hede;
        src83 <= 12'h66c;
        src84 <= 12'hed0;
        src85 <= 12'h302;
        src86 <= 12'h9f4;
        src87 <= 12'h9e6;
        src88 <= 12'h96a;
        src89 <= 12'hd10;
        src90 <= 12'h4;
        src91 <= 12'hbe6;
        src92 <= 12'h5ca;
        src93 <= 12'h385;
        src94 <= 12'h225;
        src95 <= 12'h39a;
        src96 <= 12'he4a;
        src97 <= 12'h291;
        src98 <= 12'h709;
        src99 <= 12'ha34;
        src100 <= 12'ha87;
        src101 <= 12'h2fd;
        src102 <= 12'h61e;
        src103 <= 12'hc01;
        src104 <= 12'h1cf;
        src105 <= 12'hbf6;
        src106 <= 12'h212;
        src107 <= 12'hc23;
        src108 <= 12'h80e;
        src109 <= 12'h5e2;
        src110 <= 12'h794;
        src111 <= 12'h4f7;
        src112 <= 12'h364;
        src113 <= 12'hcf6;
        src114 <= 12'hfb7;
        src115 <= 12'hf71;
        src116 <= 12'hc72;
        src117 <= 12'hfaf;
        src118 <= 12'hfae;
        src119 <= 12'h7ef;
        src120 <= 12'h859;
        src121 <= 12'h2af;
        src122 <= 12'hb53;
        src123 <= 12'haaf;
        src124 <= 12'hfcd;
        src125 <= 12'h1a5;
        src126 <= 12'heb8;
        src127 <= 12'h3e8;
        src128 <= 12'h256;
        src129 <= 12'h689;
        src130 <= 12'haa5;
        src131 <= 12'h9f2;
        src132 <= 12'h551;
        src133 <= 12'hca;
        src134 <= 12'hb2d;
        src135 <= 12'h138;
        src136 <= 12'h8ed;
        src137 <= 12'h2da;
        src138 <= 12'h5b6;
        src139 <= 12'he9;
        src140 <= 12'h3dd;
        src141 <= 12'hc4c;
        src142 <= 12'h402;
        src143 <= 12'ha10;
        src144 <= 12'h8c0;
        src145 <= 12'hee5;
        src146 <= 12'hbda;
        src147 <= 12'hc2c;
        src148 <= 12'hf0c;
        src149 <= 12'hf7e;
        src150 <= 12'hddd;
        src151 <= 12'hfc;
        src152 <= 12'hfe1;
        src153 <= 12'h95f;
        src154 <= 12'hbfc;
        src155 <= 12'he6b;
        src156 <= 12'hde3;
        src157 <= 12'hcdc;
        src158 <= 12'h3de;
        src159 <= 12'h829;
        src160 <= 12'h158;
        src161 <= 12'h15b;
        exp <= 20'h5188d;
        #1
        src0 <= 12'hab1;
        src1 <= 12'hccd;
        src2 <= 12'h35d;
        src3 <= 12'h9c8;
        src4 <= 12'h190;
        src5 <= 12'h1f;
        src6 <= 12'hac0;
        src7 <= 12'h26d;
        src8 <= 12'h821;
        src9 <= 12'h88c;
        src10 <= 12'h496;
        src11 <= 12'hc08;
        src12 <= 12'hf1c;
        src13 <= 12'h328;
        src14 <= 12'h928;
        src15 <= 12'hc4d;
        src16 <= 12'hff3;
        src17 <= 12'h398;
        src18 <= 12'h353;
        src19 <= 12'h814;
        src20 <= 12'h339;
        src21 <= 12'h2f;
        src22 <= 12'h67c;
        src23 <= 12'h536;
        src24 <= 12'h3d7;
        src25 <= 12'hf94;
        src26 <= 12'heb4;
        src27 <= 12'h145;
        src28 <= 12'hf2e;
        src29 <= 12'h23a;
        src30 <= 12'h42d;
        src31 <= 12'h645;
        src32 <= 12'hce0;
        src33 <= 12'hddf;
        src34 <= 12'h2d1;
        src35 <= 12'h92d;
        src36 <= 12'he0c;
        src37 <= 12'hb05;
        src38 <= 12'h766;
        src39 <= 12'h5cb;
        src40 <= 12'h77d;
        src41 <= 12'h11;
        src42 <= 12'h32b;
        src43 <= 12'h4d;
        src44 <= 12'h29d;
        src45 <= 12'h6e4;
        src46 <= 12'h8d5;
        src47 <= 12'haa3;
        src48 <= 12'h148;
        src49 <= 12'hfce;
        src50 <= 12'hda;
        src51 <= 12'hd70;
        src52 <= 12'h443;
        src53 <= 12'h90a;
        src54 <= 12'h615;
        src55 <= 12'hccb;
        src56 <= 12'he88;
        src57 <= 12'h9b6;
        src58 <= 12'h847;
        src59 <= 12'h33c;
        src60 <= 12'h73e;
        src61 <= 12'h8b2;
        src62 <= 12'hb5f;
        src63 <= 12'h3b6;
        src64 <= 12'hc64;
        src65 <= 12'haad;
        src66 <= 12'h1ec;
        src67 <= 12'h906;
        src68 <= 12'h325;
        src69 <= 12'h36a;
        src70 <= 12'hc95;
        src71 <= 12'h6b4;
        src72 <= 12'h3bd;
        src73 <= 12'h66e;
        src74 <= 12'h8e6;
        src75 <= 12'h8ae;
        src76 <= 12'hba4;
        src77 <= 12'he2d;
        src78 <= 12'h96b;
        src79 <= 12'h5f3;
        src80 <= 12'h788;
        src81 <= 12'hc32;
        src82 <= 12'h72d;
        src83 <= 12'h5bf;
        src84 <= 12'hd84;
        src85 <= 12'h32a;
        src86 <= 12'h5fc;
        src87 <= 12'he13;
        src88 <= 12'h785;
        src89 <= 12'h838;
        src90 <= 12'h8c9;
        src91 <= 12'h25e;
        src92 <= 12'hd5d;
        src93 <= 12'hb0f;
        src94 <= 12'h62;
        src95 <= 12'ha83;
        src96 <= 12'h50a;
        src97 <= 12'hb74;
        src98 <= 12'hd4b;
        src99 <= 12'h95a;
        src100 <= 12'h3b3;
        src101 <= 12'h5ad;
        src102 <= 12'hb11;
        src103 <= 12'h9c4;
        src104 <= 12'h7a1;
        src105 <= 12'hfd6;
        src106 <= 12'h6bc;
        src107 <= 12'h54d;
        src108 <= 12'hb38;
        src109 <= 12'h394;
        src110 <= 12'hb60;
        src111 <= 12'h40f;
        src112 <= 12'ha04;
        src113 <= 12'h326;
        src114 <= 12'h858;
        src115 <= 12'h986;
        src116 <= 12'h396;
        src117 <= 12'hfc8;
        src118 <= 12'hc17;
        src119 <= 12'h99c;
        src120 <= 12'hbca;
        src121 <= 12'h697;
        src122 <= 12'h3f7;
        src123 <= 12'h12f;
        src124 <= 12'hc70;
        src125 <= 12'h4fa;
        src126 <= 12'hf2b;
        src127 <= 12'h60a;
        src128 <= 12'hdd6;
        src129 <= 12'h4;
        src130 <= 12'h6c7;
        src131 <= 12'hba1;
        src132 <= 12'haad;
        src133 <= 12'hd6a;
        src134 <= 12'hd9f;
        src135 <= 12'h6e0;
        src136 <= 12'h34f;
        src137 <= 12'h498;
        src138 <= 12'h1fa;
        src139 <= 12'hf1e;
        src140 <= 12'h606;
        src141 <= 12'he82;
        src142 <= 12'h3c2;
        src143 <= 12'h15f;
        src144 <= 12'hd23;
        src145 <= 12'h56e;
        src146 <= 12'h672;
        src147 <= 12'h1d3;
        src148 <= 12'he0b;
        src149 <= 12'h371;
        src150 <= 12'haa1;
        src151 <= 12'h12f;
        src152 <= 12'h5a2;
        src153 <= 12'h361;
        src154 <= 12'h6be;
        src155 <= 12'h34;
        src156 <= 12'h3a0;
        src157 <= 12'hdc0;
        src158 <= 12'hce9;
        src159 <= 12'ha63;
        src160 <= 12'ha28;
        src161 <= 12'h1c8;
        exp <= 20'h4ef04;
        #1
        src0 <= 12'hf;
        src1 <= 12'h117;
        src2 <= 12'h546;
        src3 <= 12'h97b;
        src4 <= 12'h803;
        src5 <= 12'h724;
        src6 <= 12'h5f1;
        src7 <= 12'h446;
        src8 <= 12'h2e;
        src9 <= 12'h1f5;
        src10 <= 12'h3;
        src11 <= 12'hc6d;
        src12 <= 12'hc57;
        src13 <= 12'hf39;
        src14 <= 12'hfde;
        src15 <= 12'h422;
        src16 <= 12'hf31;
        src17 <= 12'h654;
        src18 <= 12'h391;
        src19 <= 12'h30b;
        src20 <= 12'hce5;
        src21 <= 12'h6af;
        src22 <= 12'h64f;
        src23 <= 12'h63f;
        src24 <= 12'h827;
        src25 <= 12'hab0;
        src26 <= 12'h4bb;
        src27 <= 12'h257;
        src28 <= 12'hdff;
        src29 <= 12'hbe1;
        src30 <= 12'h399;
        src31 <= 12'h9b8;
        src32 <= 12'h32a;
        src33 <= 12'hac;
        src34 <= 12'h373;
        src35 <= 12'hfda;
        src36 <= 12'h5f2;
        src37 <= 12'h39f;
        src38 <= 12'h476;
        src39 <= 12'h447;
        src40 <= 12'h71e;
        src41 <= 12'ha9c;
        src42 <= 12'h277;
        src43 <= 12'hed2;
        src44 <= 12'hed3;
        src45 <= 12'he1f;
        src46 <= 12'h15d;
        src47 <= 12'hd1d;
        src48 <= 12'hb2a;
        src49 <= 12'hf1c;
        src50 <= 12'h6fa;
        src51 <= 12'ha09;
        src52 <= 12'h2b5;
        src53 <= 12'h3c9;
        src54 <= 12'h8d2;
        src55 <= 12'h6d8;
        src56 <= 12'h9ad;
        src57 <= 12'h87e;
        src58 <= 12'h6d;
        src59 <= 12'hbcf;
        src60 <= 12'h39f;
        src61 <= 12'h46c;
        src62 <= 12'hf88;
        src63 <= 12'h3f3;
        src64 <= 12'h717;
        src65 <= 12'h941;
        src66 <= 12'hd3c;
        src67 <= 12'hec1;
        src68 <= 12'ha21;
        src69 <= 12'h607;
        src70 <= 12'h372;
        src71 <= 12'h41c;
        src72 <= 12'hf43;
        src73 <= 12'hbae;
        src74 <= 12'hdc1;
        src75 <= 12'h19f;
        src76 <= 12'h263;
        src77 <= 12'h465;
        src78 <= 12'h28c;
        src79 <= 12'h272;
        src80 <= 12'hae1;
        src81 <= 12'hab5;
        src82 <= 12'h1f;
        src83 <= 12'h7ac;
        src84 <= 12'hba5;
        src85 <= 12'hada;
        src86 <= 12'hef7;
        src87 <= 12'h4c8;
        src88 <= 12'h7fe;
        src89 <= 12'h7d6;
        src90 <= 12'h515;
        src91 <= 12'hd9a;
        src92 <= 12'h9c5;
        src93 <= 12'hd71;
        src94 <= 12'hc40;
        src95 <= 12'h886;
        src96 <= 12'h81b;
        src97 <= 12'h5da;
        src98 <= 12'h285;
        src99 <= 12'h6ed;
        src100 <= 12'h7ca;
        src101 <= 12'he91;
        src102 <= 12'h91;
        src103 <= 12'h648;
        src104 <= 12'h2f3;
        src105 <= 12'h231;
        src106 <= 12'h5ac;
        src107 <= 12'h812;
        src108 <= 12'h514;
        src109 <= 12'h695;
        src110 <= 12'h8d2;
        src111 <= 12'h584;
        src112 <= 12'h325;
        src113 <= 12'h3e;
        src114 <= 12'hbe0;
        src115 <= 12'hc97;
        src116 <= 12'h630;
        src117 <= 12'h710;
        src118 <= 12'hbe5;
        src119 <= 12'hddc;
        src120 <= 12'h71;
        src121 <= 12'ha38;
        src122 <= 12'hf8b;
        src123 <= 12'h16b;
        src124 <= 12'hbf8;
        src125 <= 12'hd9;
        src126 <= 12'hb;
        src127 <= 12'hcae;
        src128 <= 12'h86;
        src129 <= 12'hfa1;
        src130 <= 12'h406;
        src131 <= 12'hd7a;
        src132 <= 12'h764;
        src133 <= 12'h442;
        src134 <= 12'h31e;
        src135 <= 12'h17c;
        src136 <= 12'h62a;
        src137 <= 12'hd35;
        src138 <= 12'h92d;
        src139 <= 12'h41;
        src140 <= 12'h6f1;
        src141 <= 12'h16b;
        src142 <= 12'haa2;
        src143 <= 12'hbfb;
        src144 <= 12'h989;
        src145 <= 12'h934;
        src146 <= 12'h9e;
        src147 <= 12'hcae;
        src148 <= 12'h93;
        src149 <= 12'hd54;
        src150 <= 12'haec;
        src151 <= 12'h83e;
        src152 <= 12'h5e6;
        src153 <= 12'h55a;
        src154 <= 12'hfc8;
        src155 <= 12'h6d7;
        src156 <= 12'h951;
        src157 <= 12'hf62;
        src158 <= 12'h397;
        src159 <= 12'hc7;
        src160 <= 12'h318;
        src161 <= 12'hc61;
        exp <= 20'h4bef3;
        #1
        src0 <= 12'h7ac;
        src1 <= 12'hd03;
        src2 <= 12'h51c;
        src3 <= 12'he16;
        src4 <= 12'h3dd;
        src5 <= 12'hf1f;
        src6 <= 12'h7e0;
        src7 <= 12'h53d;
        src8 <= 12'hd03;
        src9 <= 12'ha37;
        src10 <= 12'h13d;
        src11 <= 12'ha33;
        src12 <= 12'hc84;
        src13 <= 12'hb77;
        src14 <= 12'hf35;
        src15 <= 12'h9de;
        src16 <= 12'h593;
        src17 <= 12'h59a;
        src18 <= 12'hdc4;
        src19 <= 12'h3ed;
        src20 <= 12'hdcf;
        src21 <= 12'heb7;
        src22 <= 12'had1;
        src23 <= 12'h46f;
        src24 <= 12'h590;
        src25 <= 12'ha55;
        src26 <= 12'h5e7;
        src27 <= 12'h85a;
        src28 <= 12'hd2a;
        src29 <= 12'h3a0;
        src30 <= 12'h718;
        src31 <= 12'hbbf;
        src32 <= 12'h706;
        src33 <= 12'h61a;
        src34 <= 12'hc77;
        src35 <= 12'h2fe;
        src36 <= 12'h39c;
        src37 <= 12'h2b7;
        src38 <= 12'hc0;
        src39 <= 12'h50e;
        src40 <= 12'hea3;
        src41 <= 12'h87d;
        src42 <= 12'h986;
        src43 <= 12'h81b;
        src44 <= 12'hef;
        src45 <= 12'hc68;
        src46 <= 12'had6;
        src47 <= 12'hb84;
        src48 <= 12'h53;
        src49 <= 12'h520;
        src50 <= 12'hf84;
        src51 <= 12'h615;
        src52 <= 12'h646;
        src53 <= 12'hdbe;
        src54 <= 12'h1e3;
        src55 <= 12'hd00;
        src56 <= 12'h728;
        src57 <= 12'h4a4;
        src58 <= 12'h9e1;
        src59 <= 12'h508;
        src60 <= 12'h9b0;
        src61 <= 12'ha2e;
        src62 <= 12'h8e9;
        src63 <= 12'hfed;
        src64 <= 12'h6f0;
        src65 <= 12'h33c;
        src66 <= 12'hf4c;
        src67 <= 12'h553;
        src68 <= 12'h834;
        src69 <= 12'hb8;
        src70 <= 12'hdf4;
        src71 <= 12'h41a;
        src72 <= 12'hcb6;
        src73 <= 12'h36b;
        src74 <= 12'h29e;
        src75 <= 12'he30;
        src76 <= 12'h5c9;
        src77 <= 12'h226;
        src78 <= 12'hc76;
        src79 <= 12'hf23;
        src80 <= 12'h254;
        src81 <= 12'hf77;
        src82 <= 12'hc2;
        src83 <= 12'h55;
        src84 <= 12'h9d8;
        src85 <= 12'h663;
        src86 <= 12'h70e;
        src87 <= 12'h547;
        src88 <= 12'h3bc;
        src89 <= 12'hc86;
        src90 <= 12'hee3;
        src91 <= 12'he5e;
        src92 <= 12'h395;
        src93 <= 12'h74e;
        src94 <= 12'h846;
        src95 <= 12'h223;
        src96 <= 12'h94a;
        src97 <= 12'h88;
        src98 <= 12'h72e;
        src99 <= 12'h1af;
        src100 <= 12'h18c;
        src101 <= 12'h552;
        src102 <= 12'h9a0;
        src103 <= 12'h527;
        src104 <= 12'h41a;
        src105 <= 12'h2e8;
        src106 <= 12'h1e1;
        src107 <= 12'h9eb;
        src108 <= 12'h382;
        src109 <= 12'h56a;
        src110 <= 12'h6e7;
        src111 <= 12'h763;
        src112 <= 12'hf9c;
        src113 <= 12'he9d;
        src114 <= 12'hde1;
        src115 <= 12'h249;
        src116 <= 12'h616;
        src117 <= 12'h503;
        src118 <= 12'h679;
        src119 <= 12'h54b;
        src120 <= 12'h720;
        src121 <= 12'h313;
        src122 <= 12'hc1e;
        src123 <= 12'hdc7;
        src124 <= 12'h27c;
        src125 <= 12'h81f;
        src126 <= 12'hc38;
        src127 <= 12'h740;
        src128 <= 12'h3b6;
        src129 <= 12'h25f;
        src130 <= 12'h796;
        src131 <= 12'h5f4;
        src132 <= 12'h6c6;
        src133 <= 12'h93e;
        src134 <= 12'h6a3;
        src135 <= 12'he7;
        src136 <= 12'h4bd;
        src137 <= 12'h487;
        src138 <= 12'he22;
        src139 <= 12'h6d7;
        src140 <= 12'h4b3;
        src141 <= 12'h45f;
        src142 <= 12'hadb;
        src143 <= 12'hdae;
        src144 <= 12'h2d5;
        src145 <= 12'hf33;
        src146 <= 12'hf80;
        src147 <= 12'h5cf;
        src148 <= 12'h16a;
        src149 <= 12'h808;
        src150 <= 12'h65f;
        src151 <= 12'h24f;
        src152 <= 12'heef;
        src153 <= 12'h3ec;
        src154 <= 12'h707;
        src155 <= 12'h85;
        src156 <= 12'hfa;
        src157 <= 12'hbff;
        src158 <= 12'h5c4;
        src159 <= 12'hdaf;
        src160 <= 12'hb36;
        src161 <= 12'h1c8;
        exp <= 20'h4d72e;
        #1
        src0 <= 12'h533;
        src1 <= 12'h5eb;
        src2 <= 12'hc63;
        src3 <= 12'hff8;
        src4 <= 12'he5b;
        src5 <= 12'hb86;
        src6 <= 12'h9fe;
        src7 <= 12'h342;
        src8 <= 12'h9a2;
        src9 <= 12'h4bb;
        src10 <= 12'hfb0;
        src11 <= 12'h3da;
        src12 <= 12'haa6;
        src13 <= 12'h14e;
        src14 <= 12'hc50;
        src15 <= 12'h806;
        src16 <= 12'hfa1;
        src17 <= 12'he98;
        src18 <= 12'heb3;
        src19 <= 12'h5c0;
        src20 <= 12'hc9a;
        src21 <= 12'hc58;
        src22 <= 12'h49e;
        src23 <= 12'h445;
        src24 <= 12'h1e8;
        src25 <= 12'hf2c;
        src26 <= 12'head;
        src27 <= 12'hc74;
        src28 <= 12'hcf3;
        src29 <= 12'h8ae;
        src30 <= 12'hebf;
        src31 <= 12'h38b;
        src32 <= 12'h890;
        src33 <= 12'h410;
        src34 <= 12'h90a;
        src35 <= 12'hc0;
        src36 <= 12'h188;
        src37 <= 12'h98b;
        src38 <= 12'h5da;
        src39 <= 12'h3fe;
        src40 <= 12'hf84;
        src41 <= 12'h7b2;
        src42 <= 12'hdbd;
        src43 <= 12'h381;
        src44 <= 12'h1a6;
        src45 <= 12'hbcb;
        src46 <= 12'h271;
        src47 <= 12'h5ec;
        src48 <= 12'hd7d;
        src49 <= 12'h1c9;
        src50 <= 12'h8f;
        src51 <= 12'h2f1;
        src52 <= 12'ha33;
        src53 <= 12'hac9;
        src54 <= 12'h697;
        src55 <= 12'hc24;
        src56 <= 12'h34a;
        src57 <= 12'h8e5;
        src58 <= 12'h8c;
        src59 <= 12'h10e;
        src60 <= 12'ha23;
        src61 <= 12'hbf5;
        src62 <= 12'hdbb;
        src63 <= 12'h153;
        src64 <= 12'he22;
        src65 <= 12'hec3;
        src66 <= 12'hf70;
        src67 <= 12'ha79;
        src68 <= 12'h2da;
        src69 <= 12'h93e;
        src70 <= 12'hbe0;
        src71 <= 12'hdb1;
        src72 <= 12'h8fe;
        src73 <= 12'hd39;
        src74 <= 12'h91b;
        src75 <= 12'h39b;
        src76 <= 12'h9d1;
        src77 <= 12'h24c;
        src78 <= 12'h6d;
        src79 <= 12'h69e;
        src80 <= 12'hbfa;
        src81 <= 12'h94d;
        src82 <= 12'h63d;
        src83 <= 12'h751;
        src84 <= 12'h992;
        src85 <= 12'hc3;
        src86 <= 12'h2b;
        src87 <= 12'he60;
        src88 <= 12'h136;
        src89 <= 12'h86f;
        src90 <= 12'hcfc;
        src91 <= 12'h220;
        src92 <= 12'h517;
        src93 <= 12'h5f;
        src94 <= 12'h59;
        src95 <= 12'hbb6;
        src96 <= 12'h342;
        src97 <= 12'ha89;
        src98 <= 12'h96b;
        src99 <= 12'h5cc;
        src100 <= 12'h503;
        src101 <= 12'hb25;
        src102 <= 12'h115;
        src103 <= 12'h701;
        src104 <= 12'h287;
        src105 <= 12'h481;
        src106 <= 12'h6ed;
        src107 <= 12'h491;
        src108 <= 12'h2c;
        src109 <= 12'h4c2;
        src110 <= 12'h7ae;
        src111 <= 12'hc4b;
        src112 <= 12'h584;
        src113 <= 12'h53b;
        src114 <= 12'h102;
        src115 <= 12'he6a;
        src116 <= 12'h20a;
        src117 <= 12'h12d;
        src118 <= 12'h145;
        src119 <= 12'he1a;
        src120 <= 12'hb;
        src121 <= 12'h2f8;
        src122 <= 12'hb6d;
        src123 <= 12'h666;
        src124 <= 12'hc63;
        src125 <= 12'h228;
        src126 <= 12'ha17;
        src127 <= 12'h9d4;
        src128 <= 12'hcc9;
        src129 <= 12'he73;
        src130 <= 12'h237;
        src131 <= 12'h7f8;
        src132 <= 12'h157;
        src133 <= 12'hffe;
        src134 <= 12'h556;
        src135 <= 12'h378;
        src136 <= 12'h772;
        src137 <= 12'h7ad;
        src138 <= 12'hc84;
        src139 <= 12'h341;
        src140 <= 12'hade;
        src141 <= 12'he81;
        src142 <= 12'hd6f;
        src143 <= 12'h20f;
        src144 <= 12'haec;
        src145 <= 12'ha3a;
        src146 <= 12'hd73;
        src147 <= 12'hc96;
        src148 <= 12'h38c;
        src149 <= 12'h28;
        src150 <= 12'h1ae;
        src151 <= 12'h521;
        src152 <= 12'hbdf;
        src153 <= 12'he88;
        src154 <= 12'hb4e;
        src155 <= 12'h16f;
        src156 <= 12'h251;
        src157 <= 12'hf69;
        src158 <= 12'hff7;
        src159 <= 12'h7;
        src160 <= 12'h495;
        src161 <= 12'hdb5;
        exp <= 20'h4e9d7;
        #1
        src0 <= 12'h7ef;
        src1 <= 12'h5f3;
        src2 <= 12'hd2d;
        src3 <= 12'he9a;
        src4 <= 12'h799;
        src5 <= 12'he32;
        src6 <= 12'hc15;
        src7 <= 12'hca9;
        src8 <= 12'h8ba;
        src9 <= 12'he9a;
        src10 <= 12'hdc0;
        src11 <= 12'h8d1;
        src12 <= 12'hae5;
        src13 <= 12'hb8a;
        src14 <= 12'h86;
        src15 <= 12'h26;
        src16 <= 12'h703;
        src17 <= 12'h18f;
        src18 <= 12'h630;
        src19 <= 12'he92;
        src20 <= 12'hb5;
        src21 <= 12'hcaf;
        src22 <= 12'hc62;
        src23 <= 12'h830;
        src24 <= 12'h235;
        src25 <= 12'h12f;
        src26 <= 12'h752;
        src27 <= 12'h84a;
        src28 <= 12'h666;
        src29 <= 12'hb55;
        src30 <= 12'h482;
        src31 <= 12'h5a9;
        src32 <= 12'hdbb;
        src33 <= 12'had1;
        src34 <= 12'h217;
        src35 <= 12'h5a4;
        src36 <= 12'hbbe;
        src37 <= 12'h399;
        src38 <= 12'h2aa;
        src39 <= 12'h769;
        src40 <= 12'hb72;
        src41 <= 12'h8b5;
        src42 <= 12'h219;
        src43 <= 12'h802;
        src44 <= 12'hb3;
        src45 <= 12'hb6c;
        src46 <= 12'h133;
        src47 <= 12'hc0;
        src48 <= 12'he34;
        src49 <= 12'he80;
        src50 <= 12'h87e;
        src51 <= 12'h7b9;
        src52 <= 12'h55c;
        src53 <= 12'h631;
        src54 <= 12'he1e;
        src55 <= 12'ha33;
        src56 <= 12'hbd5;
        src57 <= 12'hd4f;
        src58 <= 12'h3d7;
        src59 <= 12'h470;
        src60 <= 12'h607;
        src61 <= 12'h853;
        src62 <= 12'hbb8;
        src63 <= 12'h620;
        src64 <= 12'hb0e;
        src65 <= 12'h6dd;
        src66 <= 12'h91b;
        src67 <= 12'hc5e;
        src68 <= 12'h792;
        src69 <= 12'h998;
        src70 <= 12'hb55;
        src71 <= 12'h2a2;
        src72 <= 12'h8d1;
        src73 <= 12'h6cc;
        src74 <= 12'hc12;
        src75 <= 12'h26b;
        src76 <= 12'hc43;
        src77 <= 12'hbf8;
        src78 <= 12'h10e;
        src79 <= 12'h525;
        src80 <= 12'h8ac;
        src81 <= 12'ha0f;
        src82 <= 12'h46e;
        src83 <= 12'h189;
        src84 <= 12'h209;
        src85 <= 12'h9e8;
        src86 <= 12'h446;
        src87 <= 12'hbc0;
        src88 <= 12'h955;
        src89 <= 12'h671;
        src90 <= 12'hd98;
        src91 <= 12'h69a;
        src92 <= 12'h776;
        src93 <= 12'hb40;
        src94 <= 12'h10d;
        src95 <= 12'hfb1;
        src96 <= 12'h518;
        src97 <= 12'hca9;
        src98 <= 12'h18;
        src99 <= 12'hc2a;
        src100 <= 12'h7f7;
        src101 <= 12'h6b4;
        src102 <= 12'hdff;
        src103 <= 12'h23d;
        src104 <= 12'h898;
        src105 <= 12'h7f9;
        src106 <= 12'h11e;
        src107 <= 12'hfd5;
        src108 <= 12'h457;
        src109 <= 12'hbe3;
        src110 <= 12'h6f4;
        src111 <= 12'hc09;
        src112 <= 12'ha66;
        src113 <= 12'hea3;
        src114 <= 12'hf5f;
        src115 <= 12'hdd8;
        src116 <= 12'h3de;
        src117 <= 12'h8f9;
        src118 <= 12'h6eb;
        src119 <= 12'h20a;
        src120 <= 12'h6e2;
        src121 <= 12'hdbb;
        src122 <= 12'h3dc;
        src123 <= 12'hf5d;
        src124 <= 12'h1af;
        src125 <= 12'h8fd;
        src126 <= 12'h4c9;
        src127 <= 12'h98f;
        src128 <= 12'h1af;
        src129 <= 12'h458;
        src130 <= 12'hc9;
        src131 <= 12'h68c;
        src132 <= 12'h97f;
        src133 <= 12'h475;
        src134 <= 12'h75d;
        src135 <= 12'h704;
        src136 <= 12'h4fa;
        src137 <= 12'hf81;
        src138 <= 12'hcb4;
        src139 <= 12'h688;
        src140 <= 12'hf31;
        src141 <= 12'hde0;
        src142 <= 12'h417;
        src143 <= 12'h251;
        src144 <= 12'hf17;
        src145 <= 12'h341;
        src146 <= 12'hc8f;
        src147 <= 12'he5e;
        src148 <= 12'h283;
        src149 <= 12'hf99;
        src150 <= 12'h866;
        src151 <= 12'h82b;
        src152 <= 12'h713;
        src153 <= 12'h55c;
        src154 <= 12'h860;
        src155 <= 12'he5;
        src156 <= 12'ha7a;
        src157 <= 12'h8f5;
        src158 <= 12'h334;
        src159 <= 12'h993;
        src160 <= 12'hcb6;
        src161 <= 12'h120;
        exp <= 20'h51a0d;
        #1
        src0 <= 12'ha5e;
        src1 <= 12'h31f;
        src2 <= 12'h547;
        src3 <= 12'h8;
        src4 <= 12'h628;
        src5 <= 12'h91d;
        src6 <= 12'heee;
        src7 <= 12'h324;
        src8 <= 12'h719;
        src9 <= 12'hd04;
        src10 <= 12'hb7a;
        src11 <= 12'hde8;
        src12 <= 12'h13e;
        src13 <= 12'h386;
        src14 <= 12'hd36;
        src15 <= 12'h830;
        src16 <= 12'h2cd;
        src17 <= 12'h69b;
        src18 <= 12'h2e8;
        src19 <= 12'haf6;
        src20 <= 12'h150;
        src21 <= 12'h896;
        src22 <= 12'h474;
        src23 <= 12'ha2d;
        src24 <= 12'hc08;
        src25 <= 12'he86;
        src26 <= 12'h53f;
        src27 <= 12'h3bc;
        src28 <= 12'h213;
        src29 <= 12'hbae;
        src30 <= 12'h25f;
        src31 <= 12'h1b0;
        src32 <= 12'h41f;
        src33 <= 12'h825;
        src34 <= 12'hf12;
        src35 <= 12'h9a1;
        src36 <= 12'h52e;
        src37 <= 12'ha26;
        src38 <= 12'h19e;
        src39 <= 12'hee5;
        src40 <= 12'h98f;
        src41 <= 12'hd9;
        src42 <= 12'haaa;
        src43 <= 12'h16;
        src44 <= 12'h95e;
        src45 <= 12'h662;
        src46 <= 12'h447;
        src47 <= 12'h504;
        src48 <= 12'h49;
        src49 <= 12'hde7;
        src50 <= 12'h4d6;
        src51 <= 12'h95a;
        src52 <= 12'hd24;
        src53 <= 12'h1b3;
        src54 <= 12'h9d5;
        src55 <= 12'h2be;
        src56 <= 12'hc2c;
        src57 <= 12'hccf;
        src58 <= 12'hcbb;
        src59 <= 12'haa4;
        src60 <= 12'he52;
        src61 <= 12'h764;
        src62 <= 12'hd3f;
        src63 <= 12'h557;
        src64 <= 12'h8cc;
        src65 <= 12'hec2;
        src66 <= 12'ha80;
        src67 <= 12'hcb5;
        src68 <= 12'h6c2;
        src69 <= 12'hd49;
        src70 <= 12'h2b5;
        src71 <= 12'h659;
        src72 <= 12'h937;
        src73 <= 12'ha05;
        src74 <= 12'h14a;
        src75 <= 12'h732;
        src76 <= 12'ha32;
        src77 <= 12'h6c2;
        src78 <= 12'hf34;
        src79 <= 12'h865;
        src80 <= 12'hdf1;
        src81 <= 12'hb82;
        src82 <= 12'h83e;
        src83 <= 12'h5b3;
        src84 <= 12'h3b9;
        src85 <= 12'h6c7;
        src86 <= 12'h6a;
        src87 <= 12'hdb4;
        src88 <= 12'hc4a;
        src89 <= 12'h761;
        src90 <= 12'h8e0;
        src91 <= 12'h5e8;
        src92 <= 12'h704;
        src93 <= 12'hb34;
        src94 <= 12'h35a;
        src95 <= 12'h3a4;
        src96 <= 12'h8c5;
        src97 <= 12'hf1f;
        src98 <= 12'h999;
        src99 <= 12'h5eb;
        src100 <= 12'he2f;
        src101 <= 12'hf59;
        src102 <= 12'hbcc;
        src103 <= 12'h966;
        src104 <= 12'h98f;
        src105 <= 12'ha3c;
        src106 <= 12'h1a3;
        src107 <= 12'h973;
        src108 <= 12'h32b;
        src109 <= 12'hc4c;
        src110 <= 12'ha0b;
        src111 <= 12'ha4c;
        src112 <= 12'hfcf;
        src113 <= 12'h56c;
        src114 <= 12'ha6a;
        src115 <= 12'hd47;
        src116 <= 12'h1c6;
        src117 <= 12'hdc2;
        src118 <= 12'hd83;
        src119 <= 12'h13d;
        src120 <= 12'hfa7;
        src121 <= 12'h9a8;
        src122 <= 12'he15;
        src123 <= 12'hdee;
        src124 <= 12'h33;
        src125 <= 12'hcf6;
        src126 <= 12'hf75;
        src127 <= 12'hf7b;
        src128 <= 12'hd6d;
        src129 <= 12'ha16;
        src130 <= 12'h9;
        src131 <= 12'haf3;
        src132 <= 12'hc6f;
        src133 <= 12'ha5c;
        src134 <= 12'h6d9;
        src135 <= 12'hcdb;
        src136 <= 12'h27;
        src137 <= 12'hf2e;
        src138 <= 12'h663;
        src139 <= 12'hb4a;
        src140 <= 12'h63d;
        src141 <= 12'h661;
        src142 <= 12'h806;
        src143 <= 12'hcba;
        src144 <= 12'ha97;
        src145 <= 12'h590;
        src146 <= 12'had1;
        src147 <= 12'h7e4;
        src148 <= 12'hd9a;
        src149 <= 12'h99f;
        src150 <= 12'hc3d;
        src151 <= 12'h22;
        src152 <= 12'hf0c;
        src153 <= 12'hcd8;
        src154 <= 12'hcd7;
        src155 <= 12'h98b;
        src156 <= 12'h167;
        src157 <= 12'h1ae;
        src158 <= 12'h552;
        src159 <= 12'he30;
        src160 <= 12'hd67;
        src161 <= 12'h6d1;
        exp <= 20'h56c86;
        #1
        src0 <= 12'h73e;
        src1 <= 12'h729;
        src2 <= 12'hc9e;
        src3 <= 12'haf;
        src4 <= 12'h665;
        src5 <= 12'h14;
        src6 <= 12'hb4d;
        src7 <= 12'he14;
        src8 <= 12'hdd6;
        src9 <= 12'haca;
        src10 <= 12'ha2c;
        src11 <= 12'h517;
        src12 <= 12'h5d;
        src13 <= 12'ha18;
        src14 <= 12'h249;
        src15 <= 12'h64e;
        src16 <= 12'h5cb;
        src17 <= 12'h74a;
        src18 <= 12'h64;
        src19 <= 12'hbb5;
        src20 <= 12'hb8c;
        src21 <= 12'hf49;
        src22 <= 12'h5bb;
        src23 <= 12'hcc2;
        src24 <= 12'hbe7;
        src25 <= 12'hbc6;
        src26 <= 12'he36;
        src27 <= 12'h44d;
        src28 <= 12'h417;
        src29 <= 12'hd01;
        src30 <= 12'h71c;
        src31 <= 12'hb85;
        src32 <= 12'h641;
        src33 <= 12'h89e;
        src34 <= 12'h42d;
        src35 <= 12'hbc8;
        src36 <= 12'h48a;
        src37 <= 12'h268;
        src38 <= 12'h29e;
        src39 <= 12'h6a5;
        src40 <= 12'h8c3;
        src41 <= 12'hf1b;
        src42 <= 12'hd72;
        src43 <= 12'h3fb;
        src44 <= 12'h7a5;
        src45 <= 12'h722;
        src46 <= 12'h9ef;
        src47 <= 12'h710;
        src48 <= 12'h1a1;
        src49 <= 12'h376;
        src50 <= 12'he9a;
        src51 <= 12'h45c;
        src52 <= 12'hd5f;
        src53 <= 12'hd0f;
        src54 <= 12'h3b4;
        src55 <= 12'h49b;
        src56 <= 12'hd92;
        src57 <= 12'hea;
        src58 <= 12'hb35;
        src59 <= 12'h5dc;
        src60 <= 12'h249;
        src61 <= 12'hcdd;
        src62 <= 12'h293;
        src63 <= 12'h11f;
        src64 <= 12'h16d;
        src65 <= 12'h83e;
        src66 <= 12'h8a8;
        src67 <= 12'hec5;
        src68 <= 12'hf34;
        src69 <= 12'h234;
        src70 <= 12'h1c5;
        src71 <= 12'h9a9;
        src72 <= 12'hc0c;
        src73 <= 12'he6b;
        src74 <= 12'h968;
        src75 <= 12'h332;
        src76 <= 12'had7;
        src77 <= 12'h949;
        src78 <= 12'h16c;
        src79 <= 12'hdd6;
        src80 <= 12'ha73;
        src81 <= 12'hf25;
        src82 <= 12'hfa5;
        src83 <= 12'h400;
        src84 <= 12'h703;
        src85 <= 12'h100;
        src86 <= 12'hcde;
        src87 <= 12'h907;
        src88 <= 12'h8b;
        src89 <= 12'h4c8;
        src90 <= 12'h8ac;
        src91 <= 12'h436;
        src92 <= 12'hc5a;
        src93 <= 12'h6bd;
        src94 <= 12'hd73;
        src95 <= 12'hbd4;
        src96 <= 12'h5d1;
        src97 <= 12'he33;
        src98 <= 12'h696;
        src99 <= 12'hf0;
        src100 <= 12'hea3;
        src101 <= 12'heca;
        src102 <= 12'ha41;
        src103 <= 12'h6b7;
        src104 <= 12'hc9f;
        src105 <= 12'h330;
        src106 <= 12'hec;
        src107 <= 12'h380;
        src108 <= 12'h19;
        src109 <= 12'h80f;
        src110 <= 12'h153;
        src111 <= 12'h46b;
        src112 <= 12'hd83;
        src113 <= 12'hba1;
        src114 <= 12'hae5;
        src115 <= 12'h9cd;
        src116 <= 12'h3f2;
        src117 <= 12'hab2;
        src118 <= 12'h9ea;
        src119 <= 12'h43a;
        src120 <= 12'ha3;
        src121 <= 12'h3b;
        src122 <= 12'hb88;
        src123 <= 12'h4d2;
        src124 <= 12'hf91;
        src125 <= 12'h6e2;
        src126 <= 12'h21e;
        src127 <= 12'h465;
        src128 <= 12'hea0;
        src129 <= 12'h10a;
        src130 <= 12'h689;
        src131 <= 12'hd07;
        src132 <= 12'h3d7;
        src133 <= 12'hb04;
        src134 <= 12'ha6c;
        src135 <= 12'h9a7;
        src136 <= 12'h29d;
        src137 <= 12'h6e0;
        src138 <= 12'hde0;
        src139 <= 12'hd74;
        src140 <= 12'h519;
        src141 <= 12'ha7b;
        src142 <= 12'hf93;
        src143 <= 12'h1c7;
        src144 <= 12'h45c;
        src145 <= 12'h1c5;
        src146 <= 12'h77b;
        src147 <= 12'h911;
        src148 <= 12'ha51;
        src149 <= 12'ha38;
        src150 <= 12'h1b3;
        src151 <= 12'h3f4;
        src152 <= 12'h236;
        src153 <= 12'h1e0;
        src154 <= 12'h6d4;
        src155 <= 12'h243;
        src156 <= 12'hbb;
        src157 <= 12'h206;
        src158 <= 12'hfa2;
        src159 <= 12'hd0;
        src160 <= 12'h73c;
        src161 <= 12'h4e5;
        exp <= 20'h4d069;
        #1
        src0 <= 12'h90;
        src1 <= 12'h383;
        src2 <= 12'hf79;
        src3 <= 12'hd2d;
        src4 <= 12'hb33;
        src5 <= 12'hf35;
        src6 <= 12'hcd6;
        src7 <= 12'h48a;
        src8 <= 12'h14b;
        src9 <= 12'hc54;
        src10 <= 12'h2cb;
        src11 <= 12'hff7;
        src12 <= 12'h689;
        src13 <= 12'h649;
        src14 <= 12'hbd2;
        src15 <= 12'h6e3;
        src16 <= 12'h4bb;
        src17 <= 12'h227;
        src18 <= 12'hdc7;
        src19 <= 12'h883;
        src20 <= 12'h9f9;
        src21 <= 12'h7ed;
        src22 <= 12'hb63;
        src23 <= 12'hd2;
        src24 <= 12'h921;
        src25 <= 12'h8d6;
        src26 <= 12'h61b;
        src27 <= 12'h443;
        src28 <= 12'h544;
        src29 <= 12'hf58;
        src30 <= 12'h558;
        src31 <= 12'h12;
        src32 <= 12'h81b;
        src33 <= 12'hfd2;
        src34 <= 12'h383;
        src35 <= 12'hcba;
        src36 <= 12'heed;
        src37 <= 12'he60;
        src38 <= 12'h117;
        src39 <= 12'hd25;
        src40 <= 12'h190;
        src41 <= 12'h458;
        src42 <= 12'hbc0;
        src43 <= 12'h653;
        src44 <= 12'h1aa;
        src45 <= 12'h9d9;
        src46 <= 12'hb9;
        src47 <= 12'hcb8;
        src48 <= 12'h689;
        src49 <= 12'h10a;
        src50 <= 12'h6f8;
        src51 <= 12'hbdc;
        src52 <= 12'h76b;
        src53 <= 12'hb68;
        src54 <= 12'hd1c;
        src55 <= 12'h63d;
        src56 <= 12'h9bb;
        src57 <= 12'hb5;
        src58 <= 12'hc6c;
        src59 <= 12'h918;
        src60 <= 12'h2cf;
        src61 <= 12'h4c0;
        src62 <= 12'h40e;
        src63 <= 12'hb1c;
        src64 <= 12'hc2c;
        src65 <= 12'h46f;
        src66 <= 12'h3fc;
        src67 <= 12'hb49;
        src68 <= 12'h16f;
        src69 <= 12'h2d3;
        src70 <= 12'h4ff;
        src71 <= 12'h3ce;
        src72 <= 12'h1a5;
        src73 <= 12'h121;
        src74 <= 12'h223;
        src75 <= 12'h3e0;
        src76 <= 12'hf4a;
        src77 <= 12'hbc7;
        src78 <= 12'h6b;
        src79 <= 12'h3ff;
        src80 <= 12'habb;
        src81 <= 12'h8a4;
        src82 <= 12'hd02;
        src83 <= 12'h924;
        src84 <= 12'hdaf;
        src85 <= 12'h21e;
        src86 <= 12'h2f6;
        src87 <= 12'h863;
        src88 <= 12'h815;
        src89 <= 12'heb5;
        src90 <= 12'h600;
        src91 <= 12'h5bf;
        src92 <= 12'h41e;
        src93 <= 12'h5c;
        src94 <= 12'h86f;
        src95 <= 12'hf29;
        src96 <= 12'h580;
        src97 <= 12'h495;
        src98 <= 12'hff4;
        src99 <= 12'h894;
        src100 <= 12'hdec;
        src101 <= 12'h9f0;
        src102 <= 12'hde4;
        src103 <= 12'hdfa;
        src104 <= 12'h89e;
        src105 <= 12'he92;
        src106 <= 12'h262;
        src107 <= 12'h704;
        src108 <= 12'h347;
        src109 <= 12'had4;
        src110 <= 12'h654;
        src111 <= 12'hcba;
        src112 <= 12'h152;
        src113 <= 12'h283;
        src114 <= 12'h9b8;
        src115 <= 12'h7e1;
        src116 <= 12'h339;
        src117 <= 12'h69e;
        src118 <= 12'h5fd;
        src119 <= 12'hcd3;
        src120 <= 12'hc9b;
        src121 <= 12'hda;
        src122 <= 12'ha2;
        src123 <= 12'h389;
        src124 <= 12'h4a9;
        src125 <= 12'h94;
        src126 <= 12'h644;
        src127 <= 12'h678;
        src128 <= 12'h294;
        src129 <= 12'h80b;
        src130 <= 12'hd1c;
        src131 <= 12'h49f;
        src132 <= 12'h4af;
        src133 <= 12'hdad;
        src134 <= 12'h48;
        src135 <= 12'hffd;
        src136 <= 12'h1ad;
        src137 <= 12'hd27;
        src138 <= 12'hf3d;
        src139 <= 12'h7a1;
        src140 <= 12'h522;
        src141 <= 12'h372;
        src142 <= 12'h202;
        src143 <= 12'hdcd;
        src144 <= 12'h23c;
        src145 <= 12'he4a;
        src146 <= 12'hf2b;
        src147 <= 12'h30c;
        src148 <= 12'hf93;
        src149 <= 12'h790;
        src150 <= 12'he25;
        src151 <= 12'hec7;
        src152 <= 12'h8bf;
        src153 <= 12'h3d8;
        src154 <= 12'h793;
        src155 <= 12'hcf9;
        src156 <= 12'h975;
        src157 <= 12'h329;
        src158 <= 12'hb6f;
        src159 <= 12'h566;
        src160 <= 12'hdcd;
        src161 <= 12'hd89;
        exp <= 20'h4edf2;
        #1
        src0 <= 12'h87a;
        src1 <= 12'h1e4;
        src2 <= 12'hb5;
        src3 <= 12'hdd;
        src4 <= 12'h95d;
        src5 <= 12'hde2;
        src6 <= 12'hfc4;
        src7 <= 12'h7af;
        src8 <= 12'hf4f;
        src9 <= 12'h328;
        src10 <= 12'h2ab;
        src11 <= 12'h48b;
        src12 <= 12'hc43;
        src13 <= 12'h50c;
        src14 <= 12'h4be;
        src15 <= 12'h8bc;
        src16 <= 12'hf87;
        src17 <= 12'h53b;
        src18 <= 12'h999;
        src19 <= 12'h436;
        src20 <= 12'hade;
        src21 <= 12'h8a;
        src22 <= 12'h99;
        src23 <= 12'h946;
        src24 <= 12'h4ee;
        src25 <= 12'hb4b;
        src26 <= 12'h4a5;
        src27 <= 12'h3d;
        src28 <= 12'h20c;
        src29 <= 12'hcef;
        src30 <= 12'h8e1;
        src31 <= 12'hd4a;
        src32 <= 12'hdab;
        src33 <= 12'h9c2;
        src34 <= 12'hfc0;
        src35 <= 12'h30;
        src36 <= 12'h71d;
        src37 <= 12'h7ba;
        src38 <= 12'hf1a;
        src39 <= 12'h8db;
        src40 <= 12'h1d8;
        src41 <= 12'hb9d;
        src42 <= 12'hd72;
        src43 <= 12'h2ca;
        src44 <= 12'h54;
        src45 <= 12'hde5;
        src46 <= 12'h29e;
        src47 <= 12'hd37;
        src48 <= 12'h6fb;
        src49 <= 12'hce7;
        src50 <= 12'h483;
        src51 <= 12'h75a;
        src52 <= 12'h937;
        src53 <= 12'hd37;
        src54 <= 12'ha16;
        src55 <= 12'h89c;
        src56 <= 12'hc6c;
        src57 <= 12'hb70;
        src58 <= 12'h946;
        src59 <= 12'hed2;
        src60 <= 12'h628;
        src61 <= 12'h142;
        src62 <= 12'h43b;
        src63 <= 12'h2f3;
        src64 <= 12'hc5f;
        src65 <= 12'h6f7;
        src66 <= 12'h3ee;
        src67 <= 12'h2a;
        src68 <= 12'h86f;
        src69 <= 12'h7d3;
        src70 <= 12'hc47;
        src71 <= 12'h6ac;
        src72 <= 12'h791;
        src73 <= 12'hbe3;
        src74 <= 12'hda2;
        src75 <= 12'hc5c;
        src76 <= 12'h1cb;
        src77 <= 12'h77f;
        src78 <= 12'h26c;
        src79 <= 12'h663;
        src80 <= 12'hba6;
        src81 <= 12'hc5f;
        src82 <= 12'h65a;
        src83 <= 12'heec;
        src84 <= 12'h852;
        src85 <= 12'hfd2;
        src86 <= 12'hfd5;
        src87 <= 12'hd6a;
        src88 <= 12'had8;
        src89 <= 12'h2ad;
        src90 <= 12'h961;
        src91 <= 12'hea5;
        src92 <= 12'h547;
        src93 <= 12'hbb4;
        src94 <= 12'h7a3;
        src95 <= 12'hbd3;
        src96 <= 12'h6fe;
        src97 <= 12'hafc;
        src98 <= 12'hd84;
        src99 <= 12'hf26;
        src100 <= 12'h505;
        src101 <= 12'h4e1;
        src102 <= 12'h50;
        src103 <= 12'ha54;
        src104 <= 12'hfe2;
        src105 <= 12'hb4d;
        src106 <= 12'h807;
        src107 <= 12'h61c;
        src108 <= 12'hefd;
        src109 <= 12'h2ff;
        src110 <= 12'ha86;
        src111 <= 12'hb10;
        src112 <= 12'h383;
        src113 <= 12'h98a;
        src114 <= 12'hf17;
        src115 <= 12'h868;
        src116 <= 12'h60f;
        src117 <= 12'h5de;
        src118 <= 12'h673;
        src119 <= 12'h7fb;
        src120 <= 12'h924;
        src121 <= 12'h608;
        src122 <= 12'h37a;
        src123 <= 12'haf0;
        src124 <= 12'h4;
        src125 <= 12'h9e6;
        src126 <= 12'h9c;
        src127 <= 12'h8c5;
        src128 <= 12'ha20;
        src129 <= 12'h665;
        src130 <= 12'heb9;
        src131 <= 12'h55f;
        src132 <= 12'hd9e;
        src133 <= 12'hebf;
        src134 <= 12'hf38;
        src135 <= 12'h4d6;
        src136 <= 12'h6ea;
        src137 <= 12'h512;
        src138 <= 12'hd44;
        src139 <= 12'h9c;
        src140 <= 12'h79;
        src141 <= 12'h189;
        src142 <= 12'h353;
        src143 <= 12'h4a4;
        src144 <= 12'hbf;
        src145 <= 12'h78;
        src146 <= 12'h8a0;
        src147 <= 12'h951;
        src148 <= 12'hefb;
        src149 <= 12'h8f9;
        src150 <= 12'heed;
        src151 <= 12'ha6;
        src152 <= 12'he88;
        src153 <= 12'hc4e;
        src154 <= 12'hfa4;
        src155 <= 12'ha04;
        src156 <= 12'h533;
        src157 <= 12'h146;
        src158 <= 12'he09;
        src159 <= 12'hc76;
        src160 <= 12'h79;
        src161 <= 12'hf22;
        exp <= 20'h539d3;
        #1
        src0 <= 12'h7f5;
        src1 <= 12'h869;
        src2 <= 12'h61;
        src3 <= 12'h9fe;
        src4 <= 12'hd28;
        src5 <= 12'hcd5;
        src6 <= 12'hbb4;
        src7 <= 12'hdaa;
        src8 <= 12'h16e;
        src9 <= 12'h818;
        src10 <= 12'h47f;
        src11 <= 12'hdf1;
        src12 <= 12'h7c5;
        src13 <= 12'h6f9;
        src14 <= 12'h6db;
        src15 <= 12'hea0;
        src16 <= 12'h8f3;
        src17 <= 12'hd4d;
        src18 <= 12'h3cd;
        src19 <= 12'hb59;
        src20 <= 12'h8f4;
        src21 <= 12'h9e0;
        src22 <= 12'hadd;
        src23 <= 12'h34f;
        src24 <= 12'hd54;
        src25 <= 12'h8c5;
        src26 <= 12'h730;
        src27 <= 12'h215;
        src28 <= 12'he14;
        src29 <= 12'hf30;
        src30 <= 12'h7e3;
        src31 <= 12'ha48;
        src32 <= 12'hff;
        src33 <= 12'h9f5;
        src34 <= 12'ha03;
        src35 <= 12'h409;
        src36 <= 12'hb0e;
        src37 <= 12'he4b;
        src38 <= 12'h8de;
        src39 <= 12'hdf1;
        src40 <= 12'hdf3;
        src41 <= 12'h125;
        src42 <= 12'h2a7;
        src43 <= 12'h13c;
        src44 <= 12'h78c;
        src45 <= 12'hd57;
        src46 <= 12'h46d;
        src47 <= 12'h76a;
        src48 <= 12'hf93;
        src49 <= 12'h195;
        src50 <= 12'h344;
        src51 <= 12'h2d5;
        src52 <= 12'hc7;
        src53 <= 12'h3a2;
        src54 <= 12'h2ff;
        src55 <= 12'h3ce;
        src56 <= 12'h256;
        src57 <= 12'hee4;
        src58 <= 12'ha97;
        src59 <= 12'h83a;
        src60 <= 12'h2e;
        src61 <= 12'he2c;
        src62 <= 12'he17;
        src63 <= 12'hf8c;
        src64 <= 12'hff2;
        src65 <= 12'he47;
        src66 <= 12'hf1;
        src67 <= 12'ha3d;
        src68 <= 12'h62b;
        src69 <= 12'h8ac;
        src70 <= 12'hba4;
        src71 <= 12'hb70;
        src72 <= 12'hded;
        src73 <= 12'h7ce;
        src74 <= 12'h617;
        src75 <= 12'h1c1;
        src76 <= 12'h331;
        src77 <= 12'hb4c;
        src78 <= 12'hc88;
        src79 <= 12'hbda;
        src80 <= 12'hc5a;
        src81 <= 12'h121;
        src82 <= 12'hdb8;
        src83 <= 12'hd93;
        src84 <= 12'h960;
        src85 <= 12'h577;
        src86 <= 12'hd7b;
        src87 <= 12'h2d0;
        src88 <= 12'ha33;
        src89 <= 12'h908;
        src90 <= 12'h787;
        src91 <= 12'hd38;
        src92 <= 12'hd34;
        src93 <= 12'h5ec;
        src94 <= 12'hd9;
        src95 <= 12'h850;
        src96 <= 12'hc;
        src97 <= 12'h7e0;
        src98 <= 12'hc72;
        src99 <= 12'h2bd;
        src100 <= 12'h9f7;
        src101 <= 12'he7f;
        src102 <= 12'hf1e;
        src103 <= 12'hdfa;
        src104 <= 12'hb93;
        src105 <= 12'hb55;
        src106 <= 12'h1df;
        src107 <= 12'h7b7;
        src108 <= 12'hf17;
        src109 <= 12'hc73;
        src110 <= 12'h303;
        src111 <= 12'h132;
        src112 <= 12'hf46;
        src113 <= 12'h921;
        src114 <= 12'h473;
        src115 <= 12'hca;
        src116 <= 12'hae6;
        src117 <= 12'h9ce;
        src118 <= 12'h56e;
        src119 <= 12'hae6;
        src120 <= 12'h1ff;
        src121 <= 12'h548;
        src122 <= 12'hd0e;
        src123 <= 12'h3ee;
        src124 <= 12'h792;
        src125 <= 12'hac0;
        src126 <= 12'hbe5;
        src127 <= 12'h527;
        src128 <= 12'hc78;
        src129 <= 12'h7b4;
        src130 <= 12'h9c3;
        src131 <= 12'h1eb;
        src132 <= 12'h1e5;
        src133 <= 12'hacc;
        src134 <= 12'h993;
        src135 <= 12'h898;
        src136 <= 12'h1ac;
        src137 <= 12'h1b4;
        src138 <= 12'h51;
        src139 <= 12'hfbc;
        src140 <= 12'h9f1;
        src141 <= 12'hff1;
        src142 <= 12'h3da;
        src143 <= 12'h6f5;
        src144 <= 12'h472;
        src145 <= 12'ha97;
        src146 <= 12'hd69;
        src147 <= 12'h35e;
        src148 <= 12'hdee;
        src149 <= 12'h83c;
        src150 <= 12'h98d;
        src151 <= 12'h5a;
        src152 <= 12'hc0a;
        src153 <= 12'h9e;
        src154 <= 12'h3df;
        src155 <= 12'h9da;
        src156 <= 12'h7cf;
        src157 <= 12'hb3f;
        src158 <= 12'h2ad;
        src159 <= 12'hb9f;
        src160 <= 12'h856;
        src161 <= 12'hefa;
        exp <= 20'h547b8;
        #1
        src0 <= 12'h991;
        src1 <= 12'hd53;
        src2 <= 12'h690;
        src3 <= 12'ha68;
        src4 <= 12'h75c;
        src5 <= 12'h943;
        src6 <= 12'h7d2;
        src7 <= 12'h598;
        src8 <= 12'h7f6;
        src9 <= 12'h8a;
        src10 <= 12'h4cc;
        src11 <= 12'hc17;
        src12 <= 12'he8d;
        src13 <= 12'hbce;
        src14 <= 12'hf60;
        src15 <= 12'h9e5;
        src16 <= 12'hd66;
        src17 <= 12'h758;
        src18 <= 12'hfa3;
        src19 <= 12'h336;
        src20 <= 12'h6d1;
        src21 <= 12'h26b;
        src22 <= 12'ha7a;
        src23 <= 12'he0c;
        src24 <= 12'hd74;
        src25 <= 12'h760;
        src26 <= 12'haa7;
        src27 <= 12'h5a6;
        src28 <= 12'h63b;
        src29 <= 12'h775;
        src30 <= 12'hb61;
        src31 <= 12'h7b0;
        src32 <= 12'he51;
        src33 <= 12'hf17;
        src34 <= 12'he7f;
        src35 <= 12'h34;
        src36 <= 12'h843;
        src37 <= 12'h433;
        src38 <= 12'h986;
        src39 <= 12'h500;
        src40 <= 12'h407;
        src41 <= 12'hef0;
        src42 <= 12'hf53;
        src43 <= 12'h7c8;
        src44 <= 12'h126;
        src45 <= 12'h53b;
        src46 <= 12'h2fc;
        src47 <= 12'ha1d;
        src48 <= 12'h9a7;
        src49 <= 12'he30;
        src50 <= 12'h4a6;
        src51 <= 12'h371;
        src52 <= 12'ha9a;
        src53 <= 12'hef3;
        src54 <= 12'hac3;
        src55 <= 12'hbe5;
        src56 <= 12'h746;
        src57 <= 12'h1db;
        src58 <= 12'hd2e;
        src59 <= 12'hcc2;
        src60 <= 12'hc3c;
        src61 <= 12'h9ff;
        src62 <= 12'hf57;
        src63 <= 12'h686;
        src64 <= 12'ha90;
        src65 <= 12'hc59;
        src66 <= 12'ha6;
        src67 <= 12'h842;
        src68 <= 12'h186;
        src69 <= 12'h54;
        src70 <= 12'h675;
        src71 <= 12'he41;
        src72 <= 12'ha8d;
        src73 <= 12'h13d;
        src74 <= 12'h53c;
        src75 <= 12'hbcd;
        src76 <= 12'hef6;
        src77 <= 12'h44f;
        src78 <= 12'h5ed;
        src79 <= 12'he09;
        src80 <= 12'h3f0;
        src81 <= 12'h7af;
        src82 <= 12'h627;
        src83 <= 12'hd00;
        src84 <= 12'h681;
        src85 <= 12'hfbf;
        src86 <= 12'h982;
        src87 <= 12'hf0b;
        src88 <= 12'h729;
        src89 <= 12'hcb7;
        src90 <= 12'ha50;
        src91 <= 12'hb56;
        src92 <= 12'h4a1;
        src93 <= 12'ha03;
        src94 <= 12'h3;
        src95 <= 12'hec5;
        src96 <= 12'h664;
        src97 <= 12'ha25;
        src98 <= 12'h453;
        src99 <= 12'h75b;
        src100 <= 12'hb7e;
        src101 <= 12'h839;
        src102 <= 12'h37d;
        src103 <= 12'h491;
        src104 <= 12'hafc;
        src105 <= 12'h459;
        src106 <= 12'h5e3;
        src107 <= 12'h26e;
        src108 <= 12'h860;
        src109 <= 12'h917;
        src110 <= 12'hae1;
        src111 <= 12'h14b;
        src112 <= 12'h476;
        src113 <= 12'h90c;
        src114 <= 12'ha7a;
        src115 <= 12'hc74;
        src116 <= 12'h964;
        src117 <= 12'hab5;
        src118 <= 12'h894;
        src119 <= 12'h165;
        src120 <= 12'ha1e;
        src121 <= 12'h484;
        src122 <= 12'h4f6;
        src123 <= 12'h96e;
        src124 <= 12'h98c;
        src125 <= 12'h6b5;
        src126 <= 12'h351;
        src127 <= 12'h66;
        src128 <= 12'h387;
        src129 <= 12'h200;
        src130 <= 12'ha0c;
        src131 <= 12'hbf5;
        src132 <= 12'h102;
        src133 <= 12'h77c;
        src134 <= 12'h503;
        src135 <= 12'h59a;
        src136 <= 12'h184;
        src137 <= 12'h338;
        src138 <= 12'h681;
        src139 <= 12'hd87;
        src140 <= 12'h5ea;
        src141 <= 12'he0a;
        src142 <= 12'hd77;
        src143 <= 12'h36d;
        src144 <= 12'hd3c;
        src145 <= 12'hd66;
        src146 <= 12'h854;
        src147 <= 12'hb5;
        src148 <= 12'hb3c;
        src149 <= 12'h62;
        src150 <= 12'hbfe;
        src151 <= 12'h187;
        src152 <= 12'h2;
        src153 <= 12'hc04;
        src154 <= 12'hb6c;
        src155 <= 12'hae6;
        src156 <= 12'ha96;
        src157 <= 12'h805;
        src158 <= 12'h227;
        src159 <= 12'h84;
        src160 <= 12'h124;
        src161 <= 12'h925;
        exp <= 20'h520bf;
        #1
        src0 <= 12'hde8;
        src1 <= 12'h530;
        src2 <= 12'h730;
        src3 <= 12'hb65;
        src4 <= 12'h8b1;
        src5 <= 12'h445;
        src6 <= 12'hc5b;
        src7 <= 12'hdd3;
        src8 <= 12'hdf4;
        src9 <= 12'h526;
        src10 <= 12'hdd5;
        src11 <= 12'hd75;
        src12 <= 12'hae4;
        src13 <= 12'hef1;
        src14 <= 12'hf9d;
        src15 <= 12'h466;
        src16 <= 12'h501;
        src17 <= 12'he80;
        src18 <= 12'h7b5;
        src19 <= 12'h874;
        src20 <= 12'h9fa;
        src21 <= 12'hd91;
        src22 <= 12'h9b;
        src23 <= 12'h592;
        src24 <= 12'hf20;
        src25 <= 12'h9d8;
        src26 <= 12'h44c;
        src27 <= 12'h9c0;
        src28 <= 12'h45f;
        src29 <= 12'h776;
        src30 <= 12'h29d;
        src31 <= 12'h8e6;
        src32 <= 12'h3ff;
        src33 <= 12'h117;
        src34 <= 12'h32c;
        src35 <= 12'h94a;
        src36 <= 12'h32e;
        src37 <= 12'hb9c;
        src38 <= 12'h2de;
        src39 <= 12'h376;
        src40 <= 12'h89d;
        src41 <= 12'h8bb;
        src42 <= 12'h351;
        src43 <= 12'hbb5;
        src44 <= 12'h57f;
        src45 <= 12'hc79;
        src46 <= 12'hdf0;
        src47 <= 12'hb3f;
        src48 <= 12'h487;
        src49 <= 12'h290;
        src50 <= 12'hc51;
        src51 <= 12'hb91;
        src52 <= 12'hee8;
        src53 <= 12'hf6f;
        src54 <= 12'h161;
        src55 <= 12'hc42;
        src56 <= 12'h184;
        src57 <= 12'h667;
        src58 <= 12'hb4c;
        src59 <= 12'h46a;
        src60 <= 12'hde0;
        src61 <= 12'ha96;
        src62 <= 12'h444;
        src63 <= 12'h790;
        src64 <= 12'h162;
        src65 <= 12'hd6;
        src66 <= 12'h6e7;
        src67 <= 12'h677;
        src68 <= 12'h10c;
        src69 <= 12'hed2;
        src70 <= 12'hd65;
        src71 <= 12'h669;
        src72 <= 12'h9e2;
        src73 <= 12'h46c;
        src74 <= 12'h7ce;
        src75 <= 12'h2de;
        src76 <= 12'h9e;
        src77 <= 12'h9e0;
        src78 <= 12'he74;
        src79 <= 12'hfd1;
        src80 <= 12'h76c;
        src81 <= 12'h7ed;
        src82 <= 12'h4e6;
        src83 <= 12'h1aa;
        src84 <= 12'he6e;
        src85 <= 12'hb25;
        src86 <= 12'h2f6;
        src87 <= 12'h882;
        src88 <= 12'h184;
        src89 <= 12'hf82;
        src90 <= 12'ha15;
        src91 <= 12'h7f6;
        src92 <= 12'hd11;
        src93 <= 12'h159;
        src94 <= 12'h961;
        src95 <= 12'had8;
        src96 <= 12'hf1a;
        src97 <= 12'hb7f;
        src98 <= 12'h5cb;
        src99 <= 12'hef3;
        src100 <= 12'h6e5;
        src101 <= 12'h168;
        src102 <= 12'h5da;
        src103 <= 12'h210;
        src104 <= 12'heb;
        src105 <= 12'h90c;
        src106 <= 12'hbd2;
        src107 <= 12'h54e;
        src108 <= 12'h36b;
        src109 <= 12'hb51;
        src110 <= 12'hf50;
        src111 <= 12'hf2;
        src112 <= 12'ha8f;
        src113 <= 12'ha8c;
        src114 <= 12'h905;
        src115 <= 12'h413;
        src116 <= 12'h948;
        src117 <= 12'ha70;
        src118 <= 12'he51;
        src119 <= 12'hc3d;
        src120 <= 12'h98d;
        src121 <= 12'h71c;
        src122 <= 12'h8ad;
        src123 <= 12'hac0;
        src124 <= 12'h6ee;
        src125 <= 12'hd2d;
        src126 <= 12'h363;
        src127 <= 12'hd43;
        src128 <= 12'hd50;
        src129 <= 12'hfe4;
        src130 <= 12'h74c;
        src131 <= 12'hed4;
        src132 <= 12'h7e5;
        src133 <= 12'h28d;
        src134 <= 12'h65;
        src135 <= 12'h467;
        src136 <= 12'hf;
        src137 <= 12'h4ba;
        src138 <= 12'h3af;
        src139 <= 12'h926;
        src140 <= 12'h82e;
        src141 <= 12'h826;
        src142 <= 12'ha14;
        src143 <= 12'ha12;
        src144 <= 12'h70b;
        src145 <= 12'h3fe;
        src146 <= 12'hb59;
        src147 <= 12'h603;
        src148 <= 12'he62;
        src149 <= 12'hc23;
        src150 <= 12'h3e1;
        src151 <= 12'hd6f;
        src152 <= 12'h2a6;
        src153 <= 12'h3cc;
        src154 <= 12'h122;
        src155 <= 12'hffc;
        src156 <= 12'h56f;
        src157 <= 12'h6b3;
        src158 <= 12'h621;
        src159 <= 12'h63;
        src160 <= 12'h571;
        src161 <= 12'h48;
        exp <= 20'h51b45;
        #1
        src0 <= 12'h10f;
        src1 <= 12'h3db;
        src2 <= 12'ha6f;
        src3 <= 12'he26;
        src4 <= 12'h454;
        src5 <= 12'h473;
        src6 <= 12'h34;
        src7 <= 12'h33e;
        src8 <= 12'he03;
        src9 <= 12'h1a5;
        src10 <= 12'h48c;
        src11 <= 12'hc28;
        src12 <= 12'h976;
        src13 <= 12'h296;
        src14 <= 12'h7a;
        src15 <= 12'h1d4;
        src16 <= 12'h590;
        src17 <= 12'hcdd;
        src18 <= 12'h4d6;
        src19 <= 12'hf2;
        src20 <= 12'h4b0;
        src21 <= 12'h8a7;
        src22 <= 12'h232;
        src23 <= 12'h45b;
        src24 <= 12'hb88;
        src25 <= 12'h1b1;
        src26 <= 12'had0;
        src27 <= 12'he4a;
        src28 <= 12'h698;
        src29 <= 12'hda2;
        src30 <= 12'hb7a;
        src31 <= 12'he8e;
        src32 <= 12'hfbb;
        src33 <= 12'h354;
        src34 <= 12'hda2;
        src35 <= 12'h3d0;
        src36 <= 12'h540;
        src37 <= 12'hb57;
        src38 <= 12'h7d2;
        src39 <= 12'h452;
        src40 <= 12'h9b1;
        src41 <= 12'hde3;
        src42 <= 12'hef2;
        src43 <= 12'h6ea;
        src44 <= 12'hec7;
        src45 <= 12'h93e;
        src46 <= 12'h150;
        src47 <= 12'hb77;
        src48 <= 12'h85;
        src49 <= 12'hc81;
        src50 <= 12'h8e;
        src51 <= 12'h448;
        src52 <= 12'h625;
        src53 <= 12'hf52;
        src54 <= 12'ha72;
        src55 <= 12'h186;
        src56 <= 12'h8f4;
        src57 <= 12'hf51;
        src58 <= 12'h3fe;
        src59 <= 12'h517;
        src60 <= 12'hd5d;
        src61 <= 12'h6dc;
        src62 <= 12'h901;
        src63 <= 12'h888;
        src64 <= 12'hb31;
        src65 <= 12'h5db;
        src66 <= 12'hf22;
        src67 <= 12'hb10;
        src68 <= 12'h315;
        src69 <= 12'h6b7;
        src70 <= 12'h52c;
        src71 <= 12'he52;
        src72 <= 12'h30c;
        src73 <= 12'h6e5;
        src74 <= 12'hc1b;
        src75 <= 12'ha89;
        src76 <= 12'ha7b;
        src77 <= 12'h257;
        src78 <= 12'h6be;
        src79 <= 12'ha53;
        src80 <= 12'hc87;
        src81 <= 12'h9cb;
        src82 <= 12'hd57;
        src83 <= 12'h413;
        src84 <= 12'h20c;
        src85 <= 12'hb0e;
        src86 <= 12'h581;
        src87 <= 12'h77d;
        src88 <= 12'h371;
        src89 <= 12'h82b;
        src90 <= 12'h12e;
        src91 <= 12'h488;
        src92 <= 12'hd4f;
        src93 <= 12'h227;
        src94 <= 12'h819;
        src95 <= 12'h6ef;
        src96 <= 12'h262;
        src97 <= 12'haf4;
        src98 <= 12'hc7e;
        src99 <= 12'h64d;
        src100 <= 12'h1f7;
        src101 <= 12'hd43;
        src102 <= 12'hf07;
        src103 <= 12'h103;
        src104 <= 12'h7;
        src105 <= 12'h6fc;
        src106 <= 12'hd89;
        src107 <= 12'h893;
        src108 <= 12'he1a;
        src109 <= 12'h57b;
        src110 <= 12'ha76;
        src111 <= 12'h703;
        src112 <= 12'h325;
        src113 <= 12'he9f;
        src114 <= 12'h822;
        src115 <= 12'hf8f;
        src116 <= 12'h6be;
        src117 <= 12'he43;
        src118 <= 12'h90b;
        src119 <= 12'h4a9;
        src120 <= 12'hbe5;
        src121 <= 12'ha78;
        src122 <= 12'haa7;
        src123 <= 12'h89a;
        src124 <= 12'h970;
        src125 <= 12'hf94;
        src126 <= 12'h40e;
        src127 <= 12'h80f;
        src128 <= 12'h50d;
        src129 <= 12'h4d2;
        src130 <= 12'h7ac;
        src131 <= 12'h30;
        src132 <= 12'h4c7;
        src133 <= 12'hd1b;
        src134 <= 12'hb1b;
        src135 <= 12'h140;
        src136 <= 12'hf3d;
        src137 <= 12'h53d;
        src138 <= 12'h3ab;
        src139 <= 12'h204;
        src140 <= 12'h6bf;
        src141 <= 12'hf69;
        src142 <= 12'h2d8;
        src143 <= 12'h62f;
        src144 <= 12'h6a;
        src145 <= 12'h352;
        src146 <= 12'h676;
        src147 <= 12'h1a2;
        src148 <= 12'h401;
        src149 <= 12'h2f1;
        src150 <= 12'ha96;
        src151 <= 12'h77b;
        src152 <= 12'h8af;
        src153 <= 12'hd75;
        src154 <= 12'hee4;
        src155 <= 12'hd52;
        src156 <= 12'h6e7;
        src157 <= 12'hc89;
        src158 <= 12'h275;
        src159 <= 12'hf20;
        src160 <= 12'h4c0;
        src161 <= 12'h389;
        exp <= 20'h4e9e9;
        #1
        src0 <= 12'hd26;
        src1 <= 12'hb9b;
        src2 <= 12'h4ef;
        src3 <= 12'hbe9;
        src4 <= 12'ha9d;
        src5 <= 12'h55d;
        src6 <= 12'h656;
        src7 <= 12'h639;
        src8 <= 12'hddc;
        src9 <= 12'h40;
        src10 <= 12'h9c2;
        src11 <= 12'h29c;
        src12 <= 12'hf86;
        src13 <= 12'hc7b;
        src14 <= 12'h415;
        src15 <= 12'h3b;
        src16 <= 12'h102;
        src17 <= 12'h52f;
        src18 <= 12'h1d;
        src19 <= 12'ha08;
        src20 <= 12'hddb;
        src21 <= 12'hc4f;
        src22 <= 12'h74;
        src23 <= 12'h158;
        src24 <= 12'h7ff;
        src25 <= 12'h862;
        src26 <= 12'h8a5;
        src27 <= 12'h160;
        src28 <= 12'h71d;
        src29 <= 12'h890;
        src30 <= 12'hc7;
        src31 <= 12'h8c8;
        src32 <= 12'h4a0;
        src33 <= 12'h376;
        src34 <= 12'h5c1;
        src35 <= 12'hf16;
        src36 <= 12'hc3d;
        src37 <= 12'h37e;
        src38 <= 12'h909;
        src39 <= 12'hf8;
        src40 <= 12'h3f8;
        src41 <= 12'h71b;
        src42 <= 12'h2de;
        src43 <= 12'h270;
        src44 <= 12'h543;
        src45 <= 12'h11d;
        src46 <= 12'h86f;
        src47 <= 12'hbc8;
        src48 <= 12'h7f8;
        src49 <= 12'h458;
        src50 <= 12'hc90;
        src51 <= 12'hf04;
        src52 <= 12'hd8d;
        src53 <= 12'he8a;
        src54 <= 12'hc7c;
        src55 <= 12'h6d5;
        src56 <= 12'h3c1;
        src57 <= 12'he0b;
        src58 <= 12'haeb;
        src59 <= 12'hf2d;
        src60 <= 12'h552;
        src61 <= 12'hadd;
        src62 <= 12'h3d;
        src63 <= 12'hdc1;
        src64 <= 12'h7d0;
        src65 <= 12'h364;
        src66 <= 12'h9f3;
        src67 <= 12'hd96;
        src68 <= 12'h7b8;
        src69 <= 12'h645;
        src70 <= 12'hb76;
        src71 <= 12'h8a7;
        src72 <= 12'hcb9;
        src73 <= 12'h445;
        src74 <= 12'hc26;
        src75 <= 12'h198;
        src76 <= 12'h7d7;
        src77 <= 12'hf11;
        src78 <= 12'hc24;
        src79 <= 12'h30;
        src80 <= 12'haab;
        src81 <= 12'h8c0;
        src82 <= 12'h926;
        src83 <= 12'h57a;
        src84 <= 12'h9f3;
        src85 <= 12'h65;
        src86 <= 12'h7ce;
        src87 <= 12'h5ba;
        src88 <= 12'hfdd;
        src89 <= 12'hb32;
        src90 <= 12'h77f;
        src91 <= 12'h8e4;
        src92 <= 12'h935;
        src93 <= 12'hb72;
        src94 <= 12'h99e;
        src95 <= 12'h40b;
        src96 <= 12'h203;
        src97 <= 12'h9de;
        src98 <= 12'h321;
        src99 <= 12'hb54;
        src100 <= 12'hf19;
        src101 <= 12'h8b2;
        src102 <= 12'h8b;
        src103 <= 12'h2be;
        src104 <= 12'h246;
        src105 <= 12'hb4;
        src106 <= 12'h549;
        src107 <= 12'hbe3;
        src108 <= 12'hd50;
        src109 <= 12'h9fa;
        src110 <= 12'h5df;
        src111 <= 12'ha0e;
        src112 <= 12'habb;
        src113 <= 12'hb32;
        src114 <= 12'hb8b;
        src115 <= 12'hb7a;
        src116 <= 12'hd68;
        src117 <= 12'ha9c;
        src118 <= 12'h151;
        src119 <= 12'hae6;
        src120 <= 12'h5c9;
        src121 <= 12'h852;
        src122 <= 12'h439;
        src123 <= 12'h824;
        src124 <= 12'h2e8;
        src125 <= 12'h744;
        src126 <= 12'ha3a;
        src127 <= 12'h38d;
        src128 <= 12'hf74;
        src129 <= 12'h19a;
        src130 <= 12'h86b;
        src131 <= 12'h134;
        src132 <= 12'h1c2;
        src133 <= 12'h7ee;
        src134 <= 12'he9e;
        src135 <= 12'h44;
        src136 <= 12'h36;
        src137 <= 12'h1d1;
        src138 <= 12'h815;
        src139 <= 12'had6;
        src140 <= 12'hf2e;
        src141 <= 12'h69d;
        src142 <= 12'he69;
        src143 <= 12'h8dd;
        src144 <= 12'h617;
        src145 <= 12'h572;
        src146 <= 12'hb8c;
        src147 <= 12'h6d;
        src148 <= 12'h918;
        src149 <= 12'h223;
        src150 <= 12'h6f1;
        src151 <= 12'hfa3;
        src152 <= 12'h5c8;
        src153 <= 12'h563;
        src154 <= 12'he1d;
        src155 <= 12'h25b;
        src156 <= 12'hef;
        src157 <= 12'h232;
        src158 <= 12'he08;
        src159 <= 12'h512;
        src160 <= 12'h27a;
        src161 <= 12'h55;
        exp <= 20'h4c9f4;
        #1
        src0 <= 12'ha1c;
        src1 <= 12'hdf7;
        src2 <= 12'hafa;
        src3 <= 12'h5f9;
        src4 <= 12'h851;
        src5 <= 12'h3b7;
        src6 <= 12'h7d5;
        src7 <= 12'h916;
        src8 <= 12'hcec;
        src9 <= 12'h4d9;
        src10 <= 12'hc49;
        src11 <= 12'h9d3;
        src12 <= 12'h124;
        src13 <= 12'h740;
        src14 <= 12'hb09;
        src15 <= 12'h794;
        src16 <= 12'h512;
        src17 <= 12'h806;
        src18 <= 12'h474;
        src19 <= 12'h668;
        src20 <= 12'heeb;
        src21 <= 12'h8ba;
        src22 <= 12'h3f9;
        src23 <= 12'h2cf;
        src24 <= 12'h3f8;
        src25 <= 12'h737;
        src26 <= 12'h745;
        src27 <= 12'he20;
        src28 <= 12'h9aa;
        src29 <= 12'h294;
        src30 <= 12'h7f4;
        src31 <= 12'h6bb;
        src32 <= 12'ha2e;
        src33 <= 12'hc65;
        src34 <= 12'h8fc;
        src35 <= 12'hf0a;
        src36 <= 12'h3ec;
        src37 <= 12'ha19;
        src38 <= 12'hf52;
        src39 <= 12'h7ad;
        src40 <= 12'hc9e;
        src41 <= 12'he97;
        src42 <= 12'h795;
        src43 <= 12'hca2;
        src44 <= 12'h40a;
        src45 <= 12'h5c4;
        src46 <= 12'h897;
        src47 <= 12'h572;
        src48 <= 12'hc08;
        src49 <= 12'h50;
        src50 <= 12'hcfb;
        src51 <= 12'hcf7;
        src52 <= 12'hdd0;
        src53 <= 12'ha01;
        src54 <= 12'ha8d;
        src55 <= 12'ha06;
        src56 <= 12'hbba;
        src57 <= 12'hf47;
        src58 <= 12'h9ea;
        src59 <= 12'hfd6;
        src60 <= 12'hecf;
        src61 <= 12'h8fc;
        src62 <= 12'hfc7;
        src63 <= 12'h393;
        src64 <= 12'h72e;
        src65 <= 12'h33d;
        src66 <= 12'hb1d;
        src67 <= 12'h84f;
        src68 <= 12'h24b;
        src69 <= 12'hc45;
        src70 <= 12'h79a;
        src71 <= 12'hd95;
        src72 <= 12'h673;
        src73 <= 12'h29d;
        src74 <= 12'h28d;
        src75 <= 12'hcb2;
        src76 <= 12'hfdc;
        src77 <= 12'h501;
        src78 <= 12'h7af;
        src79 <= 12'h79a;
        src80 <= 12'hbc9;
        src81 <= 12'h81e;
        src82 <= 12'hd8b;
        src83 <= 12'h5ac;
        src84 <= 12'h711;
        src85 <= 12'h5b1;
        src86 <= 12'h685;
        src87 <= 12'hf4d;
        src88 <= 12'h325;
        src89 <= 12'h48b;
        src90 <= 12'hedc;
        src91 <= 12'h190;
        src92 <= 12'h3ef;
        src93 <= 12'h602;
        src94 <= 12'h167;
        src95 <= 12'h910;
        src96 <= 12'h12;
        src97 <= 12'h79;
        src98 <= 12'hec3;
        src99 <= 12'h250;
        src100 <= 12'h12e;
        src101 <= 12'h300;
        src102 <= 12'hb0b;
        src103 <= 12'hf70;
        src104 <= 12'hda2;
        src105 <= 12'he1b;
        src106 <= 12'h8a1;
        src107 <= 12'h846;
        src108 <= 12'hb79;
        src109 <= 12'hff4;
        src110 <= 12'hd73;
        src111 <= 12'h43f;
        src112 <= 12'hf92;
        src113 <= 12'h18f;
        src114 <= 12'h550;
        src115 <= 12'h6d2;
        src116 <= 12'h1b7;
        src117 <= 12'hc37;
        src118 <= 12'h591;
        src119 <= 12'h90c;
        src120 <= 12'h8f;
        src121 <= 12'hb5d;
        src122 <= 12'hbed;
        src123 <= 12'h37e;
        src124 <= 12'h847;
        src125 <= 12'ha75;
        src126 <= 12'ha21;
        src127 <= 12'h2ae;
        src128 <= 12'h997;
        src129 <= 12'hd78;
        src130 <= 12'hd00;
        src131 <= 12'hb94;
        src132 <= 12'hfc5;
        src133 <= 12'h110;
        src134 <= 12'h4d;
        src135 <= 12'hc03;
        src136 <= 12'hfd3;
        src137 <= 12'h2d2;
        src138 <= 12'h999;
        src139 <= 12'h4a7;
        src140 <= 12'hab1;
        src141 <= 12'hd07;
        src142 <= 12'h87e;
        src143 <= 12'hf45;
        src144 <= 12'h123;
        src145 <= 12'hc15;
        src146 <= 12'hc9e;
        src147 <= 12'h2e;
        src148 <= 12'h233;
        src149 <= 12'h10d;
        src150 <= 12'had6;
        src151 <= 12'h93b;
        src152 <= 12'ha24;
        src153 <= 12'hb58;
        src154 <= 12'he5d;
        src155 <= 12'had6;
        src156 <= 12'h6ba;
        src157 <= 12'hd62;
        src158 <= 12'h21b;
        src159 <= 12'h454;
        src160 <= 12'h1e8;
        src161 <= 12'h724;
        exp <= 20'h55bef;
        #1
        src0 <= 12'h15f;
        src1 <= 12'h45d;
        src2 <= 12'he11;
        src3 <= 12'ha25;
        src4 <= 12'hefa;
        src5 <= 12'h1e5;
        src6 <= 12'h9f6;
        src7 <= 12'h7c2;
        src8 <= 12'hc89;
        src9 <= 12'h20b;
        src10 <= 12'hd0c;
        src11 <= 12'h7c;
        src12 <= 12'h8ad;
        src13 <= 12'he68;
        src14 <= 12'hbea;
        src15 <= 12'h3c0;
        src16 <= 12'h94a;
        src17 <= 12'h4d5;
        src18 <= 12'ha22;
        src19 <= 12'h530;
        src20 <= 12'h359;
        src21 <= 12'hc4a;
        src22 <= 12'hfb5;
        src23 <= 12'h21a;
        src24 <= 12'h394;
        src25 <= 12'h5e3;
        src26 <= 12'h92;
        src27 <= 12'hf84;
        src28 <= 12'hde3;
        src29 <= 12'h1c4;
        src30 <= 12'ha48;
        src31 <= 12'h35b;
        src32 <= 12'h1fa;
        src33 <= 12'he29;
        src34 <= 12'h79e;
        src35 <= 12'hf8b;
        src36 <= 12'h9c1;
        src37 <= 12'habb;
        src38 <= 12'hbbf;
        src39 <= 12'h2b5;
        src40 <= 12'ha88;
        src41 <= 12'h36d;
        src42 <= 12'h1fa;
        src43 <= 12'hd6;
        src44 <= 12'h8fa;
        src45 <= 12'h12a;
        src46 <= 12'hbd3;
        src47 <= 12'h2fe;
        src48 <= 12'hdc3;
        src49 <= 12'h6c2;
        src50 <= 12'h843;
        src51 <= 12'h3a0;
        src52 <= 12'he82;
        src53 <= 12'hf0f;
        src54 <= 12'h1b9;
        src55 <= 12'hd92;
        src56 <= 12'hfe9;
        src57 <= 12'h631;
        src58 <= 12'hdd9;
        src59 <= 12'h243;
        src60 <= 12'hdb5;
        src61 <= 12'h76;
        src62 <= 12'he29;
        src63 <= 12'h4cb;
        src64 <= 12'h6c0;
        src65 <= 12'h28a;
        src66 <= 12'hc33;
        src67 <= 12'hd4;
        src68 <= 12'h339;
        src69 <= 12'hcd9;
        src70 <= 12'hc61;
        src71 <= 12'hfa4;
        src72 <= 12'h4fa;
        src73 <= 12'h624;
        src74 <= 12'h4bb;
        src75 <= 12'h91;
        src76 <= 12'h530;
        src77 <= 12'h992;
        src78 <= 12'hbf9;
        src79 <= 12'hef1;
        src80 <= 12'h853;
        src81 <= 12'hbd9;
        src82 <= 12'ha57;
        src83 <= 12'h86;
        src84 <= 12'hf0a;
        src85 <= 12'h509;
        src86 <= 12'hb64;
        src87 <= 12'h629;
        src88 <= 12'h1d1;
        src89 <= 12'h77d;
        src90 <= 12'h22e;
        src91 <= 12'hb63;
        src92 <= 12'hc62;
        src93 <= 12'hce5;
        src94 <= 12'hdc0;
        src95 <= 12'hc81;
        src96 <= 12'hbf5;
        src97 <= 12'hc3e;
        src98 <= 12'h9e8;
        src99 <= 12'h4;
        src100 <= 12'h8c8;
        src101 <= 12'h3a6;
        src102 <= 12'hf90;
        src103 <= 12'h6a0;
        src104 <= 12'hd80;
        src105 <= 12'hcce;
        src106 <= 12'h44d;
        src107 <= 12'h78c;
        src108 <= 12'hf42;
        src109 <= 12'h1f3;
        src110 <= 12'hb45;
        src111 <= 12'he19;
        src112 <= 12'h550;
        src113 <= 12'hda5;
        src114 <= 12'h427;
        src115 <= 12'hb34;
        src116 <= 12'hfd5;
        src117 <= 12'hbc7;
        src118 <= 12'h51a;
        src119 <= 12'h6e2;
        src120 <= 12'h3e4;
        src121 <= 12'h3d2;
        src122 <= 12'h11d;
        src123 <= 12'h4d5;
        src124 <= 12'h9a0;
        src125 <= 12'hfc0;
        src126 <= 12'h105;
        src127 <= 12'h6e1;
        src128 <= 12'hffb;
        src129 <= 12'h9dc;
        src130 <= 12'hd4f;
        src131 <= 12'h1e3;
        src132 <= 12'h4d6;
        src133 <= 12'h13c;
        src134 <= 12'h50;
        src135 <= 12'h719;
        src136 <= 12'h2d3;
        src137 <= 12'h455;
        src138 <= 12'h974;
        src139 <= 12'h25e;
        src140 <= 12'h9c9;
        src141 <= 12'h20e;
        src142 <= 12'ha70;
        src143 <= 12'h4f;
        src144 <= 12'hfb8;
        src145 <= 12'he6c;
        src146 <= 12'h8ac;
        src147 <= 12'h198;
        src148 <= 12'h1a7;
        src149 <= 12'h864;
        src150 <= 12'h137;
        src151 <= 12'hd9;
        src152 <= 12'h3b3;
        src153 <= 12'h5a4;
        src154 <= 12'h54e;
        src155 <= 12'h988;
        src156 <= 12'h554;
        src157 <= 12'h276;
        src158 <= 12'h5a4;
        src159 <= 12'h49;
        src160 <= 12'h2ff;
        src161 <= 12'hd13;
        exp <= 20'h4e615;
        #1
        src0 <= 12'hc05;
        src1 <= 12'h7c5;
        src2 <= 12'he6f;
        src3 <= 12'hb5;
        src4 <= 12'h584;
        src5 <= 12'h4b2;
        src6 <= 12'haec;
        src7 <= 12'h801;
        src8 <= 12'he43;
        src9 <= 12'ha83;
        src10 <= 12'haae;
        src11 <= 12'h308;
        src12 <= 12'hcb1;
        src13 <= 12'h28b;
        src14 <= 12'h1ee;
        src15 <= 12'h943;
        src16 <= 12'h70c;
        src17 <= 12'hd7e;
        src18 <= 12'hbd6;
        src19 <= 12'hca8;
        src20 <= 12'h507;
        src21 <= 12'he40;
        src22 <= 12'haf2;
        src23 <= 12'h54a;
        src24 <= 12'h78a;
        src25 <= 12'h51e;
        src26 <= 12'h48b;
        src27 <= 12'hd07;
        src28 <= 12'h455;
        src29 <= 12'h5e2;
        src30 <= 12'hc7;
        src31 <= 12'h8c6;
        src32 <= 12'h2c8;
        src33 <= 12'h9c1;
        src34 <= 12'hc15;
        src35 <= 12'h6db;
        src36 <= 12'hd9e;
        src37 <= 12'hcc0;
        src38 <= 12'h7ee;
        src39 <= 12'hc53;
        src40 <= 12'h7d2;
        src41 <= 12'h396;
        src42 <= 12'h791;
        src43 <= 12'h42b;
        src44 <= 12'ha45;
        src45 <= 12'h883;
        src46 <= 12'h87e;
        src47 <= 12'h8be;
        src48 <= 12'hce0;
        src49 <= 12'h39b;
        src50 <= 12'hdac;
        src51 <= 12'h582;
        src52 <= 12'hdb;
        src53 <= 12'hf57;
        src54 <= 12'hfa3;
        src55 <= 12'h370;
        src56 <= 12'h329;
        src57 <= 12'h385;
        src58 <= 12'hc13;
        src59 <= 12'h93f;
        src60 <= 12'hb57;
        src61 <= 12'h4e0;
        src62 <= 12'h576;
        src63 <= 12'hbb5;
        src64 <= 12'h680;
        src65 <= 12'h300;
        src66 <= 12'hf62;
        src67 <= 12'h400;
        src68 <= 12'hb97;
        src69 <= 12'h9b9;
        src70 <= 12'he83;
        src71 <= 12'h21f;
        src72 <= 12'hb02;
        src73 <= 12'ha35;
        src74 <= 12'h586;
        src75 <= 12'h2cd;
        src76 <= 12'h91d;
        src77 <= 12'hfae;
        src78 <= 12'hfe;
        src79 <= 12'h46c;
        src80 <= 12'he3b;
        src81 <= 12'h8ac;
        src82 <= 12'h557;
        src83 <= 12'hd0b;
        src84 <= 12'hf8e;
        src85 <= 12'h226;
        src86 <= 12'h7b0;
        src87 <= 12'h886;
        src88 <= 12'h214;
        src89 <= 12'h27;
        src90 <= 12'h7ee;
        src91 <= 12'hce0;
        src92 <= 12'he5;
        src93 <= 12'hcf1;
        src94 <= 12'h263;
        src95 <= 12'h233;
        src96 <= 12'h39d;
        src97 <= 12'hee3;
        src98 <= 12'hbe3;
        src99 <= 12'h999;
        src100 <= 12'he0e;
        src101 <= 12'h1f1;
        src102 <= 12'hb2a;
        src103 <= 12'h7f5;
        src104 <= 12'h4da;
        src105 <= 12'h2a8;
        src106 <= 12'heed;
        src107 <= 12'he35;
        src108 <= 12'h560;
        src109 <= 12'h7de;
        src110 <= 12'h6d7;
        src111 <= 12'hd4e;
        src112 <= 12'hc9e;
        src113 <= 12'h832;
        src114 <= 12'h6fc;
        src115 <= 12'h836;
        src116 <= 12'h333;
        src117 <= 12'h8a6;
        src118 <= 12'hd9f;
        src119 <= 12'h937;
        src120 <= 12'h57c;
        src121 <= 12'hed8;
        src122 <= 12'h610;
        src123 <= 12'h276;
        src124 <= 12'he74;
        src125 <= 12'h289;
        src126 <= 12'h669;
        src127 <= 12'he22;
        src128 <= 12'had9;
        src129 <= 12'h6f1;
        src130 <= 12'hba;
        src131 <= 12'h141;
        src132 <= 12'h522;
        src133 <= 12'hefc;
        src134 <= 12'h1bb;
        src135 <= 12'hcb0;
        src136 <= 12'h282;
        src137 <= 12'hd73;
        src138 <= 12'h9c0;
        src139 <= 12'hd97;
        src140 <= 12'hba1;
        src141 <= 12'ha45;
        src142 <= 12'h81c;
        src143 <= 12'hf12;
        src144 <= 12'hff9;
        src145 <= 12'hddd;
        src146 <= 12'hb77;
        src147 <= 12'h99a;
        src148 <= 12'h515;
        src149 <= 12'h28c;
        src150 <= 12'hbd0;
        src151 <= 12'h4c8;
        src152 <= 12'hb01;
        src153 <= 12'h983;
        src154 <= 12'h645;
        src155 <= 12'h28d;
        src156 <= 12'hdb5;
        src157 <= 12'h975;
        src158 <= 12'h709;
        src159 <= 12'h78f;
        src160 <= 12'h99;
        src161 <= 12'h671;
        exp <= 20'h53e72;
        #1
        src0 <= 12'h84c;
        src1 <= 12'h1d9;
        src2 <= 12'h317;
        src3 <= 12'hd34;
        src4 <= 12'hde7;
        src5 <= 12'hdbb;
        src6 <= 12'h317;
        src7 <= 12'h8d2;
        src8 <= 12'hb00;
        src9 <= 12'hefe;
        src10 <= 12'hd62;
        src11 <= 12'h553;
        src12 <= 12'hec4;
        src13 <= 12'h961;
        src14 <= 12'hf48;
        src15 <= 12'h41e;
        src16 <= 12'hd8b;
        src17 <= 12'hd5;
        src18 <= 12'h1c6;
        src19 <= 12'h448;
        src20 <= 12'h72f;
        src21 <= 12'h4ce;
        src22 <= 12'h6de;
        src23 <= 12'hb13;
        src24 <= 12'h20;
        src25 <= 12'h95c;
        src26 <= 12'h88b;
        src27 <= 12'h93a;
        src28 <= 12'h835;
        src29 <= 12'hba0;
        src30 <= 12'h524;
        src31 <= 12'h42d;
        src32 <= 12'hafb;
        src33 <= 12'h87b;
        src34 <= 12'h49d;
        src35 <= 12'hce5;
        src36 <= 12'hb59;
        src37 <= 12'h425;
        src38 <= 12'h82e;
        src39 <= 12'h7a6;
        src40 <= 12'hb5f;
        src41 <= 12'h649;
        src42 <= 12'haac;
        src43 <= 12'hc7;
        src44 <= 12'hacb;
        src45 <= 12'he03;
        src46 <= 12'h257;
        src47 <= 12'hd5b;
        src48 <= 12'h2e3;
        src49 <= 12'hfda;
        src50 <= 12'hfc2;
        src51 <= 12'he67;
        src52 <= 12'h91d;
        src53 <= 12'hf3f;
        src54 <= 12'h16e;
        src55 <= 12'hc87;
        src56 <= 12'h433;
        src57 <= 12'h812;
        src58 <= 12'h6f;
        src59 <= 12'hfa6;
        src60 <= 12'hc4e;
        src61 <= 12'hf0c;
        src62 <= 12'hfd5;
        src63 <= 12'h346;
        src64 <= 12'hbf0;
        src65 <= 12'h229;
        src66 <= 12'h87c;
        src67 <= 12'h3c6;
        src68 <= 12'h9fc;
        src69 <= 12'hbab;
        src70 <= 12'hd89;
        src71 <= 12'h9dd;
        src72 <= 12'h5ec;
        src73 <= 12'h4f6;
        src74 <= 12'h881;
        src75 <= 12'hab0;
        src76 <= 12'h92e;
        src77 <= 12'h358;
        src78 <= 12'h568;
        src79 <= 12'hf73;
        src80 <= 12'h82b;
        src81 <= 12'h5d7;
        src82 <= 12'hbc;
        src83 <= 12'h603;
        src84 <= 12'hd07;
        src85 <= 12'hadb;
        src86 <= 12'hede;
        src87 <= 12'hb4;
        src88 <= 12'he55;
        src89 <= 12'hcc7;
        src90 <= 12'h295;
        src91 <= 12'h855;
        src92 <= 12'he15;
        src93 <= 12'h589;
        src94 <= 12'h974;
        src95 <= 12'h4c5;
        src96 <= 12'h438;
        src97 <= 12'h26d;
        src98 <= 12'h71c;
        src99 <= 12'h489;
        src100 <= 12'h554;
        src101 <= 12'h7da;
        src102 <= 12'h7f;
        src103 <= 12'hf2e;
        src104 <= 12'h9d1;
        src105 <= 12'ha74;
        src106 <= 12'h5d9;
        src107 <= 12'ha46;
        src108 <= 12'hc8d;
        src109 <= 12'hfa3;
        src110 <= 12'h5e2;
        src111 <= 12'h737;
        src112 <= 12'h630;
        src113 <= 12'h824;
        src114 <= 12'h409;
        src115 <= 12'hcf0;
        src116 <= 12'hc45;
        src117 <= 12'hd2;
        src118 <= 12'h8;
        src119 <= 12'hf4f;
        src120 <= 12'h86f;
        src121 <= 12'hfb3;
        src122 <= 12'hfa9;
        src123 <= 12'h6dc;
        src124 <= 12'hae1;
        src125 <= 12'hef0;
        src126 <= 12'hb05;
        src127 <= 12'h45b;
        src128 <= 12'h174;
        src129 <= 12'h4a5;
        src130 <= 12'h47f;
        src131 <= 12'hcfd;
        src132 <= 12'h1e8;
        src133 <= 12'h486;
        src134 <= 12'h69b;
        src135 <= 12'h3d;
        src136 <= 12'hedc;
        src137 <= 12'h731;
        src138 <= 12'h999;
        src139 <= 12'h770;
        src140 <= 12'h829;
        src141 <= 12'heaf;
        src142 <= 12'h7eb;
        src143 <= 12'hb28;
        src144 <= 12'hc31;
        src145 <= 12'h7cb;
        src146 <= 12'hedd;
        src147 <= 12'h3f6;
        src148 <= 12'hbb4;
        src149 <= 12'hcc3;
        src150 <= 12'h65d;
        src151 <= 12'h7fc;
        src152 <= 12'hb50;
        src153 <= 12'hafc;
        src154 <= 12'he99;
        src155 <= 12'h86f;
        src156 <= 12'h692;
        src157 <= 12'h36a;
        src158 <= 12'hcef;
        src159 <= 12'h5a4;
        src160 <= 12'h5dd;
        src161 <= 12'h363;
        exp <= 20'h562d8;
        #1
        src0 <= 12'h810;
        src1 <= 12'h762;
        src2 <= 12'h2c9;
        src3 <= 12'h80c;
        src4 <= 12'h9eb;
        src5 <= 12'h6b8;
        src6 <= 12'h468;
        src7 <= 12'h558;
        src8 <= 12'h996;
        src9 <= 12'hb1c;
        src10 <= 12'h9a3;
        src11 <= 12'hfec;
        src12 <= 12'h23c;
        src13 <= 12'ha84;
        src14 <= 12'he4a;
        src15 <= 12'hba5;
        src16 <= 12'he6a;
        src17 <= 12'hd3c;
        src18 <= 12'ha7a;
        src19 <= 12'h206;
        src20 <= 12'h170;
        src21 <= 12'hb6f;
        src22 <= 12'h73e;
        src23 <= 12'haf6;
        src24 <= 12'hc83;
        src25 <= 12'hc59;
        src26 <= 12'h63f;
        src27 <= 12'h47f;
        src28 <= 12'h255;
        src29 <= 12'heaa;
        src30 <= 12'h603;
        src31 <= 12'h8f2;
        src32 <= 12'h1e5;
        src33 <= 12'h820;
        src34 <= 12'h7a4;
        src35 <= 12'h9be;
        src36 <= 12'h88b;
        src37 <= 12'h899;
        src38 <= 12'h83f;
        src39 <= 12'h22c;
        src40 <= 12'hcce;
        src41 <= 12'hc5e;
        src42 <= 12'hb6a;
        src43 <= 12'hc22;
        src44 <= 12'hc0d;
        src45 <= 12'h45f;
        src46 <= 12'h450;
        src47 <= 12'h20a;
        src48 <= 12'h6e6;
        src49 <= 12'h7be;
        src50 <= 12'hcde;
        src51 <= 12'h30c;
        src52 <= 12'h962;
        src53 <= 12'hb9a;
        src54 <= 12'h65a;
        src55 <= 12'hb9b;
        src56 <= 12'hee5;
        src57 <= 12'h989;
        src58 <= 12'hd59;
        src59 <= 12'hf2a;
        src60 <= 12'haa3;
        src61 <= 12'h105;
        src62 <= 12'hc29;
        src63 <= 12'h2ab;
        src64 <= 12'hd81;
        src65 <= 12'h209;
        src66 <= 12'h308;
        src67 <= 12'h6cf;
        src68 <= 12'h14b;
        src69 <= 12'hddd;
        src70 <= 12'hf4b;
        src71 <= 12'h104;
        src72 <= 12'h8cf;
        src73 <= 12'hc0e;
        src74 <= 12'h54a;
        src75 <= 12'hf2e;
        src76 <= 12'h345;
        src77 <= 12'hf99;
        src78 <= 12'h3b8;
        src79 <= 12'h963;
        src80 <= 12'he5c;
        src81 <= 12'h439;
        src82 <= 12'h995;
        src83 <= 12'hc42;
        src84 <= 12'h314;
        src85 <= 12'hfd8;
        src86 <= 12'h490;
        src87 <= 12'hb37;
        src88 <= 12'h3f4;
        src89 <= 12'hc0d;
        src90 <= 12'h1bd;
        src91 <= 12'heac;
        src92 <= 12'h419;
        src93 <= 12'hdad;
        src94 <= 12'h20a;
        src95 <= 12'h54b;
        src96 <= 12'h40;
        src97 <= 12'h32c;
        src98 <= 12'ha3b;
        src99 <= 12'h258;
        src100 <= 12'h922;
        src101 <= 12'hfb9;
        src102 <= 12'hd76;
        src103 <= 12'h35f;
        src104 <= 12'h856;
        src105 <= 12'h8c4;
        src106 <= 12'hc8c;
        src107 <= 12'h5f5;
        src108 <= 12'h8f9;
        src109 <= 12'h9c5;
        src110 <= 12'h1fd;
        src111 <= 12'h159;
        src112 <= 12'h334;
        src113 <= 12'h76c;
        src114 <= 12'h898;
        src115 <= 12'h1a8;
        src116 <= 12'ha00;
        src117 <= 12'h93;
        src118 <= 12'hcf0;
        src119 <= 12'h2fc;
        src120 <= 12'heab;
        src121 <= 12'hcbf;
        src122 <= 12'hf2e;
        src123 <= 12'h1c9;
        src124 <= 12'hb77;
        src125 <= 12'h9af;
        src126 <= 12'h620;
        src127 <= 12'h623;
        src128 <= 12'hc4a;
        src129 <= 12'h31c;
        src130 <= 12'h84b;
        src131 <= 12'h8a1;
        src132 <= 12'h772;
        src133 <= 12'h111;
        src134 <= 12'h2f5;
        src135 <= 12'h8d1;
        src136 <= 12'h82d;
        src137 <= 12'h1e4;
        src138 <= 12'h1f3;
        src139 <= 12'h789;
        src140 <= 12'hec7;
        src141 <= 12'h282;
        src142 <= 12'h738;
        src143 <= 12'h7d9;
        src144 <= 12'h6eb;
        src145 <= 12'hd56;
        src146 <= 12'h992;
        src147 <= 12'h2c3;
        src148 <= 12'h391;
        src149 <= 12'h713;
        src150 <= 12'h450;
        src151 <= 12'ha07;
        src152 <= 12'hb7f;
        src153 <= 12'h5a;
        src154 <= 12'h773;
        src155 <= 12'h6c4;
        src156 <= 12'hc0e;
        src157 <= 12'h1d5;
        src158 <= 12'h56c;
        src159 <= 12'hd79;
        src160 <= 12'h8eb;
        src161 <= 12'h6bd;
        exp <= 20'h50ba5;
        #1
        src0 <= 12'hcc9;
        src1 <= 12'hccd;
        src2 <= 12'h9a2;
        src3 <= 12'h317;
        src4 <= 12'h64b;
        src5 <= 12'h5a0;
        src6 <= 12'ha8c;
        src7 <= 12'h7ea;
        src8 <= 12'h99b;
        src9 <= 12'h35e;
        src10 <= 12'hcf3;
        src11 <= 12'hf39;
        src12 <= 12'hd92;
        src13 <= 12'h8f7;
        src14 <= 12'he6a;
        src15 <= 12'h3a4;
        src16 <= 12'ha58;
        src17 <= 12'hc9c;
        src18 <= 12'hcc3;
        src19 <= 12'hc17;
        src20 <= 12'hdf5;
        src21 <= 12'h242;
        src22 <= 12'h2f6;
        src23 <= 12'h2d7;
        src24 <= 12'ha76;
        src25 <= 12'h387;
        src26 <= 12'h7b7;
        src27 <= 12'h9cb;
        src28 <= 12'h924;
        src29 <= 12'hcf0;
        src30 <= 12'h22e;
        src31 <= 12'h9ac;
        src32 <= 12'hef9;
        src33 <= 12'hd7;
        src34 <= 12'h96d;
        src35 <= 12'had;
        src36 <= 12'he;
        src37 <= 12'hea8;
        src38 <= 12'had0;
        src39 <= 12'h235;
        src40 <= 12'hed7;
        src41 <= 12'hb92;
        src42 <= 12'h575;
        src43 <= 12'hf47;
        src44 <= 12'h9e4;
        src45 <= 12'hf15;
        src46 <= 12'h45e;
        src47 <= 12'h8e8;
        src48 <= 12'h668;
        src49 <= 12'h7b6;
        src50 <= 12'h620;
        src51 <= 12'hdb0;
        src52 <= 12'ha33;
        src53 <= 12'h6d;
        src54 <= 12'hd0c;
        src55 <= 12'hcc;
        src56 <= 12'h80b;
        src57 <= 12'hc14;
        src58 <= 12'h3c6;
        src59 <= 12'h4a6;
        src60 <= 12'h82a;
        src61 <= 12'ha70;
        src62 <= 12'h17f;
        src63 <= 12'h5ce;
        src64 <= 12'hc2b;
        src65 <= 12'h8a7;
        src66 <= 12'h440;
        src67 <= 12'h1af;
        src68 <= 12'h199;
        src69 <= 12'h77a;
        src70 <= 12'h637;
        src71 <= 12'hd7a;
        src72 <= 12'hf27;
        src73 <= 12'hc14;
        src74 <= 12'h55;
        src75 <= 12'hdfd;
        src76 <= 12'hb20;
        src77 <= 12'hf2e;
        src78 <= 12'h844;
        src79 <= 12'h88e;
        src80 <= 12'hb0;
        src81 <= 12'h6d2;
        src82 <= 12'hc4;
        src83 <= 12'h345;
        src84 <= 12'h729;
        src85 <= 12'h5e4;
        src86 <= 12'hc4c;
        src87 <= 12'h232;
        src88 <= 12'h2e7;
        src89 <= 12'h819;
        src90 <= 12'h25a;
        src91 <= 12'he26;
        src92 <= 12'h1a4;
        src93 <= 12'hfe2;
        src94 <= 12'hb67;
        src95 <= 12'hdd6;
        src96 <= 12'h76d;
        src97 <= 12'h843;
        src98 <= 12'h104;
        src99 <= 12'hfde;
        src100 <= 12'hfd4;
        src101 <= 12'ha51;
        src102 <= 12'h677;
        src103 <= 12'hc8c;
        src104 <= 12'h942;
        src105 <= 12'hade;
        src106 <= 12'h233;
        src107 <= 12'h8a2;
        src108 <= 12'hd5a;
        src109 <= 12'h57d;
        src110 <= 12'hf90;
        src111 <= 12'hcc3;
        src112 <= 12'he94;
        src113 <= 12'h60c;
        src114 <= 12'h280;
        src115 <= 12'h96a;
        src116 <= 12'he16;
        src117 <= 12'ha9a;
        src118 <= 12'h252;
        src119 <= 12'ha1d;
        src120 <= 12'h517;
        src121 <= 12'h19f;
        src122 <= 12'h630;
        src123 <= 12'hc00;
        src124 <= 12'h879;
        src125 <= 12'hc42;
        src126 <= 12'h581;
        src127 <= 12'h950;
        src128 <= 12'h812;
        src129 <= 12'h131;
        src130 <= 12'h5b2;
        src131 <= 12'h8da;
        src132 <= 12'hd4c;
        src133 <= 12'h7e1;
        src134 <= 12'hdee;
        src135 <= 12'h73b;
        src136 <= 12'h64d;
        src137 <= 12'hebf;
        src138 <= 12'h8b1;
        src139 <= 12'h6eb;
        src140 <= 12'h601;
        src141 <= 12'h5e5;
        src142 <= 12'h532;
        src143 <= 12'hccc;
        src144 <= 12'h402;
        src145 <= 12'h374;
        src146 <= 12'h283;
        src147 <= 12'h71c;
        src148 <= 12'h817;
        src149 <= 12'h5a7;
        src150 <= 12'h9da;
        src151 <= 12'h844;
        src152 <= 12'hda4;
        src153 <= 12'h91f;
        src154 <= 12'hc5c;
        src155 <= 12'h88a;
        src156 <= 12'h6df;
        src157 <= 12'hc90;
        src158 <= 12'ha60;
        src159 <= 12'hb13;
        src160 <= 12'h74d;
        src161 <= 12'ha29;
        exp <= 20'h54cae;
        #1
        src0 <= 12'h5f1;
        src1 <= 12'h7a0;
        src2 <= 12'he23;
        src3 <= 12'h20f;
        src4 <= 12'he0e;
        src5 <= 12'hcae;
        src6 <= 12'h675;
        src7 <= 12'h4e;
        src8 <= 12'ha7f;
        src9 <= 12'h5aa;
        src10 <= 12'hace;
        src11 <= 12'h12b;
        src12 <= 12'hcfa;
        src13 <= 12'h819;
        src14 <= 12'hde1;
        src15 <= 12'h4c;
        src16 <= 12'hc0f;
        src17 <= 12'h12e;
        src18 <= 12'h467;
        src19 <= 12'h89;
        src20 <= 12'h9c2;
        src21 <= 12'h3e;
        src22 <= 12'hc85;
        src23 <= 12'h8c1;
        src24 <= 12'hbb7;
        src25 <= 12'he78;
        src26 <= 12'h530;
        src27 <= 12'h77;
        src28 <= 12'hd0f;
        src29 <= 12'h2e;
        src30 <= 12'h704;
        src31 <= 12'h126;
        src32 <= 12'h8a7;
        src33 <= 12'h47d;
        src34 <= 12'h374;
        src35 <= 12'h854;
        src36 <= 12'h8a3;
        src37 <= 12'h181;
        src38 <= 12'h98;
        src39 <= 12'h6d8;
        src40 <= 12'h9c7;
        src41 <= 12'hc95;
        src42 <= 12'hc9d;
        src43 <= 12'ha8e;
        src44 <= 12'hc19;
        src45 <= 12'h992;
        src46 <= 12'hf1a;
        src47 <= 12'h1fc;
        src48 <= 12'h890;
        src49 <= 12'h50d;
        src50 <= 12'h438;
        src51 <= 12'h9c4;
        src52 <= 12'h568;
        src53 <= 12'haff;
        src54 <= 12'h86;
        src55 <= 12'h140;
        src56 <= 12'had4;
        src57 <= 12'h9df;
        src58 <= 12'h1ec;
        src59 <= 12'h786;
        src60 <= 12'h315;
        src61 <= 12'hc03;
        src62 <= 12'h404;
        src63 <= 12'h4d5;
        src64 <= 12'h138;
        src65 <= 12'h342;
        src66 <= 12'h5f;
        src67 <= 12'h6a0;
        src68 <= 12'ha53;
        src69 <= 12'hf07;
        src70 <= 12'h481;
        src71 <= 12'h971;
        src72 <= 12'h883;
        src73 <= 12'h1f9;
        src74 <= 12'h77c;
        src75 <= 12'h903;
        src76 <= 12'h244;
        src77 <= 12'h931;
        src78 <= 12'hf9b;
        src79 <= 12'h429;
        src80 <= 12'hb18;
        src81 <= 12'h9a3;
        src82 <= 12'hb68;
        src83 <= 12'he80;
        src84 <= 12'h16;
        src85 <= 12'h89d;
        src86 <= 12'ha06;
        src87 <= 12'h45b;
        src88 <= 12'h21f;
        src89 <= 12'hae9;
        src90 <= 12'hfd1;
        src91 <= 12'h40a;
        src92 <= 12'h624;
        src93 <= 12'hd7d;
        src94 <= 12'hd07;
        src95 <= 12'h82;
        src96 <= 12'hac4;
        src97 <= 12'h5af;
        src98 <= 12'hda1;
        src99 <= 12'hd85;
        src100 <= 12'hf46;
        src101 <= 12'ha6b;
        src102 <= 12'h266;
        src103 <= 12'h3e1;
        src104 <= 12'h31a;
        src105 <= 12'h2a7;
        src106 <= 12'h86;
        src107 <= 12'hc5f;
        src108 <= 12'h784;
        src109 <= 12'h3f2;
        src110 <= 12'h462;
        src111 <= 12'h245;
        src112 <= 12'h1ea;
        src113 <= 12'h964;
        src114 <= 12'hefe;
        src115 <= 12'h29c;
        src116 <= 12'h833;
        src117 <= 12'h499;
        src118 <= 12'h83;
        src119 <= 12'hb76;
        src120 <= 12'h792;
        src121 <= 12'hc2e;
        src122 <= 12'hd5;
        src123 <= 12'h81d;
        src124 <= 12'hb12;
        src125 <= 12'h292;
        src126 <= 12'h63f;
        src127 <= 12'hb0f;
        src128 <= 12'hc28;
        src129 <= 12'h8f9;
        src130 <= 12'h8ad;
        src131 <= 12'h34d;
        src132 <= 12'hc8b;
        src133 <= 12'h527;
        src134 <= 12'h778;
        src135 <= 12'h60e;
        src136 <= 12'he35;
        src137 <= 12'hd4;
        src138 <= 12'h509;
        src139 <= 12'h3b;
        src140 <= 12'hddd;
        src141 <= 12'h2b3;
        src142 <= 12'h864;
        src143 <= 12'hdb8;
        src144 <= 12'h7f7;
        src145 <= 12'h1e4;
        src146 <= 12'h979;
        src147 <= 12'h6a9;
        src148 <= 12'hc45;
        src149 <= 12'hd55;
        src150 <= 12'h56c;
        src151 <= 12'h1bd;
        src152 <= 12'h2b8;
        src153 <= 12'hacd;
        src154 <= 12'hd05;
        src155 <= 12'hc35;
        src156 <= 12'ha13;
        src157 <= 12'h529;
        src158 <= 12'ha7c;
        src159 <= 12'h166;
        src160 <= 12'hcb9;
        src161 <= 12'h843;
        exp <= 20'h4ab3f;
        #1
        src0 <= 12'h214;
        src1 <= 12'h676;
        src2 <= 12'he89;
        src3 <= 12'h42b;
        src4 <= 12'hd83;
        src5 <= 12'h3df;
        src6 <= 12'hcdc;
        src7 <= 12'hca3;
        src8 <= 12'hc56;
        src9 <= 12'h2fa;
        src10 <= 12'h491;
        src11 <= 12'he2;
        src12 <= 12'ha95;
        src13 <= 12'he2c;
        src14 <= 12'hc7b;
        src15 <= 12'h44d;
        src16 <= 12'ha10;
        src17 <= 12'hef0;
        src18 <= 12'hdbc;
        src19 <= 12'h6be;
        src20 <= 12'he8e;
        src21 <= 12'h78;
        src22 <= 12'h827;
        src23 <= 12'hca7;
        src24 <= 12'haf1;
        src25 <= 12'h91a;
        src26 <= 12'h3e8;
        src27 <= 12'h9b3;
        src28 <= 12'h90b;
        src29 <= 12'hc2d;
        src30 <= 12'h398;
        src31 <= 12'h6d5;
        src32 <= 12'h847;
        src33 <= 12'h45b;
        src34 <= 12'hc71;
        src35 <= 12'hcf4;
        src36 <= 12'hbfa;
        src37 <= 12'h5d0;
        src38 <= 12'h1fb;
        src39 <= 12'h8ec;
        src40 <= 12'hc4a;
        src41 <= 12'h749;
        src42 <= 12'hcc6;
        src43 <= 12'h6a;
        src44 <= 12'h25b;
        src45 <= 12'hcfb;
        src46 <= 12'h8f4;
        src47 <= 12'hcf5;
        src48 <= 12'h11;
        src49 <= 12'h736;
        src50 <= 12'h4d0;
        src51 <= 12'h4c9;
        src52 <= 12'h57;
        src53 <= 12'h43d;
        src54 <= 12'h3b2;
        src55 <= 12'h548;
        src56 <= 12'h7e2;
        src57 <= 12'hae9;
        src58 <= 12'h370;
        src59 <= 12'h82f;
        src60 <= 12'hdf6;
        src61 <= 12'hd93;
        src62 <= 12'h9d7;
        src63 <= 12'hb23;
        src64 <= 12'hb1a;
        src65 <= 12'h7cc;
        src66 <= 12'h11e;
        src67 <= 12'ha5b;
        src68 <= 12'h9c5;
        src69 <= 12'hf99;
        src70 <= 12'h2ae;
        src71 <= 12'h933;
        src72 <= 12'hf76;
        src73 <= 12'h42a;
        src74 <= 12'h6e3;
        src75 <= 12'h79;
        src76 <= 12'hc9d;
        src77 <= 12'h518;
        src78 <= 12'h4c6;
        src79 <= 12'h76f;
        src80 <= 12'h20b;
        src81 <= 12'ha43;
        src82 <= 12'h6c0;
        src83 <= 12'h717;
        src84 <= 12'h896;
        src85 <= 12'hb83;
        src86 <= 12'h5e4;
        src87 <= 12'ha36;
        src88 <= 12'h6f9;
        src89 <= 12'h697;
        src90 <= 12'h371;
        src91 <= 12'h1eb;
        src92 <= 12'hdb4;
        src93 <= 12'hca0;
        src94 <= 12'h6e9;
        src95 <= 12'h11;
        src96 <= 12'h7ef;
        src97 <= 12'hbcd;
        src98 <= 12'h238;
        src99 <= 12'h1a;
        src100 <= 12'h332;
        src101 <= 12'he2c;
        src102 <= 12'h27b;
        src103 <= 12'ha51;
        src104 <= 12'h272;
        src105 <= 12'h965;
        src106 <= 12'h1cb;
        src107 <= 12'h6c4;
        src108 <= 12'h901;
        src109 <= 12'hee6;
        src110 <= 12'h302;
        src111 <= 12'hda;
        src112 <= 12'hb0b;
        src113 <= 12'h865;
        src114 <= 12'h24d;
        src115 <= 12'hef4;
        src116 <= 12'h451;
        src117 <= 12'h561;
        src118 <= 12'h3ad;
        src119 <= 12'h94b;
        src120 <= 12'hfb8;
        src121 <= 12'h7c1;
        src122 <= 12'h5dc;
        src123 <= 12'hc1b;
        src124 <= 12'hb74;
        src125 <= 12'h168;
        src126 <= 12'ha8a;
        src127 <= 12'h7b1;
        src128 <= 12'hbe3;
        src129 <= 12'hef2;
        src130 <= 12'h536;
        src131 <= 12'hb3;
        src132 <= 12'hea6;
        src133 <= 12'he1d;
        src134 <= 12'h2fc;
        src135 <= 12'h8f8;
        src136 <= 12'hf37;
        src137 <= 12'h45;
        src138 <= 12'hbe2;
        src139 <= 12'h3bb;
        src140 <= 12'ha4e;
        src141 <= 12'h3f9;
        src142 <= 12'h77c;
        src143 <= 12'hf50;
        src144 <= 12'h17;
        src145 <= 12'h71;
        src146 <= 12'h9de;
        src147 <= 12'hb04;
        src148 <= 12'h654;
        src149 <= 12'h30e;
        src150 <= 12'he4b;
        src151 <= 12'he21;
        src152 <= 12'h8a5;
        src153 <= 12'h1bb;
        src154 <= 12'hb46;
        src155 <= 12'h6a2;
        src156 <= 12'haa0;
        src157 <= 12'h681;
        src158 <= 12'h46;
        src159 <= 12'haae;
        src160 <= 12'hd9;
        src161 <= 12'hbba;
        exp <= 20'h4f23b;
        #1
        src0 <= 12'h86a;
        src1 <= 12'h1f0;
        src2 <= 12'h5cb;
        src3 <= 12'h592;
        src4 <= 12'h28e;
        src5 <= 12'hd6a;
        src6 <= 12'h480;
        src7 <= 12'h252;
        src8 <= 12'had;
        src9 <= 12'h7ba;
        src10 <= 12'hf49;
        src11 <= 12'ha43;
        src12 <= 12'hda6;
        src13 <= 12'hcae;
        src14 <= 12'ha0f;
        src15 <= 12'hb5d;
        src16 <= 12'hb31;
        src17 <= 12'h8ac;
        src18 <= 12'h5b5;
        src19 <= 12'hf2d;
        src20 <= 12'ha2;
        src21 <= 12'h58b;
        src22 <= 12'h412;
        src23 <= 12'h4c6;
        src24 <= 12'h491;
        src25 <= 12'h4c9;
        src26 <= 12'h6cc;
        src27 <= 12'h4ed;
        src28 <= 12'h188;
        src29 <= 12'he55;
        src30 <= 12'h732;
        src31 <= 12'h91b;
        src32 <= 12'h539;
        src33 <= 12'hcf6;
        src34 <= 12'h3f4;
        src35 <= 12'hca2;
        src36 <= 12'h146;
        src37 <= 12'h997;
        src38 <= 12'h681;
        src39 <= 12'ha6d;
        src40 <= 12'hf32;
        src41 <= 12'haf;
        src42 <= 12'hc7d;
        src43 <= 12'hafc;
        src44 <= 12'h65d;
        src45 <= 12'h5f3;
        src46 <= 12'hade;
        src47 <= 12'hd15;
        src48 <= 12'h5ed;
        src49 <= 12'hcaa;
        src50 <= 12'he72;
        src51 <= 12'h89e;
        src52 <= 12'ha44;
        src53 <= 12'h932;
        src54 <= 12'h52a;
        src55 <= 12'h8e4;
        src56 <= 12'ha6a;
        src57 <= 12'h5d2;
        src58 <= 12'hc46;
        src59 <= 12'h34d;
        src60 <= 12'h457;
        src61 <= 12'h615;
        src62 <= 12'h638;
        src63 <= 12'h6ed;
        src64 <= 12'hc46;
        src65 <= 12'hdb6;
        src66 <= 12'h42;
        src67 <= 12'h6da;
        src68 <= 12'hc33;
        src69 <= 12'h434;
        src70 <= 12'h885;
        src71 <= 12'he93;
        src72 <= 12'h274;
        src73 <= 12'h5e7;
        src74 <= 12'hf2d;
        src75 <= 12'he10;
        src76 <= 12'hfe9;
        src77 <= 12'h292;
        src78 <= 12'h5b2;
        src79 <= 12'h1ca;
        src80 <= 12'h2e5;
        src81 <= 12'hdb0;
        src82 <= 12'h4e6;
        src83 <= 12'h1f2;
        src84 <= 12'hcc8;
        src85 <= 12'hbfe;
        src86 <= 12'hdbb;
        src87 <= 12'h851;
        src88 <= 12'hd2e;
        src89 <= 12'h5cd;
        src90 <= 12'h5ae;
        src91 <= 12'hd05;
        src92 <= 12'hbe6;
        src93 <= 12'h698;
        src94 <= 12'h6ab;
        src95 <= 12'h8bf;
        src96 <= 12'h52d;
        src97 <= 12'h4cd;
        src98 <= 12'h69d;
        src99 <= 12'h81a;
        src100 <= 12'h557;
        src101 <= 12'heea;
        src102 <= 12'h231;
        src103 <= 12'h75e;
        src104 <= 12'h34c;
        src105 <= 12'h5a7;
        src106 <= 12'ha77;
        src107 <= 12'he93;
        src108 <= 12'h719;
        src109 <= 12'hb25;
        src110 <= 12'h8ee;
        src111 <= 12'hfd2;
        src112 <= 12'ha51;
        src113 <= 12'hf00;
        src114 <= 12'h502;
        src115 <= 12'ha88;
        src116 <= 12'h2cd;
        src117 <= 12'ha47;
        src118 <= 12'he4c;
        src119 <= 12'ha20;
        src120 <= 12'h57e;
        src121 <= 12'hcc5;
        src122 <= 12'hba9;
        src123 <= 12'ha4a;
        src124 <= 12'hc28;
        src125 <= 12'hbda;
        src126 <= 12'h5df;
        src127 <= 12'h145;
        src128 <= 12'hb63;
        src129 <= 12'h4fd;
        src130 <= 12'h88a;
        src131 <= 12'hdbe;
        src132 <= 12'h5c;
        src133 <= 12'h3f1;
        src134 <= 12'hddb;
        src135 <= 12'hed3;
        src136 <= 12'hdf5;
        src137 <= 12'h7e2;
        src138 <= 12'hcf5;
        src139 <= 12'ha3a;
        src140 <= 12'he44;
        src141 <= 12'hc9f;
        src142 <= 12'hdad;
        src143 <= 12'h7da;
        src144 <= 12'hf66;
        src145 <= 12'h98;
        src146 <= 12'h1d2;
        src147 <= 12'h2a;
        src148 <= 12'h615;
        src149 <= 12'h6ec;
        src150 <= 12'ha66;
        src151 <= 12'h194;
        src152 <= 12'hb08;
        src153 <= 12'h15c;
        src154 <= 12'hff;
        src155 <= 12'h244;
        src156 <= 12'ha3d;
        src157 <= 12'h872;
        src158 <= 12'h5e5;
        src159 <= 12'hf1c;
        src160 <= 12'h1b4;
        src161 <= 12'haef;
        exp <= 20'h53b1d;
        #1
        src0 <= 12'hf92;
        src1 <= 12'h35b;
        src2 <= 12'h17d;
        src3 <= 12'hf4d;
        src4 <= 12'h677;
        src5 <= 12'h47;
        src6 <= 12'h75;
        src7 <= 12'h8ce;
        src8 <= 12'h6d1;
        src9 <= 12'h7d;
        src10 <= 12'h7d2;
        src11 <= 12'h575;
        src12 <= 12'ha0b;
        src13 <= 12'hfa2;
        src14 <= 12'hfc8;
        src15 <= 12'hafd;
        src16 <= 12'hac;
        src17 <= 12'hb1d;
        src18 <= 12'h7b4;
        src19 <= 12'hfc5;
        src20 <= 12'h968;
        src21 <= 12'h9d8;
        src22 <= 12'he77;
        src23 <= 12'haf3;
        src24 <= 12'h6ca;
        src25 <= 12'h720;
        src26 <= 12'hf00;
        src27 <= 12'hd95;
        src28 <= 12'h1;
        src29 <= 12'h38b;
        src30 <= 12'hbb0;
        src31 <= 12'ha17;
        src32 <= 12'hf23;
        src33 <= 12'h577;
        src34 <= 12'hb8b;
        src35 <= 12'h662;
        src36 <= 12'he71;
        src37 <= 12'h94c;
        src38 <= 12'h1ff;
        src39 <= 12'ha8f;
        src40 <= 12'h32e;
        src41 <= 12'he57;
        src42 <= 12'h82b;
        src43 <= 12'hf63;
        src44 <= 12'ha5c;
        src45 <= 12'h269;
        src46 <= 12'h2f3;
        src47 <= 12'ha0;
        src48 <= 12'hfa9;
        src49 <= 12'h420;
        src50 <= 12'h429;
        src51 <= 12'hac4;
        src52 <= 12'h9f0;
        src53 <= 12'hebe;
        src54 <= 12'h3a0;
        src55 <= 12'h86e;
        src56 <= 12'h549;
        src57 <= 12'hfde;
        src58 <= 12'h7d;
        src59 <= 12'h8d9;
        src60 <= 12'hedd;
        src61 <= 12'h97f;
        src62 <= 12'hcf4;
        src63 <= 12'hc99;
        src64 <= 12'hb68;
        src65 <= 12'h40d;
        src66 <= 12'h520;
        src67 <= 12'hcad;
        src68 <= 12'h931;
        src69 <= 12'h1a1;
        src70 <= 12'hd29;
        src71 <= 12'h896;
        src72 <= 12'h6e7;
        src73 <= 12'hf73;
        src74 <= 12'h886;
        src75 <= 12'hf96;
        src76 <= 12'h35c;
        src77 <= 12'h72f;
        src78 <= 12'he75;
        src79 <= 12'h3f3;
        src80 <= 12'h295;
        src81 <= 12'h1de;
        src82 <= 12'hc27;
        src83 <= 12'h571;
        src84 <= 12'hc06;
        src85 <= 12'h2d7;
        src86 <= 12'h2aa;
        src87 <= 12'h207;
        src88 <= 12'h861;
        src89 <= 12'hbe8;
        src90 <= 12'h586;
        src91 <= 12'h35f;
        src92 <= 12'h4f0;
        src93 <= 12'hb2e;
        src94 <= 12'hb3f;
        src95 <= 12'hcf9;
        src96 <= 12'hdaa;
        src97 <= 12'h8c8;
        src98 <= 12'h448;
        src99 <= 12'hcc7;
        src100 <= 12'h6ae;
        src101 <= 12'h60;
        src102 <= 12'h849;
        src103 <= 12'hb25;
        src104 <= 12'h61d;
        src105 <= 12'hf1d;
        src106 <= 12'h568;
        src107 <= 12'hbd6;
        src108 <= 12'hcce;
        src109 <= 12'h561;
        src110 <= 12'h1e9;
        src111 <= 12'hdd2;
        src112 <= 12'h2d2;
        src113 <= 12'h8e7;
        src114 <= 12'h24b;
        src115 <= 12'h38a;
        src116 <= 12'h3b;
        src117 <= 12'hcc8;
        src118 <= 12'hff7;
        src119 <= 12'h8c9;
        src120 <= 12'hdd;
        src121 <= 12'h2da;
        src122 <= 12'h258;
        src123 <= 12'h6d6;
        src124 <= 12'h721;
        src125 <= 12'hcf1;
        src126 <= 12'hd3f;
        src127 <= 12'h65;
        src128 <= 12'hb32;
        src129 <= 12'h8c7;
        src130 <= 12'h816;
        src131 <= 12'h46a;
        src132 <= 12'he70;
        src133 <= 12'hefb;
        src134 <= 12'h70a;
        src135 <= 12'h33f;
        src136 <= 12'hc85;
        src137 <= 12'hbd8;
        src138 <= 12'h81f;
        src139 <= 12'hd02;
        src140 <= 12'h386;
        src141 <= 12'h29b;
        src142 <= 12'h9e3;
        src143 <= 12'h769;
        src144 <= 12'h1aa;
        src145 <= 12'h30f;
        src146 <= 12'h567;
        src147 <= 12'h53b;
        src148 <= 12'h7dc;
        src149 <= 12'h5ce;
        src150 <= 12'hb01;
        src151 <= 12'h136;
        src152 <= 12'hcdf;
        src153 <= 12'h57c;
        src154 <= 12'hfc7;
        src155 <= 12'h761;
        src156 <= 12'h19a;
        src157 <= 12'h652;
        src158 <= 12'h173;
        src159 <= 12'h177;
        src160 <= 12'h6a9;
        src161 <= 12'h25e;
        exp <= 20'h50cea;
        #1
        src0 <= 12'h2e2;
        src1 <= 12'h3c6;
        src2 <= 12'h1d7;
        src3 <= 12'hfa0;
        src4 <= 12'hf;
        src5 <= 12'h3f9;
        src6 <= 12'had2;
        src7 <= 12'h832;
        src8 <= 12'h172;
        src9 <= 12'h37c;
        src10 <= 12'h84d;
        src11 <= 12'h40c;
        src12 <= 12'h965;
        src13 <= 12'h391;
        src14 <= 12'h7bc;
        src15 <= 12'h9bc;
        src16 <= 12'h3d3;
        src17 <= 12'h350;
        src18 <= 12'he25;
        src19 <= 12'h9e6;
        src20 <= 12'h88b;
        src21 <= 12'h538;
        src22 <= 12'h191;
        src23 <= 12'h7c5;
        src24 <= 12'h817;
        src25 <= 12'hb09;
        src26 <= 12'h120;
        src27 <= 12'hecf;
        src28 <= 12'h9f6;
        src29 <= 12'h392;
        src30 <= 12'hce;
        src31 <= 12'hd3;
        src32 <= 12'h6d5;
        src33 <= 12'h651;
        src34 <= 12'hdbc;
        src35 <= 12'hdb3;
        src36 <= 12'hb2e;
        src37 <= 12'h6a6;
        src38 <= 12'hfa9;
        src39 <= 12'h3fa;
        src40 <= 12'h94f;
        src41 <= 12'h1ed;
        src42 <= 12'h3ba;
        src43 <= 12'h8ed;
        src44 <= 12'h1a7;
        src45 <= 12'hb01;
        src46 <= 12'h79b;
        src47 <= 12'h883;
        src48 <= 12'hd1e;
        src49 <= 12'hcf6;
        src50 <= 12'h83c;
        src51 <= 12'h46a;
        src52 <= 12'h425;
        src53 <= 12'h644;
        src54 <= 12'h802;
        src55 <= 12'h3a8;
        src56 <= 12'h3f7;
        src57 <= 12'h7a3;
        src58 <= 12'hf27;
        src59 <= 12'h221;
        src60 <= 12'haab;
        src61 <= 12'h68a;
        src62 <= 12'h768;
        src63 <= 12'hef0;
        src64 <= 12'h24c;
        src65 <= 12'h2aa;
        src66 <= 12'h224;
        src67 <= 12'hf20;
        src68 <= 12'h185;
        src69 <= 12'h669;
        src70 <= 12'h5c;
        src71 <= 12'h865;
        src72 <= 12'h3a1;
        src73 <= 12'hf77;
        src74 <= 12'hd40;
        src75 <= 12'hb4d;
        src76 <= 12'hdce;
        src77 <= 12'h955;
        src78 <= 12'h537;
        src79 <= 12'h109;
        src80 <= 12'h76d;
        src81 <= 12'hdef;
        src82 <= 12'h94a;
        src83 <= 12'h1c8;
        src84 <= 12'h501;
        src85 <= 12'hfa4;
        src86 <= 12'heb;
        src87 <= 12'h6e6;
        src88 <= 12'h238;
        src89 <= 12'hef4;
        src90 <= 12'hc26;
        src91 <= 12'h46a;
        src92 <= 12'h436;
        src93 <= 12'hc67;
        src94 <= 12'h454;
        src95 <= 12'h18f;
        src96 <= 12'hc11;
        src97 <= 12'hed8;
        src98 <= 12'hf1b;
        src99 <= 12'hd7c;
        src100 <= 12'h728;
        src101 <= 12'h591;
        src102 <= 12'h3e3;
        src103 <= 12'hb9f;
        src104 <= 12'hd89;
        src105 <= 12'h564;
        src106 <= 12'h60f;
        src107 <= 12'hd8c;
        src108 <= 12'h76;
        src109 <= 12'ha1c;
        src110 <= 12'h447;
        src111 <= 12'h7f;
        src112 <= 12'hcf;
        src113 <= 12'hcc9;
        src114 <= 12'h539;
        src115 <= 12'hd24;
        src116 <= 12'hcbc;
        src117 <= 12'h47e;
        src118 <= 12'h48b;
        src119 <= 12'h6cc;
        src120 <= 12'hfcb;
        src121 <= 12'haf3;
        src122 <= 12'hd75;
        src123 <= 12'h9fb;
        src124 <= 12'h343;
        src125 <= 12'h1b0;
        src126 <= 12'hfee;
        src127 <= 12'hef0;
        src128 <= 12'hc68;
        src129 <= 12'hced;
        src130 <= 12'h3ca;
        src131 <= 12'h7d5;
        src132 <= 12'h19b;
        src133 <= 12'h3c5;
        src134 <= 12'hfaf;
        src135 <= 12'hae1;
        src136 <= 12'hfe5;
        src137 <= 12'hf85;
        src138 <= 12'h16b;
        src139 <= 12'hde9;
        src140 <= 12'h3c7;
        src141 <= 12'h39a;
        src142 <= 12'h3cc;
        src143 <= 12'ha7b;
        src144 <= 12'h495;
        src145 <= 12'h109;
        src146 <= 12'ha8a;
        src147 <= 12'hcea;
        src148 <= 12'h9e7;
        src149 <= 12'h242;
        src150 <= 12'he56;
        src151 <= 12'hd05;
        src152 <= 12'h174;
        src153 <= 12'h585;
        src154 <= 12'h8e4;
        src155 <= 12'h50e;
        src156 <= 12'h45a;
        src157 <= 12'ha40;
        src158 <= 12'h8af;
        src159 <= 12'h2b3;
        src160 <= 12'h109;
        src161 <= 12'hda9;
        exp <= 20'h4d7fa;
        #1
        src0 <= 12'he87;
        src1 <= 12'h35;
        src2 <= 12'he23;
        src3 <= 12'hf3b;
        src4 <= 12'h99b;
        src5 <= 12'hdc7;
        src6 <= 12'h6e7;
        src7 <= 12'h725;
        src8 <= 12'h22c;
        src9 <= 12'h55d;
        src10 <= 12'h50f;
        src11 <= 12'he7d;
        src12 <= 12'h3ee;
        src13 <= 12'h4d6;
        src14 <= 12'h849;
        src15 <= 12'h173;
        src16 <= 12'hfdd;
        src17 <= 12'h6b;
        src18 <= 12'h649;
        src19 <= 12'h123;
        src20 <= 12'h481;
        src21 <= 12'h1d0;
        src22 <= 12'h32;
        src23 <= 12'h5ec;
        src24 <= 12'h1d5;
        src25 <= 12'hb7d;
        src26 <= 12'h1bb;
        src27 <= 12'hd41;
        src28 <= 12'hbdb;
        src29 <= 12'hafd;
        src30 <= 12'h112;
        src31 <= 12'ha78;
        src32 <= 12'h432;
        src33 <= 12'h5d1;
        src34 <= 12'h19d;
        src35 <= 12'h733;
        src36 <= 12'he89;
        src37 <= 12'h6ba;
        src38 <= 12'hb92;
        src39 <= 12'h3f2;
        src40 <= 12'hb00;
        src41 <= 12'h4dc;
        src42 <= 12'ha43;
        src43 <= 12'h41;
        src44 <= 12'hcc9;
        src45 <= 12'h7dd;
        src46 <= 12'h4f5;
        src47 <= 12'hc51;
        src48 <= 12'h660;
        src49 <= 12'h459;
        src50 <= 12'hebf;
        src51 <= 12'h5c0;
        src52 <= 12'h78b;
        src53 <= 12'h4ac;
        src54 <= 12'h230;
        src55 <= 12'hacc;
        src56 <= 12'h25c;
        src57 <= 12'h44;
        src58 <= 12'h1d8;
        src59 <= 12'h81c;
        src60 <= 12'hb0f;
        src61 <= 12'ha53;
        src62 <= 12'hf67;
        src63 <= 12'hcd8;
        src64 <= 12'h4b7;
        src65 <= 12'hfcc;
        src66 <= 12'h743;
        src67 <= 12'h69c;
        src68 <= 12'ha2;
        src69 <= 12'h738;
        src70 <= 12'hde9;
        src71 <= 12'h3dc;
        src72 <= 12'h1a9;
        src73 <= 12'he0d;
        src74 <= 12'ha74;
        src75 <= 12'heb9;
        src76 <= 12'hcb3;
        src77 <= 12'h883;
        src78 <= 12'h89e;
        src79 <= 12'h6e2;
        src80 <= 12'hc7e;
        src81 <= 12'h30f;
        src82 <= 12'h391;
        src83 <= 12'hf0b;
        src84 <= 12'h32c;
        src85 <= 12'h1c5;
        src86 <= 12'h3bb;
        src87 <= 12'h8c;
        src88 <= 12'hf18;
        src89 <= 12'h210;
        src90 <= 12'hfde;
        src91 <= 12'hcaa;
        src92 <= 12'h911;
        src93 <= 12'hda2;
        src94 <= 12'hd9e;
        src95 <= 12'ha91;
        src96 <= 12'ha60;
        src97 <= 12'hddd;
        src98 <= 12'h9ed;
        src99 <= 12'hcf1;
        src100 <= 12'h19b;
        src101 <= 12'hebc;
        src102 <= 12'h401;
        src103 <= 12'hc;
        src104 <= 12'hc7d;
        src105 <= 12'h9e6;
        src106 <= 12'h749;
        src107 <= 12'hc5b;
        src108 <= 12'h242;
        src109 <= 12'hbbe;
        src110 <= 12'h728;
        src111 <= 12'h3ac;
        src112 <= 12'hdd7;
        src113 <= 12'h69d;
        src114 <= 12'hca0;
        src115 <= 12'he21;
        src116 <= 12'h1db;
        src117 <= 12'h667;
        src118 <= 12'h638;
        src119 <= 12'h6f3;
        src120 <= 12'h69c;
        src121 <= 12'h76e;
        src122 <= 12'hbed;
        src123 <= 12'hc84;
        src124 <= 12'hf0c;
        src125 <= 12'hbd3;
        src126 <= 12'hf88;
        src127 <= 12'h2b6;
        src128 <= 12'haf5;
        src129 <= 12'hb0e;
        src130 <= 12'h37b;
        src131 <= 12'hf06;
        src132 <= 12'h378;
        src133 <= 12'h5e8;
        src134 <= 12'hb1d;
        src135 <= 12'h5ca;
        src136 <= 12'h6b2;
        src137 <= 12'hcf1;
        src138 <= 12'h171;
        src139 <= 12'h6e9;
        src140 <= 12'hc03;
        src141 <= 12'h9f0;
        src142 <= 12'h264;
        src143 <= 12'h635;
        src144 <= 12'hd25;
        src145 <= 12'h7db;
        src146 <= 12'h3c0;
        src147 <= 12'hebf;
        src148 <= 12'h191;
        src149 <= 12'hb5e;
        src150 <= 12'hc4e;
        src151 <= 12'h9ca;
        src152 <= 12'hbee;
        src153 <= 12'h71d;
        src154 <= 12'h885;
        src155 <= 12'h62e;
        src156 <= 12'h827;
        src157 <= 12'hb04;
        src158 <= 12'hdab;
        src159 <= 12'hf60;
        src160 <= 12'h93b;
        src161 <= 12'hbbf;
        exp <= 20'h52f5f;
        #1
        src0 <= 12'h8bb;
        src1 <= 12'hcc7;
        src2 <= 12'hcc7;
        src3 <= 12'h9d5;
        src4 <= 12'h26a;
        src5 <= 12'h37a;
        src6 <= 12'h48e;
        src7 <= 12'hbe0;
        src8 <= 12'h2f9;
        src9 <= 12'hd6d;
        src10 <= 12'hafc;
        src11 <= 12'ha6c;
        src12 <= 12'hd33;
        src13 <= 12'h1ed;
        src14 <= 12'h91b;
        src15 <= 12'h7b9;
        src16 <= 12'h7f2;
        src17 <= 12'h930;
        src18 <= 12'h34c;
        src19 <= 12'h38;
        src20 <= 12'hf09;
        src21 <= 12'hd8f;
        src22 <= 12'hdcb;
        src23 <= 12'ha5f;
        src24 <= 12'h73c;
        src25 <= 12'had5;
        src26 <= 12'hc64;
        src27 <= 12'h6fa;
        src28 <= 12'h24;
        src29 <= 12'h4ae;
        src30 <= 12'ha38;
        src31 <= 12'he67;
        src32 <= 12'hff0;
        src33 <= 12'h78a;
        src34 <= 12'h6c3;
        src35 <= 12'hdf0;
        src36 <= 12'h147;
        src37 <= 12'h158;
        src38 <= 12'h2f6;
        src39 <= 12'h804;
        src40 <= 12'h2d;
        src41 <= 12'h840;
        src42 <= 12'h116;
        src43 <= 12'h7e3;
        src44 <= 12'hc8;
        src45 <= 12'h477;
        src46 <= 12'h487;
        src47 <= 12'h903;
        src48 <= 12'h12;
        src49 <= 12'h739;
        src50 <= 12'h4f;
        src51 <= 12'h889;
        src52 <= 12'h4d4;
        src53 <= 12'h319;
        src54 <= 12'h336;
        src55 <= 12'h3b4;
        src56 <= 12'h698;
        src57 <= 12'h33;
        src58 <= 12'h6c8;
        src59 <= 12'h7a7;
        src60 <= 12'ha9c;
        src61 <= 12'hf1f;
        src62 <= 12'h18c;
        src63 <= 12'h238;
        src64 <= 12'h1f6;
        src65 <= 12'hd27;
        src66 <= 12'h84a;
        src67 <= 12'h7ff;
        src68 <= 12'hcd6;
        src69 <= 12'h8bd;
        src70 <= 12'hd99;
        src71 <= 12'h2db;
        src72 <= 12'h81;
        src73 <= 12'h68e;
        src74 <= 12'he71;
        src75 <= 12'h8b0;
        src76 <= 12'h857;
        src77 <= 12'h8d5;
        src78 <= 12'h589;
        src79 <= 12'h405;
        src80 <= 12'h535;
        src81 <= 12'hb54;
        src82 <= 12'hc70;
        src83 <= 12'h4cb;
        src84 <= 12'h4fc;
        src85 <= 12'h2d8;
        src86 <= 12'h14b;
        src87 <= 12'h8a3;
        src88 <= 12'h23f;
        src89 <= 12'hb57;
        src90 <= 12'hf0d;
        src91 <= 12'h6b5;
        src92 <= 12'heb9;
        src93 <= 12'hb61;
        src94 <= 12'hc02;
        src95 <= 12'hef;
        src96 <= 12'h27f;
        src97 <= 12'h513;
        src98 <= 12'ha7;
        src99 <= 12'hb2f;
        src100 <= 12'h13b;
        src101 <= 12'h41e;
        src102 <= 12'h60f;
        src103 <= 12'haff;
        src104 <= 12'h39d;
        src105 <= 12'hf38;
        src106 <= 12'hd6a;
        src107 <= 12'hf46;
        src108 <= 12'hebb;
        src109 <= 12'h303;
        src110 <= 12'h14c;
        src111 <= 12'h333;
        src112 <= 12'h477;
        src113 <= 12'h585;
        src114 <= 12'h67a;
        src115 <= 12'hfa7;
        src116 <= 12'ha11;
        src117 <= 12'had4;
        src118 <= 12'h929;
        src119 <= 12'hf9f;
        src120 <= 12'h179;
        src121 <= 12'h987;
        src122 <= 12'hcf6;
        src123 <= 12'h7f2;
        src124 <= 12'he6e;
        src125 <= 12'hf8e;
        src126 <= 12'h73b;
        src127 <= 12'h1fa;
        src128 <= 12'h7f7;
        src129 <= 12'ha30;
        src130 <= 12'h6de;
        src131 <= 12'h82b;
        src132 <= 12'h5e1;
        src133 <= 12'h796;
        src134 <= 12'h70b;
        src135 <= 12'h48f;
        src136 <= 12'hfc6;
        src137 <= 12'h37e;
        src138 <= 12'h5dd;
        src139 <= 12'h1c0;
        src140 <= 12'h874;
        src141 <= 12'h6d5;
        src142 <= 12'he42;
        src143 <= 12'h6d1;
        src144 <= 12'hb30;
        src145 <= 12'h605;
        src146 <= 12'h87b;
        src147 <= 12'h392;
        src148 <= 12'h94c;
        src149 <= 12'hee2;
        src150 <= 12'h401;
        src151 <= 12'h59b;
        src152 <= 12'h44b;
        src153 <= 12'h4b9;
        src154 <= 12'h763;
        src155 <= 12'h9a4;
        src156 <= 12'h30d;
        src157 <= 12'hb4c;
        src158 <= 12'h28f;
        src159 <= 12'h7d4;
        src160 <= 12'h389;
        src161 <= 12'h5d7;
        exp <= 20'h4b987;
        #1
        src0 <= 12'hb3d;
        src1 <= 12'h5b0;
        src2 <= 12'h9d6;
        src3 <= 12'hb0b;
        src4 <= 12'h671;
        src5 <= 12'h98a;
        src6 <= 12'h9e0;
        src7 <= 12'h832;
        src8 <= 12'h73d;
        src9 <= 12'h7ea;
        src10 <= 12'h9c3;
        src11 <= 12'h3d6;
        src12 <= 12'h537;
        src13 <= 12'h548;
        src14 <= 12'hbaf;
        src15 <= 12'h1a;
        src16 <= 12'h39b;
        src17 <= 12'h32f;
        src18 <= 12'h9c0;
        src19 <= 12'hc5c;
        src20 <= 12'h373;
        src21 <= 12'h263;
        src22 <= 12'h528;
        src23 <= 12'hcb8;
        src24 <= 12'h824;
        src25 <= 12'h6b1;
        src26 <= 12'h1c3;
        src27 <= 12'ha5f;
        src28 <= 12'h5b3;
        src29 <= 12'h74c;
        src30 <= 12'h9c0;
        src31 <= 12'h565;
        src32 <= 12'h2e0;
        src33 <= 12'hdbb;
        src34 <= 12'h243;
        src35 <= 12'h162;
        src36 <= 12'h70c;
        src37 <= 12'h9e4;
        src38 <= 12'hfdd;
        src39 <= 12'h9e;
        src40 <= 12'h870;
        src41 <= 12'hb52;
        src42 <= 12'hb54;
        src43 <= 12'heaf;
        src44 <= 12'heaa;
        src45 <= 12'h998;
        src46 <= 12'h43e;
        src47 <= 12'h804;
        src48 <= 12'h875;
        src49 <= 12'hc09;
        src50 <= 12'h9e9;
        src51 <= 12'h545;
        src52 <= 12'hfd1;
        src53 <= 12'h904;
        src54 <= 12'h949;
        src55 <= 12'hff4;
        src56 <= 12'h804;
        src57 <= 12'h185;
        src58 <= 12'hfa5;
        src59 <= 12'h1df;
        src60 <= 12'h84b;
        src61 <= 12'h19;
        src62 <= 12'h440;
        src63 <= 12'hd5a;
        src64 <= 12'h857;
        src65 <= 12'h4c5;
        src66 <= 12'h699;
        src67 <= 12'h714;
        src68 <= 12'hc15;
        src69 <= 12'h7ec;
        src70 <= 12'h8dd;
        src71 <= 12'hc94;
        src72 <= 12'h22b;
        src73 <= 12'haec;
        src74 <= 12'h7cc;
        src75 <= 12'h233;
        src76 <= 12'h463;
        src77 <= 12'h98e;
        src78 <= 12'hf02;
        src79 <= 12'h94;
        src80 <= 12'h95d;
        src81 <= 12'h807;
        src82 <= 12'h71a;
        src83 <= 12'h2aa;
        src84 <= 12'h6c9;
        src85 <= 12'h29f;
        src86 <= 12'h3da;
        src87 <= 12'hdd8;
        src88 <= 12'h4c5;
        src89 <= 12'h5ad;
        src90 <= 12'h89f;
        src91 <= 12'hbd0;
        src92 <= 12'he39;
        src93 <= 12'h9da;
        src94 <= 12'hcad;
        src95 <= 12'hd93;
        src96 <= 12'h90e;
        src97 <= 12'h17d;
        src98 <= 12'h6c8;
        src99 <= 12'h9c4;
        src100 <= 12'h15;
        src101 <= 12'h53;
        src102 <= 12'hc13;
        src103 <= 12'h271;
        src104 <= 12'h766;
        src105 <= 12'hdc0;
        src106 <= 12'h894;
        src107 <= 12'h6a8;
        src108 <= 12'h8f6;
        src109 <= 12'ha8;
        src110 <= 12'h718;
        src111 <= 12'hc69;
        src112 <= 12'h612;
        src113 <= 12'hbf9;
        src114 <= 12'hf4c;
        src115 <= 12'ha03;
        src116 <= 12'hf66;
        src117 <= 12'hddf;
        src118 <= 12'he95;
        src119 <= 12'hd49;
        src120 <= 12'h4f5;
        src121 <= 12'hfe2;
        src122 <= 12'hfe5;
        src123 <= 12'h25a;
        src124 <= 12'h4c;
        src125 <= 12'h59c;
        src126 <= 12'h383;
        src127 <= 12'h630;
        src128 <= 12'ha99;
        src129 <= 12'hd54;
        src130 <= 12'h898;
        src131 <= 12'h840;
        src132 <= 12'he35;
        src133 <= 12'hf75;
        src134 <= 12'h1ad;
        src135 <= 12'h7ab;
        src136 <= 12'h7f0;
        src137 <= 12'hba6;
        src138 <= 12'h339;
        src139 <= 12'h6c5;
        src140 <= 12'h83a;
        src141 <= 12'hd42;
        src142 <= 12'h72f;
        src143 <= 12'h639;
        src144 <= 12'h64c;
        src145 <= 12'h7fc;
        src146 <= 12'hf68;
        src147 <= 12'h72d;
        src148 <= 12'hd39;
        src149 <= 12'h3d5;
        src150 <= 12'ha36;
        src151 <= 12'h9b7;
        src152 <= 12'hbde;
        src153 <= 12'ha42;
        src154 <= 12'h8d1;
        src155 <= 12'h3a4;
        src156 <= 12'had0;
        src157 <= 12'h942;
        src158 <= 12'hc72;
        src159 <= 12'hf73;
        src160 <= 12'hbbb;
        src161 <= 12'hf62;
        exp <= 20'h54817;
        #1
        src0 <= 12'h37;
        src1 <= 12'h791;
        src2 <= 12'hd35;
        src3 <= 12'hfd5;
        src4 <= 12'h7d7;
        src5 <= 12'h2a;
        src6 <= 12'h592;
        src7 <= 12'hf3f;
        src8 <= 12'h36b;
        src9 <= 12'h636;
        src10 <= 12'hf44;
        src11 <= 12'hb03;
        src12 <= 12'h61e;
        src13 <= 12'h7dc;
        src14 <= 12'hcd8;
        src15 <= 12'h5d0;
        src16 <= 12'h353;
        src17 <= 12'hc70;
        src18 <= 12'h7f5;
        src19 <= 12'h814;
        src20 <= 12'h8e2;
        src21 <= 12'ha5c;
        src22 <= 12'hb5c;
        src23 <= 12'h3d3;
        src24 <= 12'h824;
        src25 <= 12'h167;
        src26 <= 12'h673;
        src27 <= 12'hf1;
        src28 <= 12'h542;
        src29 <= 12'hdf1;
        src30 <= 12'h92e;
        src31 <= 12'habb;
        src32 <= 12'hf53;
        src33 <= 12'h13e;
        src34 <= 12'h27;
        src35 <= 12'h3a1;
        src36 <= 12'h6f8;
        src37 <= 12'hb16;
        src38 <= 12'h7a1;
        src39 <= 12'h34f;
        src40 <= 12'h76c;
        src41 <= 12'h2a5;
        src42 <= 12'ha33;
        src43 <= 12'hc29;
        src44 <= 12'h221;
        src45 <= 12'hea3;
        src46 <= 12'h48d;
        src47 <= 12'hff8;
        src48 <= 12'he56;
        src49 <= 12'h25a;
        src50 <= 12'hbac;
        src51 <= 12'h852;
        src52 <= 12'had1;
        src53 <= 12'hb83;
        src54 <= 12'hec8;
        src55 <= 12'h20d;
        src56 <= 12'h99c;
        src57 <= 12'h738;
        src58 <= 12'h5b3;
        src59 <= 12'h177;
        src60 <= 12'h6de;
        src61 <= 12'hc3a;
        src62 <= 12'h369;
        src63 <= 12'h4e4;
        src64 <= 12'hf96;
        src65 <= 12'h76f;
        src66 <= 12'h559;
        src67 <= 12'h4dc;
        src68 <= 12'h55c;
        src69 <= 12'h50d;
        src70 <= 12'h7b1;
        src71 <= 12'h65a;
        src72 <= 12'heaf;
        src73 <= 12'h128;
        src74 <= 12'h67e;
        src75 <= 12'hde;
        src76 <= 12'hc4b;
        src77 <= 12'h426;
        src78 <= 12'hd22;
        src79 <= 12'hb6c;
        src80 <= 12'h1f5;
        src81 <= 12'h22c;
        src82 <= 12'h9fe;
        src83 <= 12'h629;
        src84 <= 12'h2dc;
        src85 <= 12'h6b9;
        src86 <= 12'h506;
        src87 <= 12'he84;
        src88 <= 12'h43b;
        src89 <= 12'h243;
        src90 <= 12'hb08;
        src91 <= 12'h8f9;
        src92 <= 12'h72c;
        src93 <= 12'h7f8;
        src94 <= 12'h945;
        src95 <= 12'hcd1;
        src96 <= 12'hf56;
        src97 <= 12'he29;
        src98 <= 12'hc00;
        src99 <= 12'h92d;
        src100 <= 12'h4b7;
        src101 <= 12'ha06;
        src102 <= 12'hee4;
        src103 <= 12'h6be;
        src104 <= 12'hbb2;
        src105 <= 12'he6b;
        src106 <= 12'h47c;
        src107 <= 12'ha5f;
        src108 <= 12'hff4;
        src109 <= 12'h2ed;
        src110 <= 12'hbff;
        src111 <= 12'h89a;
        src112 <= 12'h7ea;
        src113 <= 12'h2d7;
        src114 <= 12'hdce;
        src115 <= 12'hba8;
        src116 <= 12'he1;
        src117 <= 12'h288;
        src118 <= 12'hb82;
        src119 <= 12'h4a;
        src120 <= 12'h382;
        src121 <= 12'hae3;
        src122 <= 12'h414;
        src123 <= 12'hd;
        src124 <= 12'h501;
        src125 <= 12'ha6;
        src126 <= 12'h650;
        src127 <= 12'hdc7;
        src128 <= 12'hbdd;
        src129 <= 12'hb0;
        src130 <= 12'hc65;
        src131 <= 12'he09;
        src132 <= 12'hc33;
        src133 <= 12'h678;
        src134 <= 12'hedc;
        src135 <= 12'hba8;
        src136 <= 12'h222;
        src137 <= 12'h2d1;
        src138 <= 12'h8fd;
        src139 <= 12'hcb7;
        src140 <= 12'ha2d;
        src141 <= 12'hb2a;
        src142 <= 12'h777;
        src143 <= 12'hd4;
        src144 <= 12'h831;
        src145 <= 12'hd16;
        src146 <= 12'h1f;
        src147 <= 12'hc30;
        src148 <= 12'he4d;
        src149 <= 12'h47b;
        src150 <= 12'h1a4;
        src151 <= 12'h9dc;
        src152 <= 12'h8a;
        src153 <= 12'h4f5;
        src154 <= 12'hbe3;
        src155 <= 12'h73;
        src156 <= 12'hae8;
        src157 <= 12'hbbb;
        src158 <= 12'hc17;
        src159 <= 12'hd44;
        src160 <= 12'hbb0;
        src161 <= 12'hf2e;
        exp <= 20'h511e8;
        #1
        src0 <= 12'h8d7;
        src1 <= 12'hfa8;
        src2 <= 12'ha6d;
        src3 <= 12'h4f2;
        src4 <= 12'hff8;
        src5 <= 12'h38a;
        src6 <= 12'hbac;
        src7 <= 12'h7ae;
        src8 <= 12'hd76;
        src9 <= 12'h2f4;
        src10 <= 12'h4ed;
        src11 <= 12'h805;
        src12 <= 12'h1d9;
        src13 <= 12'h65e;
        src14 <= 12'h956;
        src15 <= 12'ha70;
        src16 <= 12'h3ab;
        src17 <= 12'hb66;
        src18 <= 12'h153;
        src19 <= 12'hf1b;
        src20 <= 12'heb4;
        src21 <= 12'h433;
        src22 <= 12'h7dd;
        src23 <= 12'he91;
        src24 <= 12'h441;
        src25 <= 12'h776;
        src26 <= 12'h715;
        src27 <= 12'h342;
        src28 <= 12'h4ea;
        src29 <= 12'h453;
        src30 <= 12'h27c;
        src31 <= 12'h8e8;
        src32 <= 12'h794;
        src33 <= 12'h90f;
        src34 <= 12'h2d3;
        src35 <= 12'h1b3;
        src36 <= 12'h2e6;
        src37 <= 12'hde9;
        src38 <= 12'hc74;
        src39 <= 12'hbd6;
        src40 <= 12'h1a6;
        src41 <= 12'hd0d;
        src42 <= 12'h8d4;
        src43 <= 12'h7dd;
        src44 <= 12'hd19;
        src45 <= 12'h97c;
        src46 <= 12'hb46;
        src47 <= 12'h420;
        src48 <= 12'h6ac;
        src49 <= 12'h8f0;
        src50 <= 12'h1d5;
        src51 <= 12'h832;
        src52 <= 12'ha30;
        src53 <= 12'h973;
        src54 <= 12'hfeb;
        src55 <= 12'hacc;
        src56 <= 12'h385;
        src57 <= 12'hd8d;
        src58 <= 12'h6c6;
        src59 <= 12'he7d;
        src60 <= 12'h4fa;
        src61 <= 12'h2d;
        src62 <= 12'h4a8;
        src63 <= 12'hc06;
        src64 <= 12'hd3c;
        src65 <= 12'hc7c;
        src66 <= 12'h33d;
        src67 <= 12'he47;
        src68 <= 12'hfd9;
        src69 <= 12'h8c;
        src70 <= 12'h327;
        src71 <= 12'hc7c;
        src72 <= 12'h1e3;
        src73 <= 12'h8c;
        src74 <= 12'hd8d;
        src75 <= 12'h3ba;
        src76 <= 12'ha79;
        src77 <= 12'hbfc;
        src78 <= 12'h1dc;
        src79 <= 12'hb06;
        src80 <= 12'hc29;
        src81 <= 12'h681;
        src82 <= 12'hf47;
        src83 <= 12'h193;
        src84 <= 12'hbca;
        src85 <= 12'h691;
        src86 <= 12'h9d8;
        src87 <= 12'h976;
        src88 <= 12'h8ae;
        src89 <= 12'h137;
        src90 <= 12'h46a;
        src91 <= 12'hf14;
        src92 <= 12'hfc8;
        src93 <= 12'hfd9;
        src94 <= 12'h1d4;
        src95 <= 12'hbbd;
        src96 <= 12'h2df;
        src97 <= 12'h5bd;
        src98 <= 12'hc92;
        src99 <= 12'h427;
        src100 <= 12'h314;
        src101 <= 12'h3cb;
        src102 <= 12'he3b;
        src103 <= 12'ha74;
        src104 <= 12'h2e1;
        src105 <= 12'hbb2;
        src106 <= 12'hef4;
        src107 <= 12'h85f;
        src108 <= 12'h383;
        src109 <= 12'h543;
        src110 <= 12'h32;
        src111 <= 12'h88a;
        src112 <= 12'hcfa;
        src113 <= 12'h7b2;
        src114 <= 12'hec3;
        src115 <= 12'h82c;
        src116 <= 12'h1a5;
        src117 <= 12'h9e1;
        src118 <= 12'hd21;
        src119 <= 12'h6b3;
        src120 <= 12'h709;
        src121 <= 12'ha1;
        src122 <= 12'hbb0;
        src123 <= 12'hdda;
        src124 <= 12'h4c3;
        src125 <= 12'hc94;
        src126 <= 12'h304;
        src127 <= 12'hf;
        src128 <= 12'h159;
        src129 <= 12'hea3;
        src130 <= 12'h35d;
        src131 <= 12'h3db;
        src132 <= 12'hda1;
        src133 <= 12'h2e3;
        src134 <= 12'h819;
        src135 <= 12'hfe1;
        src136 <= 12'he3a;
        src137 <= 12'h4c0;
        src138 <= 12'h46c;
        src139 <= 12'h96;
        src140 <= 12'hd83;
        src141 <= 12'h68;
        src142 <= 12'hd95;
        src143 <= 12'h5b4;
        src144 <= 12'h3ed;
        src145 <= 12'hc67;
        src146 <= 12'h8c7;
        src147 <= 12'hb09;
        src148 <= 12'hc53;
        src149 <= 12'hf2d;
        src150 <= 12'h2a4;
        src151 <= 12'ha40;
        src152 <= 12'h16a;
        src153 <= 12'h10d;
        src154 <= 12'h188;
        src155 <= 12'ha92;
        src156 <= 12'hec2;
        src157 <= 12'h9eb;
        src158 <= 12'h940;
        src159 <= 12'ha30;
        src160 <= 12'hb14;
        src161 <= 12'h21e;
        exp <= 20'h51799;
        #1
        src0 <= 12'h747;
        src1 <= 12'h9a7;
        src2 <= 12'hd33;
        src3 <= 12'hf5d;
        src4 <= 12'h110;
        src5 <= 12'h39;
        src6 <= 12'h959;
        src7 <= 12'haa1;
        src8 <= 12'h8b4;
        src9 <= 12'hc4;
        src10 <= 12'hc8f;
        src11 <= 12'hc4f;
        src12 <= 12'h2ff;
        src13 <= 12'h928;
        src14 <= 12'hd4a;
        src15 <= 12'hb12;
        src16 <= 12'he97;
        src17 <= 12'h79f;
        src18 <= 12'h64;
        src19 <= 12'h4b7;
        src20 <= 12'h1e9;
        src21 <= 12'h585;
        src22 <= 12'hf0b;
        src23 <= 12'h714;
        src24 <= 12'h294;
        src25 <= 12'h2b0;
        src26 <= 12'h77c;
        src27 <= 12'hfa8;
        src28 <= 12'hc1f;
        src29 <= 12'ha3c;
        src30 <= 12'h3b7;
        src31 <= 12'hecc;
        src32 <= 12'hb09;
        src33 <= 12'h946;
        src34 <= 12'hcd4;
        src35 <= 12'hbd5;
        src36 <= 12'h265;
        src37 <= 12'h7c1;
        src38 <= 12'h856;
        src39 <= 12'h17a;
        src40 <= 12'h438;
        src41 <= 12'hb12;
        src42 <= 12'h6a;
        src43 <= 12'hb15;
        src44 <= 12'h6b0;
        src45 <= 12'hb32;
        src46 <= 12'h582;
        src47 <= 12'ha7d;
        src48 <= 12'ha96;
        src49 <= 12'h913;
        src50 <= 12'hf3d;
        src51 <= 12'h27f;
        src52 <= 12'h93c;
        src53 <= 12'h89c;
        src54 <= 12'h157;
        src55 <= 12'h9bc;
        src56 <= 12'h468;
        src57 <= 12'hf41;
        src58 <= 12'h314;
        src59 <= 12'hfb0;
        src60 <= 12'ha50;
        src61 <= 12'ha3a;
        src62 <= 12'h13b;
        src63 <= 12'h80;
        src64 <= 12'h565;
        src65 <= 12'ha21;
        src66 <= 12'h3cf;
        src67 <= 12'hae8;
        src68 <= 12'hc57;
        src69 <= 12'h2e2;
        src70 <= 12'h6ef;
        src71 <= 12'h3b4;
        src72 <= 12'h92c;
        src73 <= 12'h282;
        src74 <= 12'h782;
        src75 <= 12'h841;
        src76 <= 12'hdb2;
        src77 <= 12'h23e;
        src78 <= 12'h105;
        src79 <= 12'hb1f;
        src80 <= 12'hba9;
        src81 <= 12'h55d;
        src82 <= 12'h8ac;
        src83 <= 12'hcfc;
        src84 <= 12'h46a;
        src85 <= 12'h1d;
        src86 <= 12'hfbe;
        src87 <= 12'h467;
        src88 <= 12'heee;
        src89 <= 12'h688;
        src90 <= 12'h73f;
        src91 <= 12'h926;
        src92 <= 12'h2f7;
        src93 <= 12'h906;
        src94 <= 12'h9e0;
        src95 <= 12'h84f;
        src96 <= 12'hb98;
        src97 <= 12'hb63;
        src98 <= 12'h4e0;
        src99 <= 12'h25b;
        src100 <= 12'hbec;
        src101 <= 12'h8f9;
        src102 <= 12'h62b;
        src103 <= 12'h50b;
        src104 <= 12'h4e0;
        src105 <= 12'h40d;
        src106 <= 12'h460;
        src107 <= 12'hf85;
        src108 <= 12'h7da;
        src109 <= 12'h862;
        src110 <= 12'h1de;
        src111 <= 12'had4;
        src112 <= 12'he8e;
        src113 <= 12'hd62;
        src114 <= 12'hade;
        src115 <= 12'hc2e;
        src116 <= 12'h61f;
        src117 <= 12'h9d;
        src118 <= 12'heba;
        src119 <= 12'hc35;
        src120 <= 12'ha3c;
        src121 <= 12'h619;
        src122 <= 12'h84d;
        src123 <= 12'h395;
        src124 <= 12'he4d;
        src125 <= 12'hbf1;
        src126 <= 12'h940;
        src127 <= 12'h336;
        src128 <= 12'h24e;
        src129 <= 12'h640;
        src130 <= 12'h379;
        src131 <= 12'h527;
        src132 <= 12'h55e;
        src133 <= 12'h96c;
        src134 <= 12'h41e;
        src135 <= 12'h494;
        src136 <= 12'h1d5;
        src137 <= 12'h3bd;
        src138 <= 12'hb6;
        src139 <= 12'h4dc;
        src140 <= 12'h7c0;
        src141 <= 12'h35a;
        src142 <= 12'h9ad;
        src143 <= 12'hb1c;
        src144 <= 12'h86c;
        src145 <= 12'h87;
        src146 <= 12'h40d;
        src147 <= 12'hae3;
        src148 <= 12'hb12;
        src149 <= 12'hda4;
        src150 <= 12'hb2;
        src151 <= 12'h271;
        src152 <= 12'hf75;
        src153 <= 12'hbab;
        src154 <= 12'haaf;
        src155 <= 12'hab0;
        src156 <= 12'h6db;
        src157 <= 12'hdac;
        src158 <= 12'hd09;
        src159 <= 12'hd4c;
        src160 <= 12'h24b;
        src161 <= 12'hf1e;
        exp <= 20'h4ff2b;
        #1
        src0 <= 12'h14f;
        src1 <= 12'ha46;
        src2 <= 12'h827;
        src3 <= 12'h4ec;
        src4 <= 12'h2b4;
        src5 <= 12'h6e7;
        src6 <= 12'h140;
        src7 <= 12'h3de;
        src8 <= 12'hb78;
        src9 <= 12'hdc1;
        src10 <= 12'hcc;
        src11 <= 12'h972;
        src12 <= 12'h99c;
        src13 <= 12'hdde;
        src14 <= 12'he2a;
        src15 <= 12'h231;
        src16 <= 12'hbe1;
        src17 <= 12'hf16;
        src18 <= 12'h68b;
        src19 <= 12'hf3b;
        src20 <= 12'h77d;
        src21 <= 12'h7ee;
        src22 <= 12'h9b3;
        src23 <= 12'hd91;
        src24 <= 12'h6d3;
        src25 <= 12'hdfe;
        src26 <= 12'h9fc;
        src27 <= 12'he02;
        src28 <= 12'h682;
        src29 <= 12'h159;
        src30 <= 12'hc7d;
        src31 <= 12'hcc0;
        src32 <= 12'h4dd;
        src33 <= 12'h7a9;
        src34 <= 12'h6a2;
        src35 <= 12'hac5;
        src36 <= 12'h9c3;
        src37 <= 12'h85c;
        src38 <= 12'hb72;
        src39 <= 12'hd31;
        src40 <= 12'hbd3;
        src41 <= 12'hffa;
        src42 <= 12'hd69;
        src43 <= 12'ha6b;
        src44 <= 12'hb79;
        src45 <= 12'h544;
        src46 <= 12'he67;
        src47 <= 12'h596;
        src48 <= 12'hc73;
        src49 <= 12'hd77;
        src50 <= 12'he48;
        src51 <= 12'h6b1;
        src52 <= 12'hd09;
        src53 <= 12'hab3;
        src54 <= 12'h6b2;
        src55 <= 12'h9e8;
        src56 <= 12'h50b;
        src57 <= 12'hcd5;
        src58 <= 12'h3b2;
        src59 <= 12'h22f;
        src60 <= 12'h581;
        src61 <= 12'hc90;
        src62 <= 12'hb4a;
        src63 <= 12'h1a4;
        src64 <= 12'hb26;
        src65 <= 12'h847;
        src66 <= 12'hf60;
        src67 <= 12'hf1;
        src68 <= 12'hf6b;
        src69 <= 12'hf51;
        src70 <= 12'hfdd;
        src71 <= 12'h59;
        src72 <= 12'h487;
        src73 <= 12'h14e;
        src74 <= 12'hef7;
        src75 <= 12'h282;
        src76 <= 12'h5f1;
        src77 <= 12'h370;
        src78 <= 12'hffe;
        src79 <= 12'h1b4;
        src80 <= 12'h1c8;
        src81 <= 12'hdea;
        src82 <= 12'hb79;
        src83 <= 12'h9df;
        src84 <= 12'hd76;
        src85 <= 12'he96;
        src86 <= 12'hdf5;
        src87 <= 12'hdc2;
        src88 <= 12'hfd0;
        src89 <= 12'haad;
        src90 <= 12'h6ff;
        src91 <= 12'h7e;
        src92 <= 12'hffe;
        src93 <= 12'hfe9;
        src94 <= 12'h1f;
        src95 <= 12'h8ea;
        src96 <= 12'h45;
        src97 <= 12'ha3c;
        src98 <= 12'ha6c;
        src99 <= 12'h45e;
        src100 <= 12'hbdb;
        src101 <= 12'hefc;
        src102 <= 12'h657;
        src103 <= 12'h262;
        src104 <= 12'hcf1;
        src105 <= 12'h73e;
        src106 <= 12'hcaf;
        src107 <= 12'h8b8;
        src108 <= 12'hc0f;
        src109 <= 12'hdd2;
        src110 <= 12'hda1;
        src111 <= 12'hf56;
        src112 <= 12'h4ac;
        src113 <= 12'h54b;
        src114 <= 12'h412;
        src115 <= 12'h9a0;
        src116 <= 12'h1b0;
        src117 <= 12'h357;
        src118 <= 12'h3a;
        src119 <= 12'h2ff;
        src120 <= 12'h758;
        src121 <= 12'hcac;
        src122 <= 12'hd82;
        src123 <= 12'h899;
        src124 <= 12'hb96;
        src125 <= 12'h9a1;
        src126 <= 12'hbe2;
        src127 <= 12'h464;
        src128 <= 12'h6b2;
        src129 <= 12'h548;
        src130 <= 12'h13a;
        src131 <= 12'h5d9;
        src132 <= 12'h4f;
        src133 <= 12'h763;
        src134 <= 12'h6f;
        src135 <= 12'h258;
        src136 <= 12'h232;
        src137 <= 12'h537;
        src138 <= 12'h8fa;
        src139 <= 12'hbb6;
        src140 <= 12'hd1d;
        src141 <= 12'h379;
        src142 <= 12'hc48;
        src143 <= 12'hba2;
        src144 <= 12'he0;
        src145 <= 12'h884;
        src146 <= 12'h983;
        src147 <= 12'h106;
        src148 <= 12'hefc;
        src149 <= 12'haab;
        src150 <= 12'h375;
        src151 <= 12'h95b;
        src152 <= 12'h260;
        src153 <= 12'h535;
        src154 <= 12'h291;
        src155 <= 12'hfaa;
        src156 <= 12'ha34;
        src157 <= 12'h65b;
        src158 <= 12'h833;
        src159 <= 12'hd00;
        src160 <= 12'h271;
        src161 <= 12'h3ff;
        exp <= 20'h5631e;
        #1
        src0 <= 12'hdea;
        src1 <= 12'h778;
        src2 <= 12'hae0;
        src3 <= 12'hc15;
        src4 <= 12'he1c;
        src5 <= 12'h725;
        src6 <= 12'haad;
        src7 <= 12'h6c0;
        src8 <= 12'h5c0;
        src9 <= 12'h9ac;
        src10 <= 12'h0;
        src11 <= 12'h7e6;
        src12 <= 12'h179;
        src13 <= 12'hf44;
        src14 <= 12'h81f;
        src15 <= 12'he80;
        src16 <= 12'h8b;
        src17 <= 12'hc91;
        src18 <= 12'h145;
        src19 <= 12'he5b;
        src20 <= 12'h7a8;
        src21 <= 12'hdd1;
        src22 <= 12'h9f9;
        src23 <= 12'h936;
        src24 <= 12'he13;
        src25 <= 12'h896;
        src26 <= 12'ha62;
        src27 <= 12'h36f;
        src28 <= 12'h1c1;
        src29 <= 12'h3d5;
        src30 <= 12'hf5a;
        src31 <= 12'h614;
        src32 <= 12'hb89;
        src33 <= 12'hb35;
        src34 <= 12'h1f0;
        src35 <= 12'h519;
        src36 <= 12'h13f;
        src37 <= 12'hf67;
        src38 <= 12'h43c;
        src39 <= 12'h84b;
        src40 <= 12'h2ff;
        src41 <= 12'h1f5;
        src42 <= 12'h6cc;
        src43 <= 12'h711;
        src44 <= 12'hdb0;
        src45 <= 12'h7f6;
        src46 <= 12'h905;
        src47 <= 12'h70;
        src48 <= 12'hc0d;
        src49 <= 12'hf8b;
        src50 <= 12'hdb9;
        src51 <= 12'h276;
        src52 <= 12'ha9;
        src53 <= 12'h3b8;
        src54 <= 12'h6cd;
        src55 <= 12'hc46;
        src56 <= 12'he0e;
        src57 <= 12'h1c7;
        src58 <= 12'h8f;
        src59 <= 12'h876;
        src60 <= 12'h5ea;
        src61 <= 12'h5de;
        src62 <= 12'h361;
        src63 <= 12'h620;
        src64 <= 12'hf5f;
        src65 <= 12'h47b;
        src66 <= 12'h296;
        src67 <= 12'h7ff;
        src68 <= 12'hc6;
        src69 <= 12'hc3e;
        src70 <= 12'h465;
        src71 <= 12'h573;
        src72 <= 12'h205;
        src73 <= 12'h9a6;
        src74 <= 12'h522;
        src75 <= 12'h13;
        src76 <= 12'h807;
        src77 <= 12'h419;
        src78 <= 12'h6ea;
        src79 <= 12'h6c9;
        src80 <= 12'h9ce;
        src81 <= 12'hd99;
        src82 <= 12'hd0e;
        src83 <= 12'h51d;
        src84 <= 12'h5a5;
        src85 <= 12'h19f;
        src86 <= 12'h3c5;
        src87 <= 12'h915;
        src88 <= 12'hd18;
        src89 <= 12'he9f;
        src90 <= 12'h80c;
        src91 <= 12'h205;
        src92 <= 12'hcc7;
        src93 <= 12'h3;
        src94 <= 12'he81;
        src95 <= 12'h885;
        src96 <= 12'h2a9;
        src97 <= 12'h360;
        src98 <= 12'hd13;
        src99 <= 12'hfda;
        src100 <= 12'hdf0;
        src101 <= 12'h83b;
        src102 <= 12'haf6;
        src103 <= 12'hf18;
        src104 <= 12'h5a8;
        src105 <= 12'hf6d;
        src106 <= 12'hceb;
        src107 <= 12'h896;
        src108 <= 12'h20;
        src109 <= 12'heae;
        src110 <= 12'ha6b;
        src111 <= 12'h122;
        src112 <= 12'hc02;
        src113 <= 12'h401;
        src114 <= 12'hb67;
        src115 <= 12'h18c;
        src116 <= 12'h963;
        src117 <= 12'h157;
        src118 <= 12'hbcc;
        src119 <= 12'hc27;
        src120 <= 12'h1f2;
        src121 <= 12'h75b;
        src122 <= 12'h3f2;
        src123 <= 12'h3f2;
        src124 <= 12'h957;
        src125 <= 12'hbad;
        src126 <= 12'h6da;
        src127 <= 12'h849;
        src128 <= 12'h2b7;
        src129 <= 12'hdc9;
        src130 <= 12'h7c6;
        src131 <= 12'h9fa;
        src132 <= 12'hc0e;
        src133 <= 12'hfe2;
        src134 <= 12'h6a3;
        src135 <= 12'h7f0;
        src136 <= 12'hf2d;
        src137 <= 12'h707;
        src138 <= 12'h962;
        src139 <= 12'h8e6;
        src140 <= 12'h4b3;
        src141 <= 12'hd62;
        src142 <= 12'hda3;
        src143 <= 12'hb3;
        src144 <= 12'h8da;
        src145 <= 12'h909;
        src146 <= 12'h69a;
        src147 <= 12'h19d;
        src148 <= 12'hdd7;
        src149 <= 12'he12;
        src150 <= 12'hc29;
        src151 <= 12'h14d;
        src152 <= 12'h98a;
        src153 <= 12'hc66;
        src154 <= 12'h1bf;
        src155 <= 12'hed5;
        src156 <= 12'he2d;
        src157 <= 12'h886;
        src158 <= 12'hc;
        src159 <= 12'h9aa;
        src160 <= 12'h77f;
        src161 <= 12'h3d4;
        exp <= 20'h51497;
        #1
        src0 <= 12'h1ef;
        src1 <= 12'h5a5;
        src2 <= 12'h70a;
        src3 <= 12'h134;
        src4 <= 12'h557;
        src5 <= 12'h47e;
        src6 <= 12'h98e;
        src7 <= 12'h5b1;
        src8 <= 12'ha38;
        src9 <= 12'h2bc;
        src10 <= 12'h1a4;
        src11 <= 12'he37;
        src12 <= 12'he4b;
        src13 <= 12'hf;
        src14 <= 12'h2f;
        src15 <= 12'hd2d;
        src16 <= 12'hb25;
        src17 <= 12'h789;
        src18 <= 12'h6f2;
        src19 <= 12'h1cb;
        src20 <= 12'hfc0;
        src21 <= 12'hc1f;
        src22 <= 12'h5ff;
        src23 <= 12'h5da;
        src24 <= 12'h870;
        src25 <= 12'h7ca;
        src26 <= 12'hc8d;
        src27 <= 12'h79d;
        src28 <= 12'h9eb;
        src29 <= 12'h1c0;
        src30 <= 12'h35d;
        src31 <= 12'h4e2;
        src32 <= 12'h530;
        src33 <= 12'hdfa;
        src34 <= 12'hf67;
        src35 <= 12'hb98;
        src36 <= 12'he;
        src37 <= 12'h65c;
        src38 <= 12'h64f;
        src39 <= 12'h695;
        src40 <= 12'hdb0;
        src41 <= 12'h5ec;
        src42 <= 12'he6c;
        src43 <= 12'hcd5;
        src44 <= 12'h44b;
        src45 <= 12'h6d0;
        src46 <= 12'hb23;
        src47 <= 12'h1f1;
        src48 <= 12'h3fd;
        src49 <= 12'hede;
        src50 <= 12'h23d;
        src51 <= 12'he26;
        src52 <= 12'h855;
        src53 <= 12'hf9f;
        src54 <= 12'h8c3;
        src55 <= 12'h192;
        src56 <= 12'hf3b;
        src57 <= 12'h81;
        src58 <= 12'h85;
        src59 <= 12'h526;
        src60 <= 12'h9a6;
        src61 <= 12'h2e7;
        src62 <= 12'he45;
        src63 <= 12'hcc3;
        src64 <= 12'hfd9;
        src65 <= 12'h373;
        src66 <= 12'h116;
        src67 <= 12'h7c;
        src68 <= 12'h467;
        src69 <= 12'hce2;
        src70 <= 12'hbf6;
        src71 <= 12'hf86;
        src72 <= 12'hd37;
        src73 <= 12'h96e;
        src74 <= 12'hf;
        src75 <= 12'hfc8;
        src76 <= 12'h72b;
        src77 <= 12'ha03;
        src78 <= 12'h3d5;
        src79 <= 12'h37b;
        src80 <= 12'hd1;
        src81 <= 12'hac7;
        src82 <= 12'hb12;
        src83 <= 12'hefd;
        src84 <= 12'he0b;
        src85 <= 12'h92d;
        src86 <= 12'h1d8;
        src87 <= 12'h90;
        src88 <= 12'h3d1;
        src89 <= 12'hd8d;
        src90 <= 12'h1dc;
        src91 <= 12'h3b8;
        src92 <= 12'h663;
        src93 <= 12'h9ba;
        src94 <= 12'heef;
        src95 <= 12'h5a;
        src96 <= 12'h715;
        src97 <= 12'h250;
        src98 <= 12'h30;
        src99 <= 12'hf77;
        src100 <= 12'hedb;
        src101 <= 12'hba5;
        src102 <= 12'h2bd;
        src103 <= 12'he12;
        src104 <= 12'hefd;
        src105 <= 12'h636;
        src106 <= 12'h90;
        src107 <= 12'haaa;
        src108 <= 12'h7d2;
        src109 <= 12'h927;
        src110 <= 12'h66b;
        src111 <= 12'h6a3;
        src112 <= 12'h718;
        src113 <= 12'h98a;
        src114 <= 12'h5d8;
        src115 <= 12'hc87;
        src116 <= 12'h5a5;
        src117 <= 12'hb2c;
        src118 <= 12'h945;
        src119 <= 12'hf63;
        src120 <= 12'hf93;
        src121 <= 12'hac6;
        src122 <= 12'h53a;
        src123 <= 12'hd9c;
        src124 <= 12'hf09;
        src125 <= 12'h93d;
        src126 <= 12'h29;
        src127 <= 12'h341;
        src128 <= 12'h390;
        src129 <= 12'h5d7;
        src130 <= 12'hce3;
        src131 <= 12'h726;
        src132 <= 12'h680;
        src133 <= 12'h810;
        src134 <= 12'h992;
        src135 <= 12'h144;
        src136 <= 12'h2ae;
        src137 <= 12'h49a;
        src138 <= 12'h92a;
        src139 <= 12'hd2;
        src140 <= 12'h13c;
        src141 <= 12'he23;
        src142 <= 12'h505;
        src143 <= 12'h113;
        src144 <= 12'h430;
        src145 <= 12'h437;
        src146 <= 12'h489;
        src147 <= 12'hc4a;
        src148 <= 12'heec;
        src149 <= 12'hb2;
        src150 <= 12'hc43;
        src151 <= 12'h101;
        src152 <= 12'h4ab;
        src153 <= 12'h575;
        src154 <= 12'h499;
        src155 <= 12'hcbf;
        src156 <= 12'h63c;
        src157 <= 12'h842;
        src158 <= 12'h560;
        src159 <= 12'h1ae;
        src160 <= 12'hf5d;
        src161 <= 12'hf08;
        exp <= 20'h4d95c;
        #1
        src0 <= 12'hbce;
        src1 <= 12'h440;
        src2 <= 12'hc45;
        src3 <= 12'hd0b;
        src4 <= 12'h4a8;
        src5 <= 12'hd30;
        src6 <= 12'h667;
        src7 <= 12'h3f8;
        src8 <= 12'h4c9;
        src9 <= 12'hcb5;
        src10 <= 12'hb29;
        src11 <= 12'h2a5;
        src12 <= 12'hc88;
        src13 <= 12'hcff;
        src14 <= 12'h29c;
        src15 <= 12'h24e;
        src16 <= 12'h5b2;
        src17 <= 12'hfd8;
        src18 <= 12'h4c7;
        src19 <= 12'hd8d;
        src20 <= 12'h791;
        src21 <= 12'h592;
        src22 <= 12'h3d6;
        src23 <= 12'h852;
        src24 <= 12'h6f7;
        src25 <= 12'h22d;
        src26 <= 12'hc73;
        src27 <= 12'h301;
        src28 <= 12'hfd6;
        src29 <= 12'h36c;
        src30 <= 12'h65d;
        src31 <= 12'h2c2;
        src32 <= 12'h374;
        src33 <= 12'hd8;
        src34 <= 12'he2;
        src35 <= 12'hd4;
        src36 <= 12'h591;
        src37 <= 12'hcb8;
        src38 <= 12'ha06;
        src39 <= 12'h9d8;
        src40 <= 12'h562;
        src41 <= 12'h128;
        src42 <= 12'hf55;
        src43 <= 12'h95c;
        src44 <= 12'h7af;
        src45 <= 12'h3df;
        src46 <= 12'hb23;
        src47 <= 12'h68f;
        src48 <= 12'hc19;
        src49 <= 12'h828;
        src50 <= 12'h95d;
        src51 <= 12'hfb6;
        src52 <= 12'hbfb;
        src53 <= 12'h503;
        src54 <= 12'h9d0;
        src55 <= 12'h732;
        src56 <= 12'hb1c;
        src57 <= 12'h903;
        src58 <= 12'h709;
        src59 <= 12'h5b;
        src60 <= 12'hf45;
        src61 <= 12'h4dc;
        src62 <= 12'h19f;
        src63 <= 12'hd9c;
        src64 <= 12'he1b;
        src65 <= 12'h968;
        src66 <= 12'hed4;
        src67 <= 12'h2a2;
        src68 <= 12'h3c2;
        src69 <= 12'hbfb;
        src70 <= 12'h4c;
        src71 <= 12'h606;
        src72 <= 12'hdf5;
        src73 <= 12'h74c;
        src74 <= 12'hff9;
        src75 <= 12'ha;
        src76 <= 12'h9d1;
        src77 <= 12'h411;
        src78 <= 12'h2f2;
        src79 <= 12'h310;
        src80 <= 12'h9a3;
        src81 <= 12'haac;
        src82 <= 12'hc85;
        src83 <= 12'h16b;
        src84 <= 12'h815;
        src85 <= 12'h5cb;
        src86 <= 12'h6b8;
        src87 <= 12'h63d;
        src88 <= 12'h59c;
        src89 <= 12'h376;
        src90 <= 12'h96a;
        src91 <= 12'h8c;
        src92 <= 12'hb0b;
        src93 <= 12'h186;
        src94 <= 12'ha00;
        src95 <= 12'h51a;
        src96 <= 12'h642;
        src97 <= 12'hb6d;
        src98 <= 12'h1c7;
        src99 <= 12'ha78;
        src100 <= 12'hc93;
        src101 <= 12'h1f0;
        src102 <= 12'h64d;
        src103 <= 12'hce1;
        src104 <= 12'h6a9;
        src105 <= 12'h3fe;
        src106 <= 12'hbd1;
        src107 <= 12'h9ca;
        src108 <= 12'h28;
        src109 <= 12'h909;
        src110 <= 12'hc3f;
        src111 <= 12'h17f;
        src112 <= 12'h606;
        src113 <= 12'hc26;
        src114 <= 12'ha3d;
        src115 <= 12'h69d;
        src116 <= 12'hac2;
        src117 <= 12'h54c;
        src118 <= 12'h67c;
        src119 <= 12'he6e;
        src120 <= 12'h550;
        src121 <= 12'hbb3;
        src122 <= 12'h83c;
        src123 <= 12'hb1d;
        src124 <= 12'h7af;
        src125 <= 12'h414;
        src126 <= 12'h310;
        src127 <= 12'hff;
        src128 <= 12'h8b2;
        src129 <= 12'h2a7;
        src130 <= 12'hde2;
        src131 <= 12'hf99;
        src132 <= 12'hf25;
        src133 <= 12'hc39;
        src134 <= 12'h42e;
        src135 <= 12'h77b;
        src136 <= 12'ha87;
        src137 <= 12'he73;
        src138 <= 12'h243;
        src139 <= 12'hf6e;
        src140 <= 12'h1c8;
        src141 <= 12'h225;
        src142 <= 12'hcd1;
        src143 <= 12'hf0;
        src144 <= 12'hf1a;
        src145 <= 12'h8b7;
        src146 <= 12'h1ab;
        src147 <= 12'hd95;
        src148 <= 12'h6f0;
        src149 <= 12'h792;
        src150 <= 12'h38;
        src151 <= 12'he52;
        src152 <= 12'h715;
        src153 <= 12'hbd8;
        src154 <= 12'h62c;
        src155 <= 12'h837;
        src156 <= 12'h22d;
        src157 <= 12'hec2;
        src158 <= 12'h266;
        src159 <= 12'h5db;
        src160 <= 12'hdf8;
        src161 <= 12'h6cb;
        exp <= 20'h4e6d2;
        #1
        src0 <= 12'h5c8;
        src1 <= 12'hde3;
        src2 <= 12'hc39;
        src3 <= 12'ha9d;
        src4 <= 12'h511;
        src5 <= 12'hbc6;
        src6 <= 12'h752;
        src7 <= 12'hdb2;
        src8 <= 12'h4d4;
        src9 <= 12'h22f;
        src10 <= 12'h1b9;
        src11 <= 12'hf2f;
        src12 <= 12'h34b;
        src13 <= 12'he6f;
        src14 <= 12'he18;
        src15 <= 12'hb5d;
        src16 <= 12'haea;
        src17 <= 12'hb39;
        src18 <= 12'h74a;
        src19 <= 12'h301;
        src20 <= 12'h1d;
        src21 <= 12'haef;
        src22 <= 12'h8a6;
        src23 <= 12'h706;
        src24 <= 12'h240;
        src25 <= 12'h90e;
        src26 <= 12'heff;
        src27 <= 12'hfae;
        src28 <= 12'h48c;
        src29 <= 12'h958;
        src30 <= 12'hcaf;
        src31 <= 12'h263;
        src32 <= 12'hac;
        src33 <= 12'h425;
        src34 <= 12'ha21;
        src35 <= 12'h492;
        src36 <= 12'hfa3;
        src37 <= 12'h931;
        src38 <= 12'h70c;
        src39 <= 12'h423;
        src40 <= 12'h142;
        src41 <= 12'h7ec;
        src42 <= 12'h88;
        src43 <= 12'hb53;
        src44 <= 12'he8;
        src45 <= 12'ha65;
        src46 <= 12'hb71;
        src47 <= 12'h1d2;
        src48 <= 12'he47;
        src49 <= 12'h286;
        src50 <= 12'h4c3;
        src51 <= 12'h938;
        src52 <= 12'h76f;
        src53 <= 12'h6fa;
        src54 <= 12'h8f9;
        src55 <= 12'hd0e;
        src56 <= 12'h7e9;
        src57 <= 12'h1c0;
        src58 <= 12'heaf;
        src59 <= 12'h230;
        src60 <= 12'h859;
        src61 <= 12'h63e;
        src62 <= 12'h9bb;
        src63 <= 12'h98e;
        src64 <= 12'h525;
        src65 <= 12'h113;
        src66 <= 12'he86;
        src67 <= 12'h89a;
        src68 <= 12'hdef;
        src69 <= 12'h4c3;
        src70 <= 12'h3eb;
        src71 <= 12'h16b;
        src72 <= 12'h966;
        src73 <= 12'h793;
        src74 <= 12'hdd9;
        src75 <= 12'h7fa;
        src76 <= 12'h381;
        src77 <= 12'h851;
        src78 <= 12'h9f2;
        src79 <= 12'hd78;
        src80 <= 12'h9d2;
        src81 <= 12'h14f;
        src82 <= 12'hcf8;
        src83 <= 12'hb0f;
        src84 <= 12'h29b;
        src85 <= 12'h56;
        src86 <= 12'h9bf;
        src87 <= 12'hde6;
        src88 <= 12'h34d;
        src89 <= 12'h3c;
        src90 <= 12'he53;
        src91 <= 12'h2ef;
        src92 <= 12'h9ec;
        src93 <= 12'h510;
        src94 <= 12'h370;
        src95 <= 12'hc46;
        src96 <= 12'h88e;
        src97 <= 12'h2b5;
        src98 <= 12'h437;
        src99 <= 12'he6c;
        src100 <= 12'hc14;
        src101 <= 12'h71d;
        src102 <= 12'ha50;
        src103 <= 12'heca;
        src104 <= 12'hc27;
        src105 <= 12'h9e2;
        src106 <= 12'hb10;
        src107 <= 12'hed0;
        src108 <= 12'hfba;
        src109 <= 12'he5b;
        src110 <= 12'h2dd;
        src111 <= 12'h2d;
        src112 <= 12'h74e;
        src113 <= 12'h54b;
        src114 <= 12'h252;
        src115 <= 12'h37b;
        src116 <= 12'hbc3;
        src117 <= 12'hf75;
        src118 <= 12'h186;
        src119 <= 12'h8a1;
        src120 <= 12'hb3b;
        src121 <= 12'h341;
        src122 <= 12'h431;
        src123 <= 12'ha77;
        src124 <= 12'h3c1;
        src125 <= 12'ha92;
        src126 <= 12'h621;
        src127 <= 12'he46;
        src128 <= 12'h37c;
        src129 <= 12'hef8;
        src130 <= 12'hc6;
        src131 <= 12'h8a5;
        src132 <= 12'h69a;
        src133 <= 12'h646;
        src134 <= 12'hf9a;
        src135 <= 12'h4e0;
        src136 <= 12'hbd3;
        src137 <= 12'h520;
        src138 <= 12'hd7a;
        src139 <= 12'hb91;
        src140 <= 12'h8d4;
        src141 <= 12'hae8;
        src142 <= 12'h2be;
        src143 <= 12'hfd5;
        src144 <= 12'hdf1;
        src145 <= 12'h945;
        src146 <= 12'ha94;
        src147 <= 12'h40;
        src148 <= 12'hae;
        src149 <= 12'h3bb;
        src150 <= 12'hecb;
        src151 <= 12'h381;
        src152 <= 12'hdb8;
        src153 <= 12'h6df;
        src154 <= 12'h5d7;
        src155 <= 12'hf2d;
        src156 <= 12'h24e;
        src157 <= 12'h824;
        src158 <= 12'h9d3;
        src159 <= 12'h620;
        src160 <= 12'h96f;
        src161 <= 12'hd7e;
        exp <= 20'h51efe;
        #1
        src0 <= 12'h343;
        src1 <= 12'h71a;
        src2 <= 12'hb3b;
        src3 <= 12'hda2;
        src4 <= 12'hb6a;
        src5 <= 12'h6ac;
        src6 <= 12'h497;
        src7 <= 12'h21c;
        src8 <= 12'he98;
        src9 <= 12'hb2;
        src10 <= 12'hca6;
        src11 <= 12'h824;
        src12 <= 12'h984;
        src13 <= 12'h10e;
        src14 <= 12'h463;
        src15 <= 12'hdff;
        src16 <= 12'h2b1;
        src17 <= 12'h40;
        src18 <= 12'h6e2;
        src19 <= 12'h2c9;
        src20 <= 12'h345;
        src21 <= 12'hdc5;
        src22 <= 12'h3fe;
        src23 <= 12'hb6d;
        src24 <= 12'hf0e;
        src25 <= 12'h96a;
        src26 <= 12'hb51;
        src27 <= 12'h8b2;
        src28 <= 12'h5a0;
        src29 <= 12'h472;
        src30 <= 12'hfe4;
        src31 <= 12'he15;
        src32 <= 12'hf4;
        src33 <= 12'h6bf;
        src34 <= 12'ha3f;
        src35 <= 12'h2e;
        src36 <= 12'hb23;
        src37 <= 12'h758;
        src38 <= 12'hc84;
        src39 <= 12'hdc6;
        src40 <= 12'h9d8;
        src41 <= 12'hcd8;
        src42 <= 12'h338;
        src43 <= 12'h53b;
        src44 <= 12'hd03;
        src45 <= 12'h6be;
        src46 <= 12'hd12;
        src47 <= 12'h8d1;
        src48 <= 12'hada;
        src49 <= 12'hfc7;
        src50 <= 12'h329;
        src51 <= 12'hfb2;
        src52 <= 12'h2dc;
        src53 <= 12'h87f;
        src54 <= 12'hc4c;
        src55 <= 12'hf4f;
        src56 <= 12'h1ce;
        src57 <= 12'h62e;
        src58 <= 12'h172;
        src59 <= 12'h9e0;
        src60 <= 12'h9ee;
        src61 <= 12'h841;
        src62 <= 12'h43;
        src63 <= 12'hfb5;
        src64 <= 12'h2d1;
        src65 <= 12'h5f8;
        src66 <= 12'hbec;
        src67 <= 12'h3f1;
        src68 <= 12'h28b;
        src69 <= 12'hb36;
        src70 <= 12'h878;
        src71 <= 12'hae2;
        src72 <= 12'hfac;
        src73 <= 12'h9b;
        src74 <= 12'h82f;
        src75 <= 12'h301;
        src76 <= 12'hf3e;
        src77 <= 12'h5a4;
        src78 <= 12'h524;
        src79 <= 12'heb8;
        src80 <= 12'h44e;
        src81 <= 12'hee5;
        src82 <= 12'he2a;
        src83 <= 12'h9b2;
        src84 <= 12'he37;
        src85 <= 12'he2a;
        src86 <= 12'h6ed;
        src87 <= 12'ha95;
        src88 <= 12'hf36;
        src89 <= 12'h52e;
        src90 <= 12'hf55;
        src91 <= 12'h276;
        src92 <= 12'h935;
        src93 <= 12'hdcd;
        src94 <= 12'h707;
        src95 <= 12'h174;
        src96 <= 12'h63a;
        src97 <= 12'h61d;
        src98 <= 12'hcb2;
        src99 <= 12'h829;
        src100 <= 12'h152;
        src101 <= 12'h8ec;
        src102 <= 12'he63;
        src103 <= 12'h440;
        src104 <= 12'h5b4;
        src105 <= 12'h3e0;
        src106 <= 12'h76b;
        src107 <= 12'h2a;
        src108 <= 12'hd83;
        src109 <= 12'h313;
        src110 <= 12'he25;
        src111 <= 12'h203;
        src112 <= 12'hbf0;
        src113 <= 12'hfff;
        src114 <= 12'h32;
        src115 <= 12'he40;
        src116 <= 12'h793;
        src117 <= 12'ha2c;
        src118 <= 12'h955;
        src119 <= 12'h8e4;
        src120 <= 12'he8e;
        src121 <= 12'h104;
        src122 <= 12'hb93;
        src123 <= 12'habf;
        src124 <= 12'h225;
        src125 <= 12'h18f;
        src126 <= 12'h93e;
        src127 <= 12'h264;
        src128 <= 12'h5ec;
        src129 <= 12'h348;
        src130 <= 12'h293;
        src131 <= 12'hf72;
        src132 <= 12'h947;
        src133 <= 12'h682;
        src134 <= 12'hf68;
        src135 <= 12'h39a;
        src136 <= 12'h683;
        src137 <= 12'hf12;
        src138 <= 12'hd3f;
        src139 <= 12'h145;
        src140 <= 12'h90b;
        src141 <= 12'h617;
        src142 <= 12'h36f;
        src143 <= 12'h1cb;
        src144 <= 12'hc0e;
        src145 <= 12'h590;
        src146 <= 12'haf1;
        src147 <= 12'h5ae;
        src148 <= 12'hf2a;
        src149 <= 12'h262;
        src150 <= 12'hf98;
        src151 <= 12'h6c6;
        src152 <= 12'h8a8;
        src153 <= 12'h205;
        src154 <= 12'he53;
        src155 <= 12'he4f;
        src156 <= 12'h409;
        src157 <= 12'hc0e;
        src158 <= 12'h475;
        src159 <= 12'h146;
        src160 <= 12'h67f;
        src161 <= 12'hc3c;
        exp <= 20'h530d2;
        #1
        src0 <= 12'h97;
        src1 <= 12'h2a7;
        src2 <= 12'h71;
        src3 <= 12'hf76;
        src4 <= 12'h96a;
        src5 <= 12'hfb0;
        src6 <= 12'he75;
        src7 <= 12'h3ee;
        src8 <= 12'hfad;
        src9 <= 12'h864;
        src10 <= 12'h743;
        src11 <= 12'h436;
        src12 <= 12'h719;
        src13 <= 12'ha8f;
        src14 <= 12'h9fd;
        src15 <= 12'h74f;
        src16 <= 12'h987;
        src17 <= 12'hba1;
        src18 <= 12'h15;
        src19 <= 12'h3c0;
        src20 <= 12'h1cd;
        src21 <= 12'h91d;
        src22 <= 12'hfc1;
        src23 <= 12'hc86;
        src24 <= 12'hce1;
        src25 <= 12'h5e4;
        src26 <= 12'h959;
        src27 <= 12'hae0;
        src28 <= 12'h731;
        src29 <= 12'h38e;
        src30 <= 12'h33b;
        src31 <= 12'h3ef;
        src32 <= 12'h45b;
        src33 <= 12'h486;
        src34 <= 12'hd7e;
        src35 <= 12'ha09;
        src36 <= 12'h53e;
        src37 <= 12'h818;
        src38 <= 12'h538;
        src39 <= 12'h92a;
        src40 <= 12'h976;
        src41 <= 12'h2e2;
        src42 <= 12'h36;
        src43 <= 12'hd5c;
        src44 <= 12'h873;
        src45 <= 12'hae4;
        src46 <= 12'h21d;
        src47 <= 12'h219;
        src48 <= 12'hdff;
        src49 <= 12'h24a;
        src50 <= 12'h203;
        src51 <= 12'ha7f;
        src52 <= 12'h8c8;
        src53 <= 12'h39;
        src54 <= 12'hab;
        src55 <= 12'h4ee;
        src56 <= 12'h6aa;
        src57 <= 12'h39f;
        src58 <= 12'h0;
        src59 <= 12'h2b3;
        src60 <= 12'haac;
        src61 <= 12'h347;
        src62 <= 12'he94;
        src63 <= 12'he7a;
        src64 <= 12'h147;
        src65 <= 12'h1c7;
        src66 <= 12'h993;
        src67 <= 12'h3e2;
        src68 <= 12'h460;
        src69 <= 12'hb97;
        src70 <= 12'h33b;
        src71 <= 12'h7af;
        src72 <= 12'hf22;
        src73 <= 12'h287;
        src74 <= 12'hb2b;
        src75 <= 12'h793;
        src76 <= 12'h45f;
        src77 <= 12'h9f2;
        src78 <= 12'h3a6;
        src79 <= 12'hefc;
        src80 <= 12'hab4;
        src81 <= 12'h5ce;
        src82 <= 12'h92;
        src83 <= 12'h705;
        src84 <= 12'hb96;
        src85 <= 12'h79c;
        src86 <= 12'hfa8;
        src87 <= 12'hd00;
        src88 <= 12'h1a4;
        src89 <= 12'h970;
        src90 <= 12'h351;
        src91 <= 12'h553;
        src92 <= 12'h9ba;
        src93 <= 12'hdd7;
        src94 <= 12'h845;
        src95 <= 12'h927;
        src96 <= 12'h529;
        src97 <= 12'h6e5;
        src98 <= 12'h853;
        src99 <= 12'h5dc;
        src100 <= 12'haac;
        src101 <= 12'hbcc;
        src102 <= 12'haea;
        src103 <= 12'hce8;
        src104 <= 12'h9c4;
        src105 <= 12'h117;
        src106 <= 12'h588;
        src107 <= 12'hd9d;
        src108 <= 12'h0;
        src109 <= 12'h711;
        src110 <= 12'hace;
        src111 <= 12'hae9;
        src112 <= 12'h592;
        src113 <= 12'h3be;
        src114 <= 12'hf48;
        src115 <= 12'hddc;
        src116 <= 12'hd30;
        src117 <= 12'h446;
        src118 <= 12'hb5a;
        src119 <= 12'hc04;
        src120 <= 12'h739;
        src121 <= 12'h1ab;
        src122 <= 12'had8;
        src123 <= 12'hf7d;
        src124 <= 12'hd25;
        src125 <= 12'hbb4;
        src126 <= 12'h3de;
        src127 <= 12'he1b;
        src128 <= 12'h597;
        src129 <= 12'h1fa;
        src130 <= 12'h67f;
        src131 <= 12'he04;
        src132 <= 12'hd1f;
        src133 <= 12'hf29;
        src134 <= 12'h2b0;
        src135 <= 12'h7bf;
        src136 <= 12'h780;
        src137 <= 12'h490;
        src138 <= 12'h640;
        src139 <= 12'hed6;
        src140 <= 12'hc67;
        src141 <= 12'hd46;
        src142 <= 12'h82;
        src143 <= 12'h8d1;
        src144 <= 12'hf2d;
        src145 <= 12'hb4f;
        src146 <= 12'hf06;
        src147 <= 12'h197;
        src148 <= 12'h178;
        src149 <= 12'h179;
        src150 <= 12'h883;
        src151 <= 12'h166;
        src152 <= 12'hdb8;
        src153 <= 12'hd8e;
        src154 <= 12'h504;
        src155 <= 12'h224;
        src156 <= 12'hb8d;
        src157 <= 12'h44c;
        src158 <= 12'he4;
        src159 <= 12'h5cf;
        src160 <= 12'hb0a;
        src161 <= 12'h852;
        exp <= 20'h4f070;
        #1
        src0 <= 12'h17e;
        src1 <= 12'h71b;
        src2 <= 12'h1bc;
        src3 <= 12'h188;
        src4 <= 12'hb65;
        src5 <= 12'h83c;
        src6 <= 12'hecd;
        src7 <= 12'hea0;
        src8 <= 12'he63;
        src9 <= 12'h3e;
        src10 <= 12'h7b7;
        src11 <= 12'h2a9;
        src12 <= 12'h6cc;
        src13 <= 12'h3d4;
        src14 <= 12'h630;
        src15 <= 12'h997;
        src16 <= 12'hf10;
        src17 <= 12'hea8;
        src18 <= 12'had8;
        src19 <= 12'hbc;
        src20 <= 12'hc86;
        src21 <= 12'hbbc;
        src22 <= 12'h95a;
        src23 <= 12'h9ab;
        src24 <= 12'ha23;
        src25 <= 12'h77;
        src26 <= 12'h7fb;
        src27 <= 12'hfb9;
        src28 <= 12'h2f7;
        src29 <= 12'hdf;
        src30 <= 12'h70f;
        src31 <= 12'hd88;
        src32 <= 12'heb4;
        src33 <= 12'h65a;
        src34 <= 12'h66f;
        src35 <= 12'hcb0;
        src36 <= 12'haa0;
        src37 <= 12'hd1;
        src38 <= 12'h508;
        src39 <= 12'h64b;
        src40 <= 12'h11a;
        src41 <= 12'h315;
        src42 <= 12'ha7a;
        src43 <= 12'h9c1;
        src44 <= 12'h8cd;
        src45 <= 12'hac9;
        src46 <= 12'hfdb;
        src47 <= 12'h872;
        src48 <= 12'had6;
        src49 <= 12'hdf7;
        src50 <= 12'hb8c;
        src51 <= 12'hc67;
        src52 <= 12'h10f;
        src53 <= 12'h553;
        src54 <= 12'h233;
        src55 <= 12'h8c5;
        src56 <= 12'h98b;
        src57 <= 12'h616;
        src58 <= 12'h205;
        src59 <= 12'h1fa;
        src60 <= 12'h9d0;
        src61 <= 12'h410;
        src62 <= 12'h1e0;
        src63 <= 12'h31f;
        src64 <= 12'hc5c;
        src65 <= 12'h8e4;
        src66 <= 12'h57b;
        src67 <= 12'hd7e;
        src68 <= 12'he3e;
        src69 <= 12'h72;
        src70 <= 12'hc12;
        src71 <= 12'h6c7;
        src72 <= 12'h8f0;
        src73 <= 12'h83e;
        src74 <= 12'haeb;
        src75 <= 12'hac0;
        src76 <= 12'hc75;
        src77 <= 12'h684;
        src78 <= 12'h8d5;
        src79 <= 12'haa0;
        src80 <= 12'hfdc;
        src81 <= 12'h9e9;
        src82 <= 12'h407;
        src83 <= 12'h53a;
        src84 <= 12'hfc5;
        src85 <= 12'h244;
        src86 <= 12'haa1;
        src87 <= 12'hada;
        src88 <= 12'h674;
        src89 <= 12'haf8;
        src90 <= 12'h16d;
        src91 <= 12'hc17;
        src92 <= 12'h855;
        src93 <= 12'h534;
        src94 <= 12'h3cf;
        src95 <= 12'hcc3;
        src96 <= 12'h30a;
        src97 <= 12'h66e;
        src98 <= 12'hb4;
        src99 <= 12'h3c9;
        src100 <= 12'ha4;
        src101 <= 12'hf8f;
        src102 <= 12'he1e;
        src103 <= 12'h8b5;
        src104 <= 12'h119;
        src105 <= 12'h5fd;
        src106 <= 12'h35f;
        src107 <= 12'he;
        src108 <= 12'h6dc;
        src109 <= 12'h711;
        src110 <= 12'hbc7;
        src111 <= 12'ha06;
        src112 <= 12'h7b9;
        src113 <= 12'h2d3;
        src114 <= 12'h519;
        src115 <= 12'h8a;
        src116 <= 12'h7aa;
        src117 <= 12'h24f;
        src118 <= 12'h4d2;
        src119 <= 12'h9ef;
        src120 <= 12'he07;
        src121 <= 12'he04;
        src122 <= 12'h446;
        src123 <= 12'h2c2;
        src124 <= 12'hf3;
        src125 <= 12'h6c4;
        src126 <= 12'h6c9;
        src127 <= 12'h101;
        src128 <= 12'h21e;
        src129 <= 12'h620;
        src130 <= 12'h56f;
        src131 <= 12'hab8;
        src132 <= 12'hade;
        src133 <= 12'hf09;
        src134 <= 12'h1a4;
        src135 <= 12'h156;
        src136 <= 12'h866;
        src137 <= 12'h1f4;
        src138 <= 12'h46b;
        src139 <= 12'h36;
        src140 <= 12'he2f;
        src141 <= 12'h79d;
        src142 <= 12'h237;
        src143 <= 12'hd73;
        src144 <= 12'h284;
        src145 <= 12'he68;
        src146 <= 12'h874;
        src147 <= 12'h162;
        src148 <= 12'h8c8;
        src149 <= 12'hf14;
        src150 <= 12'h332;
        src151 <= 12'h432;
        src152 <= 12'hba9;
        src153 <= 12'had0;
        src154 <= 12'h144;
        src155 <= 12'h47d;
        src156 <= 12'h441;
        src157 <= 12'hd44;
        src158 <= 12'hb56;
        src159 <= 12'ha19;
        src160 <= 12'he5b;
        src161 <= 12'h876;
        exp <= 20'h4c683;
        #1
        src0 <= 12'h8e3;
        src1 <= 12'h69f;
        src2 <= 12'hd6e;
        src3 <= 12'hedc;
        src4 <= 12'h8e2;
        src5 <= 12'hbbc;
        src6 <= 12'hc05;
        src7 <= 12'ha76;
        src8 <= 12'h4c2;
        src9 <= 12'h961;
        src10 <= 12'h3e0;
        src11 <= 12'hbfc;
        src12 <= 12'hf87;
        src13 <= 12'hc4e;
        src14 <= 12'he62;
        src15 <= 12'h4f7;
        src16 <= 12'h978;
        src17 <= 12'h6a3;
        src18 <= 12'h693;
        src19 <= 12'h570;
        src20 <= 12'h376;
        src21 <= 12'ha5e;
        src22 <= 12'hae;
        src23 <= 12'h9bc;
        src24 <= 12'h722;
        src25 <= 12'h957;
        src26 <= 12'h1b1;
        src27 <= 12'h20e;
        src28 <= 12'ha5f;
        src29 <= 12'he76;
        src30 <= 12'hec1;
        src31 <= 12'h431;
        src32 <= 12'h797;
        src33 <= 12'h6fe;
        src34 <= 12'h5c2;
        src35 <= 12'h8e3;
        src36 <= 12'h674;
        src37 <= 12'h8c8;
        src38 <= 12'hfa8;
        src39 <= 12'h2d2;
        src40 <= 12'hf1a;
        src41 <= 12'h1d2;
        src42 <= 12'h8e;
        src43 <= 12'h5f4;
        src44 <= 12'hd88;
        src45 <= 12'h4c6;
        src46 <= 12'h213;
        src47 <= 12'he3;
        src48 <= 12'h4d4;
        src49 <= 12'h716;
        src50 <= 12'h2ff;
        src51 <= 12'h333;
        src52 <= 12'hbe;
        src53 <= 12'h100;
        src54 <= 12'hfa0;
        src55 <= 12'h569;
        src56 <= 12'hbc6;
        src57 <= 12'hf6b;
        src58 <= 12'h77f;
        src59 <= 12'h51;
        src60 <= 12'h5e7;
        src61 <= 12'h2c8;
        src62 <= 12'h3ef;
        src63 <= 12'hf88;
        src64 <= 12'h740;
        src65 <= 12'hf59;
        src66 <= 12'hbd2;
        src67 <= 12'h410;
        src68 <= 12'h123;
        src69 <= 12'h521;
        src70 <= 12'h389;
        src71 <= 12'h8ef;
        src72 <= 12'hf86;
        src73 <= 12'h8d2;
        src74 <= 12'h66c;
        src75 <= 12'h6e9;
        src76 <= 12'hbb8;
        src77 <= 12'h967;
        src78 <= 12'h613;
        src79 <= 12'hdaa;
        src80 <= 12'h390;
        src81 <= 12'h9c6;
        src82 <= 12'h7e2;
        src83 <= 12'ha30;
        src84 <= 12'hdac;
        src85 <= 12'hade;
        src86 <= 12'he1d;
        src87 <= 12'hbb4;
        src88 <= 12'hf5;
        src89 <= 12'hf4;
        src90 <= 12'h5bb;
        src91 <= 12'hb7d;
        src92 <= 12'h9bf;
        src93 <= 12'h50;
        src94 <= 12'h6c9;
        src95 <= 12'hf17;
        src96 <= 12'h70d;
        src97 <= 12'h5f8;
        src98 <= 12'hfcf;
        src99 <= 12'hfc4;
        src100 <= 12'h4c5;
        src101 <= 12'ha3a;
        src102 <= 12'haf1;
        src103 <= 12'h290;
        src104 <= 12'h3f8;
        src105 <= 12'hc0e;
        src106 <= 12'h545;
        src107 <= 12'h151;
        src108 <= 12'h222;
        src109 <= 12'hd51;
        src110 <= 12'ha4e;
        src111 <= 12'h80b;
        src112 <= 12'hf73;
        src113 <= 12'h714;
        src114 <= 12'h2ec;
        src115 <= 12'hbdb;
        src116 <= 12'hc08;
        src117 <= 12'h71e;
        src118 <= 12'h1eb;
        src119 <= 12'hf47;
        src120 <= 12'h7a5;
        src121 <= 12'hece;
        src122 <= 12'h8da;
        src123 <= 12'h508;
        src124 <= 12'hfbc;
        src125 <= 12'he52;
        src126 <= 12'h1db;
        src127 <= 12'hc12;
        src128 <= 12'he0c;
        src129 <= 12'hcd2;
        src130 <= 12'h98;
        src131 <= 12'h6ec;
        src132 <= 12'he7;
        src133 <= 12'hf91;
        src134 <= 12'hbab;
        src135 <= 12'hd43;
        src136 <= 12'hf56;
        src137 <= 12'h2bf;
        src138 <= 12'h14c;
        src139 <= 12'h5fd;
        src140 <= 12'h8bf;
        src141 <= 12'h15a;
        src142 <= 12'hb9f;
        src143 <= 12'he91;
        src144 <= 12'hb18;
        src145 <= 12'hc4d;
        src146 <= 12'hd6;
        src147 <= 12'hf61;
        src148 <= 12'h584;
        src149 <= 12'h4d7;
        src150 <= 12'h1d0;
        src151 <= 12'h626;
        src152 <= 12'h73f;
        src153 <= 12'h22;
        src154 <= 12'h6ff;
        src155 <= 12'h49c;
        src156 <= 12'h984;
        src157 <= 12'h971;
        src158 <= 12'h450;
        src159 <= 12'hfc4;
        src160 <= 12'h7f9;
        src161 <= 12'h244;
        exp <= 20'h51bc0;
        #1
        src0 <= 12'hdcb;
        src1 <= 12'hac9;
        src2 <= 12'hfc2;
        src3 <= 12'h4f9;
        src4 <= 12'h8b;
        src5 <= 12'hd38;
        src6 <= 12'h8a0;
        src7 <= 12'h880;
        src8 <= 12'h26e;
        src9 <= 12'h30d;
        src10 <= 12'hc5f;
        src11 <= 12'h35f;
        src12 <= 12'hbe;
        src13 <= 12'h67c;
        src14 <= 12'hd28;
        src15 <= 12'h266;
        src16 <= 12'h5a5;
        src17 <= 12'h2f2;
        src18 <= 12'hec9;
        src19 <= 12'h89c;
        src20 <= 12'ha5f;
        src21 <= 12'h36e;
        src22 <= 12'h267;
        src23 <= 12'h46e;
        src24 <= 12'hbf1;
        src25 <= 12'h7da;
        src26 <= 12'hdc4;
        src27 <= 12'h3ff;
        src28 <= 12'hb2f;
        src29 <= 12'hc7a;
        src30 <= 12'h29f;
        src31 <= 12'h5cd;
        src32 <= 12'hcaa;
        src33 <= 12'h59a;
        src34 <= 12'h202;
        src35 <= 12'h42d;
        src36 <= 12'hccc;
        src37 <= 12'he7b;
        src38 <= 12'h527;
        src39 <= 12'h864;
        src40 <= 12'h6b;
        src41 <= 12'hfdb;
        src42 <= 12'h63c;
        src43 <= 12'h48a;
        src44 <= 12'hf78;
        src45 <= 12'h9e2;
        src46 <= 12'h5cc;
        src47 <= 12'ha67;
        src48 <= 12'h5f0;
        src49 <= 12'h90e;
        src50 <= 12'h5c3;
        src51 <= 12'hf82;
        src52 <= 12'h933;
        src53 <= 12'h5dc;
        src54 <= 12'h9d;
        src55 <= 12'h402;
        src56 <= 12'h21d;
        src57 <= 12'hf38;
        src58 <= 12'hc02;
        src59 <= 12'h96b;
        src60 <= 12'hd7a;
        src61 <= 12'hf77;
        src62 <= 12'h9a0;
        src63 <= 12'hde9;
        src64 <= 12'hfbd;
        src65 <= 12'h52b;
        src66 <= 12'h404;
        src67 <= 12'h89a;
        src68 <= 12'he0f;
        src69 <= 12'haa3;
        src70 <= 12'h9d8;
        src71 <= 12'h2d;
        src72 <= 12'hcf2;
        src73 <= 12'he93;
        src74 <= 12'hecb;
        src75 <= 12'h68c;
        src76 <= 12'he4a;
        src77 <= 12'h19c;
        src78 <= 12'ha70;
        src79 <= 12'h147;
        src80 <= 12'hd28;
        src81 <= 12'h6d9;
        src82 <= 12'h97e;
        src83 <= 12'hca9;
        src84 <= 12'hefe;
        src85 <= 12'hd72;
        src86 <= 12'h729;
        src87 <= 12'h444;
        src88 <= 12'heb9;
        src89 <= 12'h838;
        src90 <= 12'h8a2;
        src91 <= 12'hbd4;
        src92 <= 12'ha6b;
        src93 <= 12'h872;
        src94 <= 12'h9f7;
        src95 <= 12'h821;
        src96 <= 12'h1e2;
        src97 <= 12'h4af;
        src98 <= 12'h22e;
        src99 <= 12'h64d;
        src100 <= 12'h734;
        src101 <= 12'h446;
        src102 <= 12'h537;
        src103 <= 12'h503;
        src104 <= 12'h765;
        src105 <= 12'hfd0;
        src106 <= 12'he90;
        src107 <= 12'hbde;
        src108 <= 12'ha74;
        src109 <= 12'h158;
        src110 <= 12'h32f;
        src111 <= 12'he0d;
        src112 <= 12'h319;
        src113 <= 12'h56e;
        src114 <= 12'hbfa;
        src115 <= 12'h5d3;
        src116 <= 12'h959;
        src117 <= 12'h330;
        src118 <= 12'h569;
        src119 <= 12'h9f1;
        src120 <= 12'h640;
        src121 <= 12'h278;
        src122 <= 12'h2f2;
        src123 <= 12'h792;
        src124 <= 12'hc07;
        src125 <= 12'h1b3;
        src126 <= 12'h58c;
        src127 <= 12'h9a6;
        src128 <= 12'h12b;
        src129 <= 12'hed9;
        src130 <= 12'hc63;
        src131 <= 12'h98d;
        src132 <= 12'h8c2;
        src133 <= 12'h19c;
        src134 <= 12'hf27;
        src135 <= 12'h72;
        src136 <= 12'h934;
        src137 <= 12'h2f2;
        src138 <= 12'he2a;
        src139 <= 12'haa2;
        src140 <= 12'h74f;
        src141 <= 12'hbf6;
        src142 <= 12'h55e;
        src143 <= 12'h479;
        src144 <= 12'he25;
        src145 <= 12'h839;
        src146 <= 12'hefb;
        src147 <= 12'hbc4;
        src148 <= 12'h9a1;
        src149 <= 12'hfd0;
        src150 <= 12'ha51;
        src151 <= 12'h138;
        src152 <= 12'h66;
        src153 <= 12'hb02;
        src154 <= 12'hc56;
        src155 <= 12'h75a;
        src156 <= 12'h837;
        src157 <= 12'hc4a;
        src158 <= 12'h34e;
        src159 <= 12'hfaa;
        src160 <= 12'h41a;
        src161 <= 12'h678;
        exp <= 20'h54193;
        #1
        src0 <= 12'hdb2;
        src1 <= 12'hb6c;
        src2 <= 12'h49b;
        src3 <= 12'hfe6;
        src4 <= 12'he8b;
        src5 <= 12'he;
        src6 <= 12'h2eb;
        src7 <= 12'h43f;
        src8 <= 12'hb78;
        src9 <= 12'h20b;
        src10 <= 12'h37c;
        src11 <= 12'hdc0;
        src12 <= 12'h500;
        src13 <= 12'h241;
        src14 <= 12'h1ce;
        src15 <= 12'h930;
        src16 <= 12'hdc2;
        src17 <= 12'h321;
        src18 <= 12'h13d;
        src19 <= 12'hd38;
        src20 <= 12'h40;
        src21 <= 12'he9d;
        src22 <= 12'h133;
        src23 <= 12'h997;
        src24 <= 12'h99a;
        src25 <= 12'heeb;
        src26 <= 12'hd7c;
        src27 <= 12'hd79;
        src28 <= 12'he1f;
        src29 <= 12'hc7b;
        src30 <= 12'hf2;
        src31 <= 12'hd47;
        src32 <= 12'h4da;
        src33 <= 12'h4d4;
        src34 <= 12'h440;
        src35 <= 12'h8b4;
        src36 <= 12'h4a8;
        src37 <= 12'h9a1;
        src38 <= 12'h2e5;
        src39 <= 12'h50f;
        src40 <= 12'h814;
        src41 <= 12'h563;
        src42 <= 12'h8df;
        src43 <= 12'he0c;
        src44 <= 12'h2ae;
        src45 <= 12'h83;
        src46 <= 12'hca5;
        src47 <= 12'hf79;
        src48 <= 12'hcd6;
        src49 <= 12'hea4;
        src50 <= 12'h618;
        src51 <= 12'hc27;
        src52 <= 12'he37;
        src53 <= 12'h832;
        src54 <= 12'h709;
        src55 <= 12'h13f;
        src56 <= 12'h55b;
        src57 <= 12'hb7a;
        src58 <= 12'ha1a;
        src59 <= 12'h32d;
        src60 <= 12'hc5e;
        src61 <= 12'h455;
        src62 <= 12'h5f7;
        src63 <= 12'h444;
        src64 <= 12'h504;
        src65 <= 12'hb06;
        src66 <= 12'h70b;
        src67 <= 12'hbf3;
        src68 <= 12'h687;
        src69 <= 12'ha67;
        src70 <= 12'hf05;
        src71 <= 12'hea4;
        src72 <= 12'h7f8;
        src73 <= 12'hd0a;
        src74 <= 12'hb65;
        src75 <= 12'hef1;
        src76 <= 12'ha60;
        src77 <= 12'hdaa;
        src78 <= 12'h203;
        src79 <= 12'h98a;
        src80 <= 12'h9fd;
        src81 <= 12'hfa1;
        src82 <= 12'ha43;
        src83 <= 12'hf4;
        src84 <= 12'he76;
        src85 <= 12'hea;
        src86 <= 12'h77b;
        src87 <= 12'he91;
        src88 <= 12'ha04;
        src89 <= 12'h75b;
        src90 <= 12'haf0;
        src91 <= 12'h950;
        src92 <= 12'h538;
        src93 <= 12'hd38;
        src94 <= 12'h642;
        src95 <= 12'h496;
        src96 <= 12'ha23;
        src97 <= 12'hf12;
        src98 <= 12'h845;
        src99 <= 12'hce1;
        src100 <= 12'h156;
        src101 <= 12'h540;
        src102 <= 12'h4ab;
        src103 <= 12'hec;
        src104 <= 12'hd4;
        src105 <= 12'hd2;
        src106 <= 12'h17a;
        src107 <= 12'hf58;
        src108 <= 12'hf1d;
        src109 <= 12'ha82;
        src110 <= 12'h17a;
        src111 <= 12'h433;
        src112 <= 12'h7bd;
        src113 <= 12'hec3;
        src114 <= 12'h64b;
        src115 <= 12'hb93;
        src116 <= 12'h93e;
        src117 <= 12'hdfc;
        src118 <= 12'h701;
        src119 <= 12'hcd6;
        src120 <= 12'h7bb;
        src121 <= 12'hc36;
        src122 <= 12'h328;
        src123 <= 12'h23b;
        src124 <= 12'he90;
        src125 <= 12'h4df;
        src126 <= 12'h4cb;
        src127 <= 12'hed8;
        src128 <= 12'h29a;
        src129 <= 12'h6ba;
        src130 <= 12'h8f7;
        src131 <= 12'hdd8;
        src132 <= 12'hcf1;
        src133 <= 12'h265;
        src134 <= 12'hce2;
        src135 <= 12'h269;
        src136 <= 12'h613;
        src137 <= 12'hf86;
        src138 <= 12'hd76;
        src139 <= 12'h545;
        src140 <= 12'h63b;
        src141 <= 12'he25;
        src142 <= 12'h619;
        src143 <= 12'heb8;
        src144 <= 12'he4d;
        src145 <= 12'hb8e;
        src146 <= 12'hf8f;
        src147 <= 12'h332;
        src148 <= 12'h7c8;
        src149 <= 12'h6d8;
        src150 <= 12'h210;
        src151 <= 12'he31;
        src152 <= 12'hc1d;
        src153 <= 12'h8c3;
        src154 <= 12'hd3a;
        src155 <= 12'hafe;
        src156 <= 12'hdd;
        src157 <= 12'h1c7;
        src158 <= 12'h5d0;
        src159 <= 12'hfe0;
        src160 <= 12'hfad;
        src161 <= 12'h667;
        exp <= 20'h568cd;
        #1
        src0 <= 12'h385;
        src1 <= 12'hd44;
        src2 <= 12'he2d;
        src3 <= 12'h178;
        src4 <= 12'h657;
        src5 <= 12'h1dd;
        src6 <= 12'hbdb;
        src7 <= 12'h350;
        src8 <= 12'h9ad;
        src9 <= 12'hd14;
        src10 <= 12'hd2d;
        src11 <= 12'hd52;
        src12 <= 12'h7a7;
        src13 <= 12'h99;
        src14 <= 12'h8ef;
        src15 <= 12'h34b;
        src16 <= 12'hb68;
        src17 <= 12'h2e4;
        src18 <= 12'h6d3;
        src19 <= 12'hceb;
        src20 <= 12'hb40;
        src21 <= 12'he29;
        src22 <= 12'he14;
        src23 <= 12'h7e7;
        src24 <= 12'h53f;
        src25 <= 12'h74;
        src26 <= 12'h8c3;
        src27 <= 12'h916;
        src28 <= 12'h95d;
        src29 <= 12'ha84;
        src30 <= 12'hbda;
        src31 <= 12'hda7;
        src32 <= 12'h274;
        src33 <= 12'hb88;
        src34 <= 12'hc8f;
        src35 <= 12'hf9f;
        src36 <= 12'hc4e;
        src37 <= 12'he1d;
        src38 <= 12'h8a;
        src39 <= 12'hb84;
        src40 <= 12'h76;
        src41 <= 12'h476;
        src42 <= 12'h422;
        src43 <= 12'h640;
        src44 <= 12'h84b;
        src45 <= 12'h3bf;
        src46 <= 12'hfb9;
        src47 <= 12'h5d2;
        src48 <= 12'h64a;
        src49 <= 12'hebc;
        src50 <= 12'h18d;
        src51 <= 12'h6c3;
        src52 <= 12'habe;
        src53 <= 12'h820;
        src54 <= 12'hc81;
        src55 <= 12'h6d9;
        src56 <= 12'h9f5;
        src57 <= 12'hcea;
        src58 <= 12'h41e;
        src59 <= 12'h5bb;
        src60 <= 12'h4f0;
        src61 <= 12'h7d5;
        src62 <= 12'h306;
        src63 <= 12'h5ab;
        src64 <= 12'hd45;
        src65 <= 12'h21d;
        src66 <= 12'hd7;
        src67 <= 12'h964;
        src68 <= 12'h83e;
        src69 <= 12'h81d;
        src70 <= 12'h3d5;
        src71 <= 12'h705;
        src72 <= 12'hc1e;
        src73 <= 12'hc40;
        src74 <= 12'h10f;
        src75 <= 12'h2f0;
        src76 <= 12'h78f;
        src77 <= 12'ha33;
        src78 <= 12'h8db;
        src79 <= 12'hb72;
        src80 <= 12'h2e9;
        src81 <= 12'h897;
        src82 <= 12'h148;
        src83 <= 12'hd95;
        src84 <= 12'h9a5;
        src85 <= 12'h4f4;
        src86 <= 12'h54f;
        src87 <= 12'h7e0;
        src88 <= 12'h862;
        src89 <= 12'hd22;
        src90 <= 12'hb0e;
        src91 <= 12'h6ba;
        src92 <= 12'h227;
        src93 <= 12'h2c4;
        src94 <= 12'h8e;
        src95 <= 12'hd4d;
        src96 <= 12'h52;
        src97 <= 12'h80d;
        src98 <= 12'hfd;
        src99 <= 12'ha;
        src100 <= 12'ha14;
        src101 <= 12'h2b6;
        src102 <= 12'hb68;
        src103 <= 12'h544;
        src104 <= 12'h885;
        src105 <= 12'hc53;
        src106 <= 12'he27;
        src107 <= 12'h3a0;
        src108 <= 12'h9ec;
        src109 <= 12'h923;
        src110 <= 12'hd64;
        src111 <= 12'h2b7;
        src112 <= 12'hc05;
        src113 <= 12'h26a;
        src114 <= 12'h7a4;
        src115 <= 12'h837;
        src116 <= 12'h3cb;
        src117 <= 12'ha3d;
        src118 <= 12'h84c;
        src119 <= 12'heed;
        src120 <= 12'h98b;
        src121 <= 12'h6f3;
        src122 <= 12'h99b;
        src123 <= 12'h800;
        src124 <= 12'h489;
        src125 <= 12'hc46;
        src126 <= 12'h5d1;
        src127 <= 12'ha8;
        src128 <= 12'hdc1;
        src129 <= 12'hbb0;
        src130 <= 12'hfb0;
        src131 <= 12'hf66;
        src132 <= 12'hfc4;
        src133 <= 12'hc7a;
        src134 <= 12'h898;
        src135 <= 12'h426;
        src136 <= 12'he7e;
        src137 <= 12'h3a3;
        src138 <= 12'h957;
        src139 <= 12'he02;
        src140 <= 12'h77e;
        src141 <= 12'ha43;
        src142 <= 12'h5d7;
        src143 <= 12'h350;
        src144 <= 12'h40d;
        src145 <= 12'hde2;
        src146 <= 12'hdee;
        src147 <= 12'hecf;
        src148 <= 12'h302;
        src149 <= 12'h923;
        src150 <= 12'hbff;
        src151 <= 12'h5fc;
        src152 <= 12'h495;
        src153 <= 12'h7e7;
        src154 <= 12'h127;
        src155 <= 12'h9c6;
        src156 <= 12'h69a;
        src157 <= 12'hcad;
        src158 <= 12'hd72;
        src159 <= 12'h600;
        src160 <= 12'h9b7;
        src161 <= 12'haf1;
        exp <= 20'h529a6;
        #1
        src0 <= 12'h49a;
        src1 <= 12'h2b9;
        src2 <= 12'h350;
        src3 <= 12'h28e;
        src4 <= 12'hb4d;
        src5 <= 12'h35;
        src6 <= 12'h29c;
        src7 <= 12'h807;
        src8 <= 12'hda0;
        src9 <= 12'hde5;
        src10 <= 12'h987;
        src11 <= 12'h1b6;
        src12 <= 12'hed6;
        src13 <= 12'hdf9;
        src14 <= 12'h392;
        src15 <= 12'he09;
        src16 <= 12'h144;
        src17 <= 12'h525;
        src18 <= 12'hbcc;
        src19 <= 12'h67e;
        src20 <= 12'h6c9;
        src21 <= 12'h785;
        src22 <= 12'h69;
        src23 <= 12'h9da;
        src24 <= 12'h614;
        src25 <= 12'h1bf;
        src26 <= 12'ha2f;
        src27 <= 12'h8a7;
        src28 <= 12'h5d;
        src29 <= 12'hc3a;
        src30 <= 12'h424;
        src31 <= 12'hba9;
        src32 <= 12'h4d;
        src33 <= 12'h76f;
        src34 <= 12'h3c8;
        src35 <= 12'h1d5;
        src36 <= 12'hc2d;
        src37 <= 12'h7c;
        src38 <= 12'h6e7;
        src39 <= 12'h4d8;
        src40 <= 12'ha16;
        src41 <= 12'h174;
        src42 <= 12'ha08;
        src43 <= 12'he97;
        src44 <= 12'h955;
        src45 <= 12'h9d1;
        src46 <= 12'h617;
        src47 <= 12'h56a;
        src48 <= 12'h6e5;
        src49 <= 12'hd7f;
        src50 <= 12'haac;
        src51 <= 12'hb;
        src52 <= 12'hac2;
        src53 <= 12'h529;
        src54 <= 12'h4a6;
        src55 <= 12'ha0d;
        src56 <= 12'hc70;
        src57 <= 12'hb00;
        src58 <= 12'h722;
        src59 <= 12'h455;
        src60 <= 12'he61;
        src61 <= 12'hd00;
        src62 <= 12'h900;
        src63 <= 12'h32f;
        src64 <= 12'h7bc;
        src65 <= 12'hf0;
        src66 <= 12'h362;
        src67 <= 12'he02;
        src68 <= 12'h43;
        src69 <= 12'h3eb;
        src70 <= 12'hbfc;
        src71 <= 12'h1fd;
        src72 <= 12'hae5;
        src73 <= 12'hd7c;
        src74 <= 12'h769;
        src75 <= 12'h45c;
        src76 <= 12'h332;
        src77 <= 12'hcfd;
        src78 <= 12'h374;
        src79 <= 12'h323;
        src80 <= 12'hb27;
        src81 <= 12'hd08;
        src82 <= 12'h2f;
        src83 <= 12'h523;
        src84 <= 12'hda5;
        src85 <= 12'h220;
        src86 <= 12'h490;
        src87 <= 12'he87;
        src88 <= 12'he1a;
        src89 <= 12'hedb;
        src90 <= 12'hf46;
        src91 <= 12'he8c;
        src92 <= 12'h64d;
        src93 <= 12'hea2;
        src94 <= 12'hc13;
        src95 <= 12'h2e9;
        src96 <= 12'h97a;
        src97 <= 12'h399;
        src98 <= 12'hdeb;
        src99 <= 12'he6c;
        src100 <= 12'h3b1;
        src101 <= 12'h35e;
        src102 <= 12'h9c9;
        src103 <= 12'h867;
        src104 <= 12'h7ce;
        src105 <= 12'hdb7;
        src106 <= 12'h260;
        src107 <= 12'h5dc;
        src108 <= 12'hf7f;
        src109 <= 12'h476;
        src110 <= 12'h180;
        src111 <= 12'hceb;
        src112 <= 12'hfdd;
        src113 <= 12'h952;
        src114 <= 12'h3b7;
        src115 <= 12'h2d7;
        src116 <= 12'h99a;
        src117 <= 12'h6c;
        src118 <= 12'h609;
        src119 <= 12'h10b;
        src120 <= 12'h962;
        src121 <= 12'h84c;
        src122 <= 12'h417;
        src123 <= 12'ha8a;
        src124 <= 12'hf45;
        src125 <= 12'hb13;
        src126 <= 12'h593;
        src127 <= 12'h3ad;
        src128 <= 12'had5;
        src129 <= 12'h32c;
        src130 <= 12'hd2;
        src131 <= 12'hc1d;
        src132 <= 12'hf5;
        src133 <= 12'h87a;
        src134 <= 12'h79d;
        src135 <= 12'he34;
        src136 <= 12'hfe7;
        src137 <= 12'h822;
        src138 <= 12'h8bc;
        src139 <= 12'h1ce;
        src140 <= 12'h7c8;
        src141 <= 12'he0c;
        src142 <= 12'h3d9;
        src143 <= 12'hc2f;
        src144 <= 12'h692;
        src145 <= 12'he00;
        src146 <= 12'h8ee;
        src147 <= 12'ha3a;
        src148 <= 12'h46b;
        src149 <= 12'h170;
        src150 <= 12'hf54;
        src151 <= 12'h8c1;
        src152 <= 12'h9b5;
        src153 <= 12'h150;
        src154 <= 12'he20;
        src155 <= 12'h939;
        src156 <= 12'h1e7;
        src157 <= 12'hf48;
        src158 <= 12'hef3;
        src159 <= 12'he9d;
        src160 <= 12'h18b;
        src161 <= 12'h7aa;
        exp <= 20'h4f1e9;
        #1
        src0 <= 12'hbc8;
        src1 <= 12'h1e0;
        src2 <= 12'hab1;
        src3 <= 12'h962;
        src4 <= 12'h8e2;
        src5 <= 12'ha8d;
        src6 <= 12'he62;
        src7 <= 12'h5ad;
        src8 <= 12'ha80;
        src9 <= 12'h54e;
        src10 <= 12'hc92;
        src11 <= 12'h39d;
        src12 <= 12'h554;
        src13 <= 12'h570;
        src14 <= 12'h3d;
        src15 <= 12'h5a0;
        src16 <= 12'h9dd;
        src17 <= 12'h7b3;
        src18 <= 12'hb0c;
        src19 <= 12'he8f;
        src20 <= 12'h5a4;
        src21 <= 12'hc97;
        src22 <= 12'hacf;
        src23 <= 12'h2d1;
        src24 <= 12'h8be;
        src25 <= 12'he25;
        src26 <= 12'h555;
        src27 <= 12'h21b;
        src28 <= 12'h8f8;
        src29 <= 12'h453;
        src30 <= 12'h6a7;
        src31 <= 12'hf07;
        src32 <= 12'haf3;
        src33 <= 12'h178;
        src34 <= 12'haca;
        src35 <= 12'ha15;
        src36 <= 12'hc21;
        src37 <= 12'hd00;
        src38 <= 12'hd19;
        src39 <= 12'h8f;
        src40 <= 12'h23c;
        src41 <= 12'hc7a;
        src42 <= 12'h77;
        src43 <= 12'h53;
        src44 <= 12'h2a7;
        src45 <= 12'ha6c;
        src46 <= 12'h45f;
        src47 <= 12'h215;
        src48 <= 12'hee2;
        src49 <= 12'ha2;
        src50 <= 12'h6a1;
        src51 <= 12'h374;
        src52 <= 12'h192;
        src53 <= 12'h960;
        src54 <= 12'h1ec;
        src55 <= 12'h10a;
        src56 <= 12'h935;
        src57 <= 12'hfc3;
        src58 <= 12'hbd3;
        src59 <= 12'h8c5;
        src60 <= 12'hf3;
        src61 <= 12'h768;
        src62 <= 12'hdc9;
        src63 <= 12'h421;
        src64 <= 12'ha50;
        src65 <= 12'h130;
        src66 <= 12'h9d0;
        src67 <= 12'h102;
        src68 <= 12'h4e6;
        src69 <= 12'h816;
        src70 <= 12'h78a;
        src71 <= 12'h2a5;
        src72 <= 12'hbc5;
        src73 <= 12'h576;
        src74 <= 12'h239;
        src75 <= 12'h7e4;
        src76 <= 12'h47d;
        src77 <= 12'h189;
        src78 <= 12'he0b;
        src79 <= 12'h854;
        src80 <= 12'h94a;
        src81 <= 12'h854;
        src82 <= 12'hbb4;
        src83 <= 12'h5d4;
        src84 <= 12'hd71;
        src85 <= 12'h82f;
        src86 <= 12'h425;
        src87 <= 12'h355;
        src88 <= 12'h567;
        src89 <= 12'hf25;
        src90 <= 12'h7bb;
        src91 <= 12'hd1b;
        src92 <= 12'h5d3;
        src93 <= 12'h6b6;
        src94 <= 12'h3f8;
        src95 <= 12'hb91;
        src96 <= 12'hbfa;
        src97 <= 12'h30c;
        src98 <= 12'hadb;
        src99 <= 12'he6e;
        src100 <= 12'h5e6;
        src101 <= 12'h59c;
        src102 <= 12'hf81;
        src103 <= 12'hc73;
        src104 <= 12'ha5b;
        src105 <= 12'h23f;
        src106 <= 12'h3f4;
        src107 <= 12'h786;
        src108 <= 12'hc38;
        src109 <= 12'h8f1;
        src110 <= 12'h646;
        src111 <= 12'h22b;
        src112 <= 12'h711;
        src113 <= 12'h431;
        src114 <= 12'h12e;
        src115 <= 12'hee9;
        src116 <= 12'h25a;
        src117 <= 12'hc7d;
        src118 <= 12'h2df;
        src119 <= 12'h1e8;
        src120 <= 12'h214;
        src121 <= 12'h43;
        src122 <= 12'h518;
        src123 <= 12'he42;
        src124 <= 12'h362;
        src125 <= 12'h736;
        src126 <= 12'h2f9;
        src127 <= 12'h5bd;
        src128 <= 12'hdee;
        src129 <= 12'hd38;
        src130 <= 12'hb3c;
        src131 <= 12'h40c;
        src132 <= 12'h360;
        src133 <= 12'h4d9;
        src134 <= 12'hcab;
        src135 <= 12'h161;
        src136 <= 12'hd86;
        src137 <= 12'h623;
        src138 <= 12'h733;
        src139 <= 12'hcb6;
        src140 <= 12'h540;
        src141 <= 12'hd48;
        src142 <= 12'h4e2;
        src143 <= 12'he7f;
        src144 <= 12'h9d2;
        src145 <= 12'h8ee;
        src146 <= 12'ha1b;
        src147 <= 12'h289;
        src148 <= 12'h26f;
        src149 <= 12'h446;
        src150 <= 12'h989;
        src151 <= 12'hf16;
        src152 <= 12'h63a;
        src153 <= 12'h374;
        src154 <= 12'hdef;
        src155 <= 12'h69;
        src156 <= 12'h77f;
        src157 <= 12'h74;
        src158 <= 12'h51;
        src159 <= 12'h131;
        src160 <= 12'h427;
        src161 <= 12'hc8c;
        exp <= 20'h4a804;
        #1
        src0 <= 12'h5d6;
        src1 <= 12'hafb;
        src2 <= 12'h39e;
        src3 <= 12'ha12;
        src4 <= 12'h9ef;
        src5 <= 12'h7f;
        src6 <= 12'h48d;
        src7 <= 12'hf;
        src8 <= 12'h773;
        src9 <= 12'h37b;
        src10 <= 12'ha2b;
        src11 <= 12'h772;
        src12 <= 12'h37;
        src13 <= 12'h618;
        src14 <= 12'h553;
        src15 <= 12'h40d;
        src16 <= 12'h605;
        src17 <= 12'h31d;
        src18 <= 12'h711;
        src19 <= 12'hfd9;
        src20 <= 12'h924;
        src21 <= 12'hc6b;
        src22 <= 12'hf67;
        src23 <= 12'hc49;
        src24 <= 12'h60b;
        src25 <= 12'h139;
        src26 <= 12'h721;
        src27 <= 12'hddf;
        src28 <= 12'h8aa;
        src29 <= 12'h126;
        src30 <= 12'ha36;
        src31 <= 12'h668;
        src32 <= 12'hd93;
        src33 <= 12'h7a;
        src34 <= 12'hdb1;
        src35 <= 12'ha45;
        src36 <= 12'h4ca;
        src37 <= 12'h5e7;
        src38 <= 12'hb7a;
        src39 <= 12'h2e3;
        src40 <= 12'hcd0;
        src41 <= 12'h809;
        src42 <= 12'hf83;
        src43 <= 12'hee0;
        src44 <= 12'h850;
        src45 <= 12'h67f;
        src46 <= 12'h3f7;
        src47 <= 12'ha20;
        src48 <= 12'h4d5;
        src49 <= 12'h484;
        src50 <= 12'hd8e;
        src51 <= 12'h32d;
        src52 <= 12'hea5;
        src53 <= 12'hbc3;
        src54 <= 12'h2ef;
        src55 <= 12'h4e4;
        src56 <= 12'h550;
        src57 <= 12'hd37;
        src58 <= 12'h518;
        src59 <= 12'he57;
        src60 <= 12'h1c5;
        src61 <= 12'h924;
        src62 <= 12'h3b4;
        src63 <= 12'h953;
        src64 <= 12'h34a;
        src65 <= 12'h6c5;
        src66 <= 12'h113;
        src67 <= 12'h61;
        src68 <= 12'h750;
        src69 <= 12'hf53;
        src70 <= 12'h6ec;
        src71 <= 12'h413;
        src72 <= 12'h9f;
        src73 <= 12'hde;
        src74 <= 12'h6ca;
        src75 <= 12'h406;
        src76 <= 12'hd4c;
        src77 <= 12'h61;
        src78 <= 12'hd0c;
        src79 <= 12'h948;
        src80 <= 12'h90f;
        src81 <= 12'hc47;
        src82 <= 12'h162;
        src83 <= 12'hd46;
        src84 <= 12'haa7;
        src85 <= 12'ha72;
        src86 <= 12'hae0;
        src87 <= 12'h114;
        src88 <= 12'hd94;
        src89 <= 12'h632;
        src90 <= 12'h834;
        src91 <= 12'ha30;
        src92 <= 12'h58;
        src93 <= 12'h37b;
        src94 <= 12'h8f1;
        src95 <= 12'h596;
        src96 <= 12'h89b;
        src97 <= 12'hc42;
        src98 <= 12'hfc5;
        src99 <= 12'ha28;
        src100 <= 12'haec;
        src101 <= 12'h464;
        src102 <= 12'h649;
        src103 <= 12'h313;
        src104 <= 12'h228;
        src105 <= 12'hf73;
        src106 <= 12'hd25;
        src107 <= 12'hc64;
        src108 <= 12'h48;
        src109 <= 12'h332;
        src110 <= 12'hc15;
        src111 <= 12'hca5;
        src112 <= 12'h41b;
        src113 <= 12'h113;
        src114 <= 12'h8a4;
        src115 <= 12'hf66;
        src116 <= 12'h5eb;
        src117 <= 12'h573;
        src118 <= 12'hc3;
        src119 <= 12'h6f8;
        src120 <= 12'h143;
        src121 <= 12'h349;
        src122 <= 12'hd2d;
        src123 <= 12'hc4b;
        src124 <= 12'h7b6;
        src125 <= 12'ha2;
        src126 <= 12'h354;
        src127 <= 12'h8a6;
        src128 <= 12'h938;
        src129 <= 12'h79;
        src130 <= 12'hdbb;
        src131 <= 12'h487;
        src132 <= 12'hd9;
        src133 <= 12'h7af;
        src134 <= 12'h848;
        src135 <= 12'h648;
        src136 <= 12'h9a6;
        src137 <= 12'h69f;
        src138 <= 12'h3e9;
        src139 <= 12'h52f;
        src140 <= 12'hfb;
        src141 <= 12'h6da;
        src142 <= 12'hc66;
        src143 <= 12'hac;
        src144 <= 12'h835;
        src145 <= 12'hadb;
        src146 <= 12'h8e4;
        src147 <= 12'h889;
        src148 <= 12'he2b;
        src149 <= 12'h40e;
        src150 <= 12'h654;
        src151 <= 12'h7fe;
        src152 <= 12'hb0;
        src153 <= 12'h4da;
        src154 <= 12'h47a;
        src155 <= 12'hd84;
        src156 <= 12'h69a;
        src157 <= 12'he04;
        src158 <= 12'ha32;
        src159 <= 12'hf5a;
        src160 <= 12'h546;
        src161 <= 12'h15;
        exp <= 20'h4a905;
        #1
        src0 <= 12'ha83;
        src1 <= 12'hc84;
        src2 <= 12'hb64;
        src3 <= 12'h54b;
        src4 <= 12'h7b6;
        src5 <= 12'hf6c;
        src6 <= 12'hc41;
        src7 <= 12'hcb8;
        src8 <= 12'h536;
        src9 <= 12'ha06;
        src10 <= 12'hd1d;
        src11 <= 12'hee4;
        src12 <= 12'hdbd;
        src13 <= 12'h8fd;
        src14 <= 12'h716;
        src15 <= 12'h8fc;
        src16 <= 12'hbe3;
        src17 <= 12'h71;
        src18 <= 12'h1ba;
        src19 <= 12'hefe;
        src20 <= 12'h9bb;
        src21 <= 12'hc2c;
        src22 <= 12'h16e;
        src23 <= 12'hd6;
        src24 <= 12'h204;
        src25 <= 12'hb93;
        src26 <= 12'hc05;
        src27 <= 12'h303;
        src28 <= 12'h9be;
        src29 <= 12'hafc;
        src30 <= 12'h1ad;
        src31 <= 12'hb97;
        src32 <= 12'h9e4;
        src33 <= 12'he42;
        src34 <= 12'h45c;
        src35 <= 12'hb04;
        src36 <= 12'h37c;
        src37 <= 12'h8b4;
        src38 <= 12'hf25;
        src39 <= 12'h151;
        src40 <= 12'hdb1;
        src41 <= 12'hc73;
        src42 <= 12'h96f;
        src43 <= 12'h67c;
        src44 <= 12'h6c3;
        src45 <= 12'h77;
        src46 <= 12'h1fd;
        src47 <= 12'hb1f;
        src48 <= 12'hd41;
        src49 <= 12'h4ef;
        src50 <= 12'hed8;
        src51 <= 12'h3b3;
        src52 <= 12'h2c9;
        src53 <= 12'hb52;
        src54 <= 12'hc69;
        src55 <= 12'he4f;
        src56 <= 12'h5b;
        src57 <= 12'h100;
        src58 <= 12'h72b;
        src59 <= 12'h670;
        src60 <= 12'h507;
        src61 <= 12'hd99;
        src62 <= 12'h78c;
        src63 <= 12'h4f4;
        src64 <= 12'h1ac;
        src65 <= 12'h94;
        src66 <= 12'h6aa;
        src67 <= 12'hb1e;
        src68 <= 12'h34b;
        src69 <= 12'h860;
        src70 <= 12'h693;
        src71 <= 12'h7d6;
        src72 <= 12'h2af;
        src73 <= 12'ha96;
        src74 <= 12'hbb6;
        src75 <= 12'h2fe;
        src76 <= 12'h26;
        src77 <= 12'h396;
        src78 <= 12'h71;
        src79 <= 12'hc31;
        src80 <= 12'hcfc;
        src81 <= 12'h17b;
        src82 <= 12'h375;
        src83 <= 12'hbd8;
        src84 <= 12'hc51;
        src85 <= 12'hc75;
        src86 <= 12'h246;
        src87 <= 12'h272;
        src88 <= 12'h84d;
        src89 <= 12'h94a;
        src90 <= 12'h108;
        src91 <= 12'hbf4;
        src92 <= 12'h8b1;
        src93 <= 12'h801;
        src94 <= 12'h180;
        src95 <= 12'h6dc;
        src96 <= 12'hfe6;
        src97 <= 12'h84;
        src98 <= 12'hce7;
        src99 <= 12'h72c;
        src100 <= 12'h910;
        src101 <= 12'h57b;
        src102 <= 12'h5d;
        src103 <= 12'hb0a;
        src104 <= 12'h9e4;
        src105 <= 12'h3c4;
        src106 <= 12'hdaf;
        src107 <= 12'h8d1;
        src108 <= 12'h4fe;
        src109 <= 12'hf6;
        src110 <= 12'h636;
        src111 <= 12'h6e3;
        src112 <= 12'h9a4;
        src113 <= 12'h8b4;
        src114 <= 12'ha07;
        src115 <= 12'h704;
        src116 <= 12'h6fc;
        src117 <= 12'h86f;
        src118 <= 12'h37f;
        src119 <= 12'h949;
        src120 <= 12'h76;
        src121 <= 12'h990;
        src122 <= 12'h9c4;
        src123 <= 12'h609;
        src124 <= 12'ha35;
        src125 <= 12'ha5e;
        src126 <= 12'h198;
        src127 <= 12'h934;
        src128 <= 12'ha22;
        src129 <= 12'ha51;
        src130 <= 12'h6e;
        src131 <= 12'h3b3;
        src132 <= 12'h95c;
        src133 <= 12'h60d;
        src134 <= 12'h433;
        src135 <= 12'hd49;
        src136 <= 12'h813;
        src137 <= 12'h14f;
        src138 <= 12'hd4a;
        src139 <= 12'h941;
        src140 <= 12'h3b0;
        src141 <= 12'h4e;
        src142 <= 12'h8e6;
        src143 <= 12'ha8d;
        src144 <= 12'h8e;
        src145 <= 12'h62e;
        src146 <= 12'h4cc;
        src147 <= 12'h8d1;
        src148 <= 12'h36b;
        src149 <= 12'h609;
        src150 <= 12'h78;
        src151 <= 12'heef;
        src152 <= 12'h373;
        src153 <= 12'h264;
        src154 <= 12'hc9c;
        src155 <= 12'haab;
        src156 <= 12'hf81;
        src157 <= 12'hbf0;
        src158 <= 12'h118;
        src159 <= 12'h899;
        src160 <= 12'h502;
        src161 <= 12'hd01;
        exp <= 20'h4c9f3;
        #1
        $finish;
    end
endmodule

