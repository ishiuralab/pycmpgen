module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    compressor2_1_54_32 compressor2_1_54_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_54_32(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [0:0] comp_out37;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37)
    );
    rowadder2_1_38 rowadder2_1inst(
        .src0({comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [0:0] dst37);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [15:0] stage1_0;
   wire [16:0] stage1_1;
   wire [21:0] stage1_2;
   wire [21:0] stage1_3;
   wire [32:0] stage1_4;
   wire [26:0] stage1_5;
   wire [32:0] stage1_6;
   wire [20:0] stage1_7;
   wire [25:0] stage1_8;
   wire [35:0] stage1_9;
   wire [17:0] stage1_10;
   wire [28:0] stage1_11;
   wire [23:0] stage1_12;
   wire [31:0] stage1_13;
   wire [30:0] stage1_14;
   wire [27:0] stage1_15;
   wire [24:0] stage1_16;
   wire [19:0] stage1_17;
   wire [29:0] stage1_18;
   wire [31:0] stage1_19;
   wire [22:0] stage1_20;
   wire [29:0] stage1_21;
   wire [21:0] stage1_22;
   wire [28:0] stage1_23;
   wire [23:0] stage1_24;
   wire [22:0] stage1_25;
   wire [17:0] stage1_26;
   wire [24:0] stage1_27;
   wire [25:0] stage1_28;
   wire [24:0] stage1_29;
   wire [17:0] stage1_30;
   wire [23:0] stage1_31;
   wire [16:0] stage1_32;
   wire [7:0] stage1_33;
   wire [9:0] stage2_0;
   wire [11:0] stage2_1;
   wire [16:0] stage2_2;
   wire [10:0] stage2_3;
   wire [9:0] stage2_4;
   wire [11:0] stage2_5;
   wire [11:0] stage2_6;
   wire [15:0] stage2_7;
   wire [16:0] stage2_8;
   wire [9:0] stage2_9;
   wire [8:0] stage2_10;
   wire [9:0] stage2_11;
   wire [15:0] stage2_12;
   wire [18:0] stage2_13;
   wire [9:0] stage2_14;
   wire [11:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [13:0] stage2_18;
   wire [9:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [16:0] stage2_22;
   wire [16:0] stage2_23;
   wire [17:0] stage2_24;
   wire [11:0] stage2_25;
   wire [8:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [10:0] stage2_30;
   wire [9:0] stage2_31;
   wire [6:0] stage2_32;
   wire [6:0] stage2_33;
   wire [3:0] stage2_34;
   wire [1:0] stage2_35;
   wire [1:0] stage3_0;
   wire [11:0] stage3_1;
   wire [2:0] stage3_2;
   wire [12:0] stage3_3;
   wire [4:0] stage3_4;
   wire [2:0] stage3_5;
   wire [4:0] stage3_6;
   wire [8:0] stage3_7;
   wire [8:0] stage3_8;
   wire [7:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [5:0] stage3_12;
   wire [6:0] stage3_13;
   wire [5:0] stage3_14;
   wire [5:0] stage3_15;
   wire [8:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [6:0] stage3_19;
   wire [7:0] stage3_20;
   wire [6:0] stage3_21;
   wire [7:0] stage3_22;
   wire [6:0] stage3_23;
   wire [4:0] stage3_24;
   wire [5:0] stage3_25;
   wire [9:0] stage3_26;
   wire [2:0] stage3_27;
   wire [3:0] stage3_28;
   wire [18:0] stage3_29;
   wire [2:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [4:0] stage3_34;
   wire [3:0] stage3_35;
   wire [1:0] stage4_0;
   wire [3:0] stage4_1;
   wire [2:0] stage4_2;
   wire [2:0] stage4_3;
   wire [2:0] stage4_4;
   wire [2:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [4:0] stage4_8;
   wire [3:0] stage4_9;
   wire [4:0] stage4_10;
   wire [2:0] stage4_11;
   wire [1:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [3:0] stage4_15;
   wire [5:0] stage4_16;
   wire [1:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [2:0] stage4_21;
   wire [5:0] stage4_22;
   wire [2:0] stage4_23;
   wire [1:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [0:0] stage4_27;
   wire [1:0] stage4_28;
   wire [5:0] stage4_29;
   wire [4:0] stage4_30;
   wire [5:0] stage4_31;
   wire [3:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [0:0] stage4_37;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [0:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [0:0] stage5_37;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[15]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_1[16]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7]},
      {stage1_6[0],stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15]}
   );
   gpc606_5 gpc16 (
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13]},
      {stage1_6[1],stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc606_5 gpc17 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage1_6[2],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc606_5 gpc18 (
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage0_4[20]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[2],stage1_6[5],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[3],stage1_6[6],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[4],stage1_6[7],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[5],stage1_6[8],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[4],stage1_7[6],stage1_6[9],stage1_5[15]}
   );
   gpc606_5 gpc25 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[5],stage1_7[7],stage1_6[10],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[6],stage1_7[8],stage1_6[11],stage1_5[17]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[7],stage1_7[9],stage1_6[12],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[8],stage1_7[10],stage1_6[13],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[9],stage1_7[11],stage1_6[14],stage1_5[20]}
   );
   gpc615_5 gpc30 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28]},
      {stage0_7[36]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[6],stage1_8[10],stage1_7[12],stage1_6[15]}
   );
   gpc615_5 gpc31 (
      {stage0_6[29], stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33]},
      {stage0_7[37]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[7],stage1_8[11],stage1_7[13],stage1_6[16]}
   );
   gpc615_5 gpc32 (
      {stage0_6[34], stage0_6[35], stage0_6[36], stage0_6[37], stage0_6[38]},
      {stage0_7[38]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[8],stage1_8[12],stage1_7[14],stage1_6[17]}
   );
   gpc606_5 gpc33 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43], stage0_7[44]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[9],stage1_8[13],stage1_7[15]}
   );
   gpc615_5 gpc34 (
      {stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49]},
      {stage0_8[18]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[10],stage1_8[14],stage1_7[16]}
   );
   gpc1163_5 gpc35 (
      {stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_10[0]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[11],stage1_8[15]}
   );
   gpc606_5 gpc36 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[12],stage1_8[16]}
   );
   gpc606_5 gpc37 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[13],stage1_8[17]}
   );
   gpc615_5 gpc38 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[18]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[14],stage1_8[18]}
   );
   gpc615_5 gpc39 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[19]},
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[15],stage1_8[19]}
   );
   gpc615_5 gpc40 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[20]},
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[16],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[17]}
   );
   gpc606_5 gpc42 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[18]}
   );
   gpc615_5 gpc43 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_10[31]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[19]}
   );
   gpc606_5 gpc44 (
      {stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[9],stage1_11[11],stage1_10[14]}
   );
   gpc606_5 gpc45 (
      {stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[10],stage1_11[12],stage1_10[15]}
   );
   gpc615_5 gpc46 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[19]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[11],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc47 (
      {stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_11[20]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[12],stage1_11[14],stage1_10[17]}
   );
   gpc606_5 gpc48 (
      {stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[4],stage1_13[7],stage1_12[13],stage1_11[15]}
   );
   gpc606_5 gpc49 (
      {stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[5],stage1_13[8],stage1_12[14],stage1_11[16]}
   );
   gpc606_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[6],stage1_13[9],stage1_12[15],stage1_11[17]}
   );
   gpc615_5 gpc51 (
      {stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43]},
      {stage0_12[24]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[7],stage1_13[10],stage1_12[16],stage1_11[18]}
   );
   gpc1423_5 gpc52 (
      {stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage0_13[24], stage0_13[25]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[4],stage1_14[8],stage1_13[11],stage1_12[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9]},
      {stage1_16[1],stage1_15[5],stage1_14[9],stage1_13[12],stage1_12[18]}
   );
   gpc606_5 gpc54 (
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage1_16[2],stage1_15[6],stage1_14[10],stage1_13[13],stage1_12[19]}
   );
   gpc606_5 gpc55 (
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21]},
      {stage1_16[3],stage1_15[7],stage1_14[11],stage1_13[14],stage1_12[20]}
   );
   gpc606_5 gpc56 (
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage1_16[4],stage1_15[8],stage1_14[12],stage1_13[15],stage1_12[21]}
   );
   gpc615_5 gpc57 (
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30]},
      {stage0_14[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[5],stage1_15[9],stage1_14[13],stage1_13[16]}
   );
   gpc615_5 gpc58 (
      {stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_14[29]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[1],stage1_16[6],stage1_15[10],stage1_14[14],stage1_13[17]}
   );
   gpc615_5 gpc59 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_14[30]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[2],stage1_16[7],stage1_15[11],stage1_14[15],stage1_13[18]}
   );
   gpc615_5 gpc60 (
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_15[19]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[8],stage1_15[12],stage1_14[16]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[20]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[9],stage1_15[13],stage1_14[17]}
   );
   gpc606_5 gpc62 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25], stage0_15[26]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[2],stage1_17[5],stage1_16[10],stage1_15[14]}
   );
   gpc606_5 gpc63 (
      {stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30], stage0_15[31], stage0_15[32]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[3],stage1_17[6],stage1_16[11],stage1_15[15]}
   );
   gpc606_5 gpc64 (
      {stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36], stage0_15[37], stage0_15[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[4],stage1_17[7],stage1_16[12],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[39], stage0_15[40], stage0_15[41], stage0_15[42], stage0_15[43]},
      {stage0_16[12]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[5],stage1_17[8],stage1_16[13],stage1_15[17]}
   );
   gpc606_5 gpc66 (
      {stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[4],stage1_18[6],stage1_17[9],stage1_16[14]}
   );
   gpc606_5 gpc67 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[5],stage1_18[7],stage1_17[10],stage1_16[15]}
   );
   gpc606_5 gpc68 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[6],stage1_18[8],stage1_17[11],stage1_16[16]}
   );
   gpc606_5 gpc69 (
      {stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[7],stage1_18[9],stage1_17[12],stage1_16[17]}
   );
   gpc606_5 gpc70 (
      {stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[8],stage1_18[10],stage1_17[13],stage1_16[18]}
   );
   gpc606_5 gpc71 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[9],stage1_18[11],stage1_17[14],stage1_16[19]}
   );
   gpc606_5 gpc72 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[6],stage1_19[10],stage1_18[12],stage1_17[15]}
   );
   gpc606_5 gpc73 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[7],stage1_19[11],stage1_18[13],stage1_17[16]}
   );
   gpc606_5 gpc74 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[8],stage1_19[12],stage1_18[14],stage1_17[17]}
   );
   gpc606_5 gpc75 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[9],stage1_19[13],stage1_18[15],stage1_17[18]}
   );
   gpc606_5 gpc76 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[10],stage1_19[14],stage1_18[16],stage1_17[19]}
   );
   gpc606_5 gpc77 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[5],stage1_20[11],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc78 (
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34]},
      {stage0_20[6]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[1],stage1_21[6],stage1_20[12],stage1_19[16]}
   );
   gpc615_5 gpc79 (
      {stage0_19[35], stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39]},
      {stage0_20[7]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[2],stage1_21[7],stage1_20[13],stage1_19[17]}
   );
   gpc606_5 gpc80 (
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[3],stage1_21[8],stage1_20[14]}
   );
   gpc606_5 gpc81 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[4],stage1_21[9],stage1_20[15]}
   );
   gpc606_5 gpc82 (
      {stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[5],stage1_21[10],stage1_20[16]}
   );
   gpc606_5 gpc83 (
      {stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[6],stage1_21[11],stage1_20[17]}
   );
   gpc606_5 gpc84 (
      {stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[7],stage1_21[12],stage1_20[18]}
   );
   gpc615_5 gpc85 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[12]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[8],stage1_21[13],stage1_20[19]}
   );
   gpc615_5 gpc86 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[13]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[9],stage1_21[14],stage1_20[20]}
   );
   gpc615_5 gpc87 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[14]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[10],stage1_21[15],stage1_20[21]}
   );
   gpc606_5 gpc88 (
      {stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[8],stage1_23[10],stage1_22[11],stage1_21[16]}
   );
   gpc606_5 gpc89 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[9],stage1_23[11],stage1_22[12],stage1_21[17]}
   );
   gpc606_5 gpc90 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[10],stage1_23[12],stage1_22[13],stage1_21[18]}
   );
   gpc606_5 gpc91 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[11],stage1_23[13],stage1_22[14],stage1_21[19]}
   );
   gpc606_5 gpc92 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[12],stage1_23[14],stage1_22[15],stage1_21[20]}
   );
   gpc606_5 gpc93 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[5],stage1_24[13],stage1_23[15]}
   );
   gpc606_5 gpc94 (
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[6],stage1_24[14],stage1_23[16]}
   );
   gpc606_5 gpc95 (
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[2],stage1_25[7],stage1_24[15]}
   );
   gpc606_5 gpc96 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[3],stage1_25[8],stage1_24[16]}
   );
   gpc606_5 gpc97 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[4],stage1_25[9],stage1_24[17]}
   );
   gpc606_5 gpc98 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[5],stage1_25[10],stage1_24[18]}
   );
   gpc606_5 gpc99 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[6],stage1_25[11],stage1_24[19]}
   );
   gpc606_5 gpc100 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[7],stage1_25[12],stage1_24[20]}
   );
   gpc606_5 gpc101 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[8],stage1_25[13],stage1_24[21]}
   );
   gpc606_5 gpc102 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[9],stage1_25[14],stage1_24[22]}
   );
   gpc606_5 gpc103 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[10],stage1_26[10],stage1_25[15],stage1_24[23]}
   );
   gpc606_5 gpc104 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[9],stage1_27[11],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc105 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[10],stage1_27[12],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc106 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[11],stage1_27[13],stage1_26[13],stage1_25[18]}
   );
   gpc606_5 gpc107 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[12],stage1_27[14],stage1_26[14],stage1_25[19]}
   );
   gpc606_5 gpc108 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[13],stage1_27[15],stage1_26[15],stage1_25[20]}
   );
   gpc606_5 gpc109 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[14],stage1_27[16],stage1_26[16],stage1_25[21]}
   );
   gpc606_5 gpc110 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[15],stage1_27[17],stage1_26[17],stage1_25[22]}
   );
   gpc606_5 gpc111 (
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[7],stage1_28[16],stage1_27[18]}
   );
   gpc606_5 gpc112 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[1],stage1_30[1],stage1_29[8],stage1_28[17]}
   );
   gpc606_5 gpc113 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[2],stage1_30[2],stage1_29[9],stage1_28[18]}
   );
   gpc606_5 gpc114 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[3],stage1_30[3],stage1_29[10],stage1_28[19]}
   );
   gpc606_5 gpc115 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[4],stage1_30[4],stage1_29[11],stage1_28[20]}
   );
   gpc606_5 gpc116 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[5],stage1_30[5],stage1_29[12],stage1_28[21]}
   );
   gpc606_5 gpc117 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[6],stage1_30[6],stage1_29[13],stage1_28[22]}
   );
   gpc606_5 gpc118 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[7],stage1_30[7],stage1_29[14],stage1_28[23]}
   );
   gpc606_5 gpc119 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[8],stage1_30[8],stage1_29[15],stage1_28[24]}
   );
   gpc606_5 gpc120 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[9],stage1_30[9],stage1_29[16],stage1_28[25]}
   );
   gpc606_5 gpc121 (
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[10],stage1_30[10],stage1_29[17]}
   );
   gpc606_5 gpc122 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[11],stage1_30[11],stage1_29[18]}
   );
   gpc606_5 gpc123 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[12],stage1_30[12],stage1_29[19]}
   );
   gpc606_5 gpc124 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[13],stage1_30[13],stage1_29[20]}
   );
   gpc606_5 gpc125 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[14],stage1_30[14],stage1_29[21]}
   );
   gpc606_5 gpc126 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[15],stage1_30[15],stage1_29[22]}
   );
   gpc606_5 gpc127 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[16],stage1_30[16],stage1_29[23]}
   );
   gpc606_5 gpc128 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[17],stage1_30[17],stage1_29[24]}
   );
   gpc1_1 gpc129 (
      {stage0_0[47]},
      {stage1_0[9]}
   );
   gpc1_1 gpc130 (
      {stage0_0[48]},
      {stage1_0[10]}
   );
   gpc1_1 gpc131 (
      {stage0_0[49]},
      {stage1_0[11]}
   );
   gpc1_1 gpc132 (
      {stage0_0[50]},
      {stage1_0[12]}
   );
   gpc1_1 gpc133 (
      {stage0_0[51]},
      {stage1_0[13]}
   );
   gpc1_1 gpc134 (
      {stage0_0[52]},
      {stage1_0[14]}
   );
   gpc1_1 gpc135 (
      {stage0_0[53]},
      {stage1_0[15]}
   );
   gpc1_1 gpc136 (
      {stage0_1[52]},
      {stage1_1[15]}
   );
   gpc1_1 gpc137 (
      {stage0_1[53]},
      {stage1_1[16]}
   );
   gpc1_1 gpc138 (
      {stage0_2[50]},
      {stage1_2[18]}
   );
   gpc1_1 gpc139 (
      {stage0_2[51]},
      {stage1_2[19]}
   );
   gpc1_1 gpc140 (
      {stage0_2[52]},
      {stage1_2[20]}
   );
   gpc1_1 gpc141 (
      {stage0_2[53]},
      {stage1_2[21]}
   );
   gpc1_1 gpc142 (
      {stage0_3[52]},
      {stage1_3[20]}
   );
   gpc1_1 gpc143 (
      {stage0_3[53]},
      {stage1_3[21]}
   );
   gpc1_1 gpc144 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc145 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc146 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc147 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc148 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc149 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc150 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc151 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc152 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc153 (
      {stage0_5[48]},
      {stage1_5[21]}
   );
   gpc1_1 gpc154 (
      {stage0_5[49]},
      {stage1_5[22]}
   );
   gpc1_1 gpc155 (
      {stage0_5[50]},
      {stage1_5[23]}
   );
   gpc1_1 gpc156 (
      {stage0_5[51]},
      {stage1_5[24]}
   );
   gpc1_1 gpc157 (
      {stage0_5[52]},
      {stage1_5[25]}
   );
   gpc1_1 gpc158 (
      {stage0_5[53]},
      {stage1_5[26]}
   );
   gpc1_1 gpc159 (
      {stage0_6[39]},
      {stage1_6[18]}
   );
   gpc1_1 gpc160 (
      {stage0_6[40]},
      {stage1_6[19]}
   );
   gpc1_1 gpc161 (
      {stage0_6[41]},
      {stage1_6[20]}
   );
   gpc1_1 gpc162 (
      {stage0_6[42]},
      {stage1_6[21]}
   );
   gpc1_1 gpc163 (
      {stage0_6[43]},
      {stage1_6[22]}
   );
   gpc1_1 gpc164 (
      {stage0_6[44]},
      {stage1_6[23]}
   );
   gpc1_1 gpc165 (
      {stage0_6[45]},
      {stage1_6[24]}
   );
   gpc1_1 gpc166 (
      {stage0_6[46]},
      {stage1_6[25]}
   );
   gpc1_1 gpc167 (
      {stage0_6[47]},
      {stage1_6[26]}
   );
   gpc1_1 gpc168 (
      {stage0_6[48]},
      {stage1_6[27]}
   );
   gpc1_1 gpc169 (
      {stage0_6[49]},
      {stage1_6[28]}
   );
   gpc1_1 gpc170 (
      {stage0_6[50]},
      {stage1_6[29]}
   );
   gpc1_1 gpc171 (
      {stage0_6[51]},
      {stage1_6[30]}
   );
   gpc1_1 gpc172 (
      {stage0_6[52]},
      {stage1_6[31]}
   );
   gpc1_1 gpc173 (
      {stage0_6[53]},
      {stage1_6[32]}
   );
   gpc1_1 gpc174 (
      {stage0_7[50]},
      {stage1_7[17]}
   );
   gpc1_1 gpc175 (
      {stage0_7[51]},
      {stage1_7[18]}
   );
   gpc1_1 gpc176 (
      {stage0_7[52]},
      {stage1_7[19]}
   );
   gpc1_1 gpc177 (
      {stage0_7[53]},
      {stage1_7[20]}
   );
   gpc1_1 gpc178 (
      {stage0_8[49]},
      {stage1_8[21]}
   );
   gpc1_1 gpc179 (
      {stage0_8[50]},
      {stage1_8[22]}
   );
   gpc1_1 gpc180 (
      {stage0_8[51]},
      {stage1_8[23]}
   );
   gpc1_1 gpc181 (
      {stage0_8[52]},
      {stage1_8[24]}
   );
   gpc1_1 gpc182 (
      {stage0_8[53]},
      {stage1_8[25]}
   );
   gpc1_1 gpc183 (
      {stage0_9[38]},
      {stage1_9[20]}
   );
   gpc1_1 gpc184 (
      {stage0_9[39]},
      {stage1_9[21]}
   );
   gpc1_1 gpc185 (
      {stage0_9[40]},
      {stage1_9[22]}
   );
   gpc1_1 gpc186 (
      {stage0_9[41]},
      {stage1_9[23]}
   );
   gpc1_1 gpc187 (
      {stage0_9[42]},
      {stage1_9[24]}
   );
   gpc1_1 gpc188 (
      {stage0_9[43]},
      {stage1_9[25]}
   );
   gpc1_1 gpc189 (
      {stage0_9[44]},
      {stage1_9[26]}
   );
   gpc1_1 gpc190 (
      {stage0_9[45]},
      {stage1_9[27]}
   );
   gpc1_1 gpc191 (
      {stage0_9[46]},
      {stage1_9[28]}
   );
   gpc1_1 gpc192 (
      {stage0_9[47]},
      {stage1_9[29]}
   );
   gpc1_1 gpc193 (
      {stage0_9[48]},
      {stage1_9[30]}
   );
   gpc1_1 gpc194 (
      {stage0_9[49]},
      {stage1_9[31]}
   );
   gpc1_1 gpc195 (
      {stage0_9[50]},
      {stage1_9[32]}
   );
   gpc1_1 gpc196 (
      {stage0_9[51]},
      {stage1_9[33]}
   );
   gpc1_1 gpc197 (
      {stage0_9[52]},
      {stage1_9[34]}
   );
   gpc1_1 gpc198 (
      {stage0_9[53]},
      {stage1_9[35]}
   );
   gpc1_1 gpc199 (
      {stage0_11[44]},
      {stage1_11[19]}
   );
   gpc1_1 gpc200 (
      {stage0_11[45]},
      {stage1_11[20]}
   );
   gpc1_1 gpc201 (
      {stage0_11[46]},
      {stage1_11[21]}
   );
   gpc1_1 gpc202 (
      {stage0_11[47]},
      {stage1_11[22]}
   );
   gpc1_1 gpc203 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc204 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc205 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc206 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc207 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc208 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc209 (
      {stage0_12[52]},
      {stage1_12[22]}
   );
   gpc1_1 gpc210 (
      {stage0_12[53]},
      {stage1_12[23]}
   );
   gpc1_1 gpc211 (
      {stage0_13[41]},
      {stage1_13[19]}
   );
   gpc1_1 gpc212 (
      {stage0_13[42]},
      {stage1_13[20]}
   );
   gpc1_1 gpc213 (
      {stage0_13[43]},
      {stage1_13[21]}
   );
   gpc1_1 gpc214 (
      {stage0_13[44]},
      {stage1_13[22]}
   );
   gpc1_1 gpc215 (
      {stage0_13[45]},
      {stage1_13[23]}
   );
   gpc1_1 gpc216 (
      {stage0_13[46]},
      {stage1_13[24]}
   );
   gpc1_1 gpc217 (
      {stage0_13[47]},
      {stage1_13[25]}
   );
   gpc1_1 gpc218 (
      {stage0_13[48]},
      {stage1_13[26]}
   );
   gpc1_1 gpc219 (
      {stage0_13[49]},
      {stage1_13[27]}
   );
   gpc1_1 gpc220 (
      {stage0_13[50]},
      {stage1_13[28]}
   );
   gpc1_1 gpc221 (
      {stage0_13[51]},
      {stage1_13[29]}
   );
   gpc1_1 gpc222 (
      {stage0_13[52]},
      {stage1_13[30]}
   );
   gpc1_1 gpc223 (
      {stage0_13[53]},
      {stage1_13[31]}
   );
   gpc1_1 gpc224 (
      {stage0_14[41]},
      {stage1_14[18]}
   );
   gpc1_1 gpc225 (
      {stage0_14[42]},
      {stage1_14[19]}
   );
   gpc1_1 gpc226 (
      {stage0_14[43]},
      {stage1_14[20]}
   );
   gpc1_1 gpc227 (
      {stage0_14[44]},
      {stage1_14[21]}
   );
   gpc1_1 gpc228 (
      {stage0_14[45]},
      {stage1_14[22]}
   );
   gpc1_1 gpc229 (
      {stage0_14[46]},
      {stage1_14[23]}
   );
   gpc1_1 gpc230 (
      {stage0_14[47]},
      {stage1_14[24]}
   );
   gpc1_1 gpc231 (
      {stage0_14[48]},
      {stage1_14[25]}
   );
   gpc1_1 gpc232 (
      {stage0_14[49]},
      {stage1_14[26]}
   );
   gpc1_1 gpc233 (
      {stage0_14[50]},
      {stage1_14[27]}
   );
   gpc1_1 gpc234 (
      {stage0_14[51]},
      {stage1_14[28]}
   );
   gpc1_1 gpc235 (
      {stage0_14[52]},
      {stage1_14[29]}
   );
   gpc1_1 gpc236 (
      {stage0_14[53]},
      {stage1_14[30]}
   );
   gpc1_1 gpc237 (
      {stage0_15[44]},
      {stage1_15[18]}
   );
   gpc1_1 gpc238 (
      {stage0_15[45]},
      {stage1_15[19]}
   );
   gpc1_1 gpc239 (
      {stage0_15[46]},
      {stage1_15[20]}
   );
   gpc1_1 gpc240 (
      {stage0_15[47]},
      {stage1_15[21]}
   );
   gpc1_1 gpc241 (
      {stage0_15[48]},
      {stage1_15[22]}
   );
   gpc1_1 gpc242 (
      {stage0_15[49]},
      {stage1_15[23]}
   );
   gpc1_1 gpc243 (
      {stage0_15[50]},
      {stage1_15[24]}
   );
   gpc1_1 gpc244 (
      {stage0_15[51]},
      {stage1_15[25]}
   );
   gpc1_1 gpc245 (
      {stage0_15[52]},
      {stage1_15[26]}
   );
   gpc1_1 gpc246 (
      {stage0_15[53]},
      {stage1_15[27]}
   );
   gpc1_1 gpc247 (
      {stage0_16[49]},
      {stage1_16[20]}
   );
   gpc1_1 gpc248 (
      {stage0_16[50]},
      {stage1_16[21]}
   );
   gpc1_1 gpc249 (
      {stage0_16[51]},
      {stage1_16[22]}
   );
   gpc1_1 gpc250 (
      {stage0_16[52]},
      {stage1_16[23]}
   );
   gpc1_1 gpc251 (
      {stage0_16[53]},
      {stage1_16[24]}
   );
   gpc1_1 gpc252 (
      {stage0_18[42]},
      {stage1_18[18]}
   );
   gpc1_1 gpc253 (
      {stage0_18[43]},
      {stage1_18[19]}
   );
   gpc1_1 gpc254 (
      {stage0_18[44]},
      {stage1_18[20]}
   );
   gpc1_1 gpc255 (
      {stage0_18[45]},
      {stage1_18[21]}
   );
   gpc1_1 gpc256 (
      {stage0_18[46]},
      {stage1_18[22]}
   );
   gpc1_1 gpc257 (
      {stage0_18[47]},
      {stage1_18[23]}
   );
   gpc1_1 gpc258 (
      {stage0_18[48]},
      {stage1_18[24]}
   );
   gpc1_1 gpc259 (
      {stage0_18[49]},
      {stage1_18[25]}
   );
   gpc1_1 gpc260 (
      {stage0_18[50]},
      {stage1_18[26]}
   );
   gpc1_1 gpc261 (
      {stage0_18[51]},
      {stage1_18[27]}
   );
   gpc1_1 gpc262 (
      {stage0_18[52]},
      {stage1_18[28]}
   );
   gpc1_1 gpc263 (
      {stage0_18[53]},
      {stage1_18[29]}
   );
   gpc1_1 gpc264 (
      {stage0_19[40]},
      {stage1_19[18]}
   );
   gpc1_1 gpc265 (
      {stage0_19[41]},
      {stage1_19[19]}
   );
   gpc1_1 gpc266 (
      {stage0_19[42]},
      {stage1_19[20]}
   );
   gpc1_1 gpc267 (
      {stage0_19[43]},
      {stage1_19[21]}
   );
   gpc1_1 gpc268 (
      {stage0_19[44]},
      {stage1_19[22]}
   );
   gpc1_1 gpc269 (
      {stage0_19[45]},
      {stage1_19[23]}
   );
   gpc1_1 gpc270 (
      {stage0_19[46]},
      {stage1_19[24]}
   );
   gpc1_1 gpc271 (
      {stage0_19[47]},
      {stage1_19[25]}
   );
   gpc1_1 gpc272 (
      {stage0_19[48]},
      {stage1_19[26]}
   );
   gpc1_1 gpc273 (
      {stage0_19[49]},
      {stage1_19[27]}
   );
   gpc1_1 gpc274 (
      {stage0_19[50]},
      {stage1_19[28]}
   );
   gpc1_1 gpc275 (
      {stage0_19[51]},
      {stage1_19[29]}
   );
   gpc1_1 gpc276 (
      {stage0_19[52]},
      {stage1_19[30]}
   );
   gpc1_1 gpc277 (
      {stage0_19[53]},
      {stage1_19[31]}
   );
   gpc1_1 gpc278 (
      {stage0_20[53]},
      {stage1_20[22]}
   );
   gpc1_1 gpc279 (
      {stage0_21[45]},
      {stage1_21[21]}
   );
   gpc1_1 gpc280 (
      {stage0_21[46]},
      {stage1_21[22]}
   );
   gpc1_1 gpc281 (
      {stage0_21[47]},
      {stage1_21[23]}
   );
   gpc1_1 gpc282 (
      {stage0_21[48]},
      {stage1_21[24]}
   );
   gpc1_1 gpc283 (
      {stage0_21[49]},
      {stage1_21[25]}
   );
   gpc1_1 gpc284 (
      {stage0_21[50]},
      {stage1_21[26]}
   );
   gpc1_1 gpc285 (
      {stage0_21[51]},
      {stage1_21[27]}
   );
   gpc1_1 gpc286 (
      {stage0_21[52]},
      {stage1_21[28]}
   );
   gpc1_1 gpc287 (
      {stage0_21[53]},
      {stage1_21[29]}
   );
   gpc1_1 gpc288 (
      {stage0_22[48]},
      {stage1_22[16]}
   );
   gpc1_1 gpc289 (
      {stage0_22[49]},
      {stage1_22[17]}
   );
   gpc1_1 gpc290 (
      {stage0_22[50]},
      {stage1_22[18]}
   );
   gpc1_1 gpc291 (
      {stage0_22[51]},
      {stage1_22[19]}
   );
   gpc1_1 gpc292 (
      {stage0_22[52]},
      {stage1_22[20]}
   );
   gpc1_1 gpc293 (
      {stage0_22[53]},
      {stage1_22[21]}
   );
   gpc1_1 gpc294 (
      {stage0_23[42]},
      {stage1_23[17]}
   );
   gpc1_1 gpc295 (
      {stage0_23[43]},
      {stage1_23[18]}
   );
   gpc1_1 gpc296 (
      {stage0_23[44]},
      {stage1_23[19]}
   );
   gpc1_1 gpc297 (
      {stage0_23[45]},
      {stage1_23[20]}
   );
   gpc1_1 gpc298 (
      {stage0_23[46]},
      {stage1_23[21]}
   );
   gpc1_1 gpc299 (
      {stage0_23[47]},
      {stage1_23[22]}
   );
   gpc1_1 gpc300 (
      {stage0_23[48]},
      {stage1_23[23]}
   );
   gpc1_1 gpc301 (
      {stage0_23[49]},
      {stage1_23[24]}
   );
   gpc1_1 gpc302 (
      {stage0_23[50]},
      {stage1_23[25]}
   );
   gpc1_1 gpc303 (
      {stage0_23[51]},
      {stage1_23[26]}
   );
   gpc1_1 gpc304 (
      {stage0_23[52]},
      {stage1_23[27]}
   );
   gpc1_1 gpc305 (
      {stage0_23[53]},
      {stage1_23[28]}
   );
   gpc1_1 gpc306 (
      {stage0_27[48]},
      {stage1_27[19]}
   );
   gpc1_1 gpc307 (
      {stage0_27[49]},
      {stage1_27[20]}
   );
   gpc1_1 gpc308 (
      {stage0_27[50]},
      {stage1_27[21]}
   );
   gpc1_1 gpc309 (
      {stage0_27[51]},
      {stage1_27[22]}
   );
   gpc1_1 gpc310 (
      {stage0_27[52]},
      {stage1_27[23]}
   );
   gpc1_1 gpc311 (
      {stage0_27[53]},
      {stage1_27[24]}
   );
   gpc1_1 gpc312 (
      {stage0_31[48]},
      {stage1_31[18]}
   );
   gpc1_1 gpc313 (
      {stage0_31[49]},
      {stage1_31[19]}
   );
   gpc1_1 gpc314 (
      {stage0_31[50]},
      {stage1_31[20]}
   );
   gpc1_1 gpc315 (
      {stage0_31[51]},
      {stage1_31[21]}
   );
   gpc1_1 gpc316 (
      {stage0_31[52]},
      {stage1_31[22]}
   );
   gpc1_1 gpc317 (
      {stage0_31[53]},
      {stage1_31[23]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc319 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[6]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc320 (
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc321 (
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc615_5 gpc322 (
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage1_4[2]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4],stage2_3[4]}
   );
   gpc606_5 gpc323 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc324 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc325 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[5],stage2_4[7]}
   );
   gpc606_5 gpc326 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[6],stage2_4[8]}
   );
   gpc606_5 gpc327 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[7],stage2_4[9]}
   );
   gpc606_5 gpc328 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[5],stage2_7[8],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc329 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc330 (
      {stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc331 (
      {stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6], stage1_8[7]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[2],stage2_9[3],stage2_8[8]}
   );
   gpc606_5 gpc332 (
      {stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[3],stage2_9[4],stage2_8[9]}
   );
   gpc606_5 gpc333 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[4],stage2_10[4],stage2_9[5],stage2_8[10]}
   );
   gpc606_5 gpc334 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[3],stage2_11[5],stage2_10[5],stage2_9[6]}
   );
   gpc606_5 gpc335 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[4],stage2_11[6],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc336 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[5],stage2_11[7],stage2_10[7],stage2_9[8]}
   );
   gpc606_5 gpc337 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[6],stage2_11[8],stage2_10[8],stage2_9[9]}
   );
   gpc615_5 gpc338 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[4],stage2_12[7],stage2_11[9]}
   );
   gpc606_5 gpc339 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[5],stage2_12[8]}
   );
   gpc606_5 gpc340 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[6],stage2_12[9]}
   );
   gpc606_5 gpc341 (
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[7],stage2_12[10]}
   );
   gpc606_5 gpc342 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[4],stage2_13[8]}
   );
   gpc606_5 gpc343 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[5],stage2_13[9]}
   );
   gpc606_5 gpc344 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[6],stage2_13[10]}
   );
   gpc1163_5 gpc345 (
      {stage1_14[18], stage1_14[19], stage1_14[20]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[7]}
   );
   gpc615_5 gpc346 (
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage1_15[24]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[1],stage2_17[4],stage2_16[7],stage2_15[8],stage2_14[8]}
   );
   gpc615_5 gpc347 (
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage1_15[25]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[2],stage2_17[5],stage2_16[8],stage2_15[9],stage2_14[9]}
   );
   gpc606_5 gpc348 (
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[3],stage2_17[6],stage2_16[9]}
   );
   gpc606_5 gpc349 (
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[4],stage2_17[7],stage2_16[10]}
   );
   gpc606_5 gpc350 (
      {stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[5],stage2_17[8]}
   );
   gpc606_5 gpc351 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[6],stage2_17[9]}
   );
   gpc606_5 gpc352 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[7],stage2_17[10]}
   );
   gpc615_5 gpc353 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16]},
      {stage1_19[18]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[8]}
   );
   gpc615_5 gpc354 (
      {stage1_18[17], stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21]},
      {stage1_19[19]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[9]}
   );
   gpc615_5 gpc355 (
      {stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26]},
      {stage1_19[20]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[10]}
   );
   gpc606_5 gpc356 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25], stage1_19[26]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[6],stage2_20[8],stage2_19[8]}
   );
   gpc606_5 gpc357 (
      {stage1_19[27], stage1_19[28], stage1_19[29], stage1_19[30], stage1_19[31], 1'b0},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[7],stage2_20[9],stage2_19[9]}
   );
   gpc606_5 gpc358 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], 1'b0},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[2],stage2_22[5],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc359 (
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[3],stage2_22[6],stage2_21[9]}
   );
   gpc606_5 gpc360 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[4],stage2_22[7],stage2_21[10]}
   );
   gpc606_5 gpc361 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[5],stage2_22[8],stage2_21[11]}
   );
   gpc615_5 gpc362 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10]},
      {stage1_23[18]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[3],stage2_24[4],stage2_23[6],stage2_22[9]}
   );
   gpc615_5 gpc363 (
      {stage1_22[11], stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15]},
      {stage1_23[19]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[4],stage2_24[5],stage2_23[7],stage2_22[10]}
   );
   gpc1415_5 gpc364 (
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4]},
      {stage1_26[0]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3]},
      {stage1_28[0]},
      {stage2_29[0],stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[5]}
   );
   gpc615_5 gpc365 (
      {stage1_25[5], stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9]},
      {stage1_26[1]},
      {stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage2_29[1],stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[6]}
   );
   gpc615_5 gpc366 (
      {stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13], stage1_25[14]},
      {stage1_26[2]},
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15]},
      {stage2_29[2],stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[7]}
   );
   gpc615_5 gpc367 (
      {stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18], stage1_25[19]},
      {stage1_26[3]},
      {stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21]},
      {stage2_29[3],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[8]}
   );
   gpc615_5 gpc368 (
      {stage1_26[4], stage1_26[5], stage1_26[6], stage1_26[7], stage1_26[8]},
      {stage1_27[22]},
      {stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5], stage1_28[6]},
      {stage2_30[0],stage2_29[4],stage2_28[4],stage2_27[4],stage2_26[6]}
   );
   gpc615_5 gpc369 (
      {stage1_26[9], stage1_26[10], stage1_26[11], stage1_26[12], stage1_26[13]},
      {stage1_27[23]},
      {stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12]},
      {stage2_30[1],stage2_29[5],stage2_28[5],stage2_27[5],stage2_26[7]}
   );
   gpc615_5 gpc370 (
      {stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17], 1'b0},
      {stage1_27[24]},
      {stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18]},
      {stage2_30[2],stage2_29[6],stage2_28[6],stage2_27[6],stage2_26[8]}
   );
   gpc2135_5 gpc371 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage1_32[0], stage1_32[1]},
      {stage2_33[0],stage2_32[0],stage2_31[0],stage2_30[3],stage2_29[7]}
   );
   gpc1406_5 gpc372 (
      {stage1_29[5], stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10]},
      {stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4]},
      {stage1_32[2]},
      {stage2_33[1],stage2_32[1],stage2_31[1],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc373 (
      {stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10]},
      {stage2_33[2],stage2_32[2],stage2_31[2],stage2_30[5],stage2_29[9]}
   );
   gpc606_5 gpc374 (
      {stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8]},
      {stage2_34[0],stage2_33[3],stage2_32[3],stage2_31[3],stage2_30[6]}
   );
   gpc606_5 gpc375 (
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14]},
      {stage2_34[1],stage2_33[4],stage2_32[4],stage2_31[4],stage2_30[7]}
   );
   gpc615_5 gpc376 (
      {stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_32[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[5],stage2_32[5],stage2_31[5]}
   );
   gpc615_5 gpc377 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20]},
      {stage1_32[16]},
      {stage1_33[6], stage1_33[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_35[1],stage2_34[3],stage2_33[6],stage2_32[6],stage2_31[6]}
   );
   gpc1_1 gpc378 (
      {stage1_0[8]},
      {stage2_0[2]}
   );
   gpc1_1 gpc379 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc380 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc381 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc382 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc383 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc384 (
      {stage1_0[14]},
      {stage2_0[8]}
   );
   gpc1_1 gpc385 (
      {stage1_0[15]},
      {stage2_0[9]}
   );
   gpc1_1 gpc386 (
      {stage1_1[7]},
      {stage2_1[2]}
   );
   gpc1_1 gpc387 (
      {stage1_1[8]},
      {stage2_1[3]}
   );
   gpc1_1 gpc388 (
      {stage1_1[9]},
      {stage2_1[4]}
   );
   gpc1_1 gpc389 (
      {stage1_1[10]},
      {stage2_1[5]}
   );
   gpc1_1 gpc390 (
      {stage1_1[11]},
      {stage2_1[6]}
   );
   gpc1_1 gpc391 (
      {stage1_1[12]},
      {stage2_1[7]}
   );
   gpc1_1 gpc392 (
      {stage1_1[13]},
      {stage2_1[8]}
   );
   gpc1_1 gpc393 (
      {stage1_1[14]},
      {stage2_1[9]}
   );
   gpc1_1 gpc394 (
      {stage1_1[15]},
      {stage2_1[10]}
   );
   gpc1_1 gpc395 (
      {stage1_1[16]},
      {stage2_1[11]}
   );
   gpc1_1 gpc396 (
      {stage1_2[7]},
      {stage2_2[2]}
   );
   gpc1_1 gpc397 (
      {stage1_2[8]},
      {stage2_2[3]}
   );
   gpc1_1 gpc398 (
      {stage1_2[9]},
      {stage2_2[4]}
   );
   gpc1_1 gpc399 (
      {stage1_2[10]},
      {stage2_2[5]}
   );
   gpc1_1 gpc400 (
      {stage1_2[11]},
      {stage2_2[6]}
   );
   gpc1_1 gpc401 (
      {stage1_2[12]},
      {stage2_2[7]}
   );
   gpc1_1 gpc402 (
      {stage1_2[13]},
      {stage2_2[8]}
   );
   gpc1_1 gpc403 (
      {stage1_2[14]},
      {stage2_2[9]}
   );
   gpc1_1 gpc404 (
      {stage1_2[15]},
      {stage2_2[10]}
   );
   gpc1_1 gpc405 (
      {stage1_2[16]},
      {stage2_2[11]}
   );
   gpc1_1 gpc406 (
      {stage1_2[17]},
      {stage2_2[12]}
   );
   gpc1_1 gpc407 (
      {stage1_2[18]},
      {stage2_2[13]}
   );
   gpc1_1 gpc408 (
      {stage1_2[19]},
      {stage2_2[14]}
   );
   gpc1_1 gpc409 (
      {stage1_2[20]},
      {stage2_2[15]}
   );
   gpc1_1 gpc410 (
      {stage1_2[21]},
      {stage2_2[16]}
   );
   gpc1_1 gpc411 (
      {stage1_3[16]},
      {stage2_3[5]}
   );
   gpc1_1 gpc412 (
      {stage1_3[17]},
      {stage2_3[6]}
   );
   gpc1_1 gpc413 (
      {stage1_3[18]},
      {stage2_3[7]}
   );
   gpc1_1 gpc414 (
      {stage1_3[19]},
      {stage2_3[8]}
   );
   gpc1_1 gpc415 (
      {stage1_3[20]},
      {stage2_3[9]}
   );
   gpc1_1 gpc416 (
      {stage1_3[21]},
      {stage2_3[10]}
   );
   gpc1_1 gpc417 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc418 (
      {stage1_5[25]},
      {stage2_5[10]}
   );
   gpc1_1 gpc419 (
      {stage1_5[26]},
      {stage2_5[11]}
   );
   gpc1_1 gpc420 (
      {stage1_6[30]},
      {stage2_6[9]}
   );
   gpc1_1 gpc421 (
      {stage1_6[31]},
      {stage2_6[10]}
   );
   gpc1_1 gpc422 (
      {stage1_6[32]},
      {stage2_6[11]}
   );
   gpc1_1 gpc423 (
      {stage1_7[16]},
      {stage2_7[11]}
   );
   gpc1_1 gpc424 (
      {stage1_7[17]},
      {stage2_7[12]}
   );
   gpc1_1 gpc425 (
      {stage1_7[18]},
      {stage2_7[13]}
   );
   gpc1_1 gpc426 (
      {stage1_7[19]},
      {stage2_7[14]}
   );
   gpc1_1 gpc427 (
      {stage1_7[20]},
      {stage2_7[15]}
   );
   gpc1_1 gpc428 (
      {stage1_8[20]},
      {stage2_8[11]}
   );
   gpc1_1 gpc429 (
      {stage1_8[21]},
      {stage2_8[12]}
   );
   gpc1_1 gpc430 (
      {stage1_8[22]},
      {stage2_8[13]}
   );
   gpc1_1 gpc431 (
      {stage1_8[23]},
      {stage2_8[14]}
   );
   gpc1_1 gpc432 (
      {stage1_8[24]},
      {stage2_8[15]}
   );
   gpc1_1 gpc433 (
      {stage1_8[25]},
      {stage2_8[16]}
   );
   gpc1_1 gpc434 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc435 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc436 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc437 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc438 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc439 (
      {stage1_13[24]},
      {stage2_13[11]}
   );
   gpc1_1 gpc440 (
      {stage1_13[25]},
      {stage2_13[12]}
   );
   gpc1_1 gpc441 (
      {stage1_13[26]},
      {stage2_13[13]}
   );
   gpc1_1 gpc442 (
      {stage1_13[27]},
      {stage2_13[14]}
   );
   gpc1_1 gpc443 (
      {stage1_13[28]},
      {stage2_13[15]}
   );
   gpc1_1 gpc444 (
      {stage1_13[29]},
      {stage2_13[16]}
   );
   gpc1_1 gpc445 (
      {stage1_13[30]},
      {stage2_13[17]}
   );
   gpc1_1 gpc446 (
      {stage1_13[31]},
      {stage2_13[18]}
   );
   gpc1_1 gpc447 (
      {stage1_15[26]},
      {stage2_15[10]}
   );
   gpc1_1 gpc448 (
      {stage1_15[27]},
      {stage2_15[11]}
   );
   gpc1_1 gpc449 (
      {stage1_17[19]},
      {stage2_17[11]}
   );
   gpc1_1 gpc450 (
      {stage1_18[27]},
      {stage2_18[11]}
   );
   gpc1_1 gpc451 (
      {stage1_18[28]},
      {stage2_18[12]}
   );
   gpc1_1 gpc452 (
      {stage1_18[29]},
      {stage2_18[13]}
   );
   gpc1_1 gpc453 (
      {stage1_22[16]},
      {stage2_22[11]}
   );
   gpc1_1 gpc454 (
      {stage1_22[17]},
      {stage2_22[12]}
   );
   gpc1_1 gpc455 (
      {stage1_22[18]},
      {stage2_22[13]}
   );
   gpc1_1 gpc456 (
      {stage1_22[19]},
      {stage2_22[14]}
   );
   gpc1_1 gpc457 (
      {stage1_22[20]},
      {stage2_22[15]}
   );
   gpc1_1 gpc458 (
      {stage1_22[21]},
      {stage2_22[16]}
   );
   gpc1_1 gpc459 (
      {stage1_23[20]},
      {stage2_23[8]}
   );
   gpc1_1 gpc460 (
      {stage1_23[21]},
      {stage2_23[9]}
   );
   gpc1_1 gpc461 (
      {stage1_23[22]},
      {stage2_23[10]}
   );
   gpc1_1 gpc462 (
      {stage1_23[23]},
      {stage2_23[11]}
   );
   gpc1_1 gpc463 (
      {stage1_23[24]},
      {stage2_23[12]}
   );
   gpc1_1 gpc464 (
      {stage1_23[25]},
      {stage2_23[13]}
   );
   gpc1_1 gpc465 (
      {stage1_23[26]},
      {stage2_23[14]}
   );
   gpc1_1 gpc466 (
      {stage1_23[27]},
      {stage2_23[15]}
   );
   gpc1_1 gpc467 (
      {stage1_23[28]},
      {stage2_23[16]}
   );
   gpc1_1 gpc468 (
      {stage1_24[12]},
      {stage2_24[6]}
   );
   gpc1_1 gpc469 (
      {stage1_24[13]},
      {stage2_24[7]}
   );
   gpc1_1 gpc470 (
      {stage1_24[14]},
      {stage2_24[8]}
   );
   gpc1_1 gpc471 (
      {stage1_24[15]},
      {stage2_24[9]}
   );
   gpc1_1 gpc472 (
      {stage1_24[16]},
      {stage2_24[10]}
   );
   gpc1_1 gpc473 (
      {stage1_24[17]},
      {stage2_24[11]}
   );
   gpc1_1 gpc474 (
      {stage1_24[18]},
      {stage2_24[12]}
   );
   gpc1_1 gpc475 (
      {stage1_24[19]},
      {stage2_24[13]}
   );
   gpc1_1 gpc476 (
      {stage1_24[20]},
      {stage2_24[14]}
   );
   gpc1_1 gpc477 (
      {stage1_24[21]},
      {stage2_24[15]}
   );
   gpc1_1 gpc478 (
      {stage1_24[22]},
      {stage2_24[16]}
   );
   gpc1_1 gpc479 (
      {stage1_24[23]},
      {stage2_24[17]}
   );
   gpc1_1 gpc480 (
      {stage1_25[20]},
      {stage2_25[9]}
   );
   gpc1_1 gpc481 (
      {stage1_25[21]},
      {stage2_25[10]}
   );
   gpc1_1 gpc482 (
      {stage1_25[22]},
      {stage2_25[11]}
   );
   gpc1_1 gpc483 (
      {stage1_28[19]},
      {stage2_28[7]}
   );
   gpc1_1 gpc484 (
      {stage1_28[20]},
      {stage2_28[8]}
   );
   gpc1_1 gpc485 (
      {stage1_28[21]},
      {stage2_28[9]}
   );
   gpc1_1 gpc486 (
      {stage1_28[22]},
      {stage2_28[10]}
   );
   gpc1_1 gpc487 (
      {stage1_28[23]},
      {stage2_28[11]}
   );
   gpc1_1 gpc488 (
      {stage1_28[24]},
      {stage2_28[12]}
   );
   gpc1_1 gpc489 (
      {stage1_28[25]},
      {stage2_28[13]}
   );
   gpc1_1 gpc490 (
      {stage1_29[17]},
      {stage2_29[10]}
   );
   gpc1_1 gpc491 (
      {stage1_29[18]},
      {stage2_29[11]}
   );
   gpc1_1 gpc492 (
      {stage1_29[19]},
      {stage2_29[12]}
   );
   gpc1_1 gpc493 (
      {stage1_29[20]},
      {stage2_29[13]}
   );
   gpc1_1 gpc494 (
      {stage1_29[21]},
      {stage2_29[14]}
   );
   gpc1_1 gpc495 (
      {stage1_29[22]},
      {stage2_29[15]}
   );
   gpc1_1 gpc496 (
      {stage1_29[23]},
      {stage2_29[16]}
   );
   gpc1_1 gpc497 (
      {stage1_29[24]},
      {stage2_29[17]}
   );
   gpc1_1 gpc498 (
      {stage1_30[15]},
      {stage2_30[8]}
   );
   gpc1_1 gpc499 (
      {stage1_30[16]},
      {stage2_30[9]}
   );
   gpc1_1 gpc500 (
      {stage1_30[17]},
      {stage2_30[10]}
   );
   gpc1_1 gpc501 (
      {stage1_31[21]},
      {stage2_31[7]}
   );
   gpc1_1 gpc502 (
      {stage1_31[22]},
      {stage2_31[8]}
   );
   gpc1_1 gpc503 (
      {stage1_31[23]},
      {stage2_31[9]}
   );
   gpc615_5 gpc504 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc505 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc506 (
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc507 (
      {stage2_4[6], stage2_4[7], stage2_4[8]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0]},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc606_5 gpc508 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[2]}
   );
   gpc606_5 gpc509 (
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[2],stage3_7[2],stage3_6[3]}
   );
   gpc606_5 gpc510 (
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], 1'b0},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[3],stage3_7[3],stage3_6[4]}
   );
   gpc615_5 gpc511 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[3],stage3_8[4],stage3_7[4]}
   );
   gpc606_5 gpc512 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[3]}
   );
   gpc615_5 gpc513 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[1],stage3_11[2]}
   );
   gpc615_5 gpc514 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage2_12[7]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[2],stage3_11[3]}
   );
   gpc606_5 gpc515 (
      {stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[3],stage3_13[3],stage3_12[3]}
   );
   gpc135_4 gpc516 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16]},
      {stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage2_15[0]},
      {stage3_16[1],stage3_15[3],stage3_14[4],stage3_13[4]}
   );
   gpc606_5 gpc517 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[4]}
   );
   gpc615_5 gpc518 (
      {stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[1],stage3_17[1],stage3_16[3],stage3_15[5]}
   );
   gpc606_5 gpc519 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[2],stage3_17[2],stage3_16[4]}
   );
   gpc1343_5 gpc520 (
      {stage2_18[6], stage2_18[7], stage2_18[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[3]}
   );
   gpc1343_5 gpc521 (
      {stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[4]}
   );
   gpc606_5 gpc522 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[2]}
   );
   gpc615_5 gpc523 (
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4]},
      {stage2_23[6]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3]}
   );
   gpc615_5 gpc524 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9]},
      {stage2_23[7]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4]}
   );
   gpc615_5 gpc525 (
      {stage2_22[10], stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14]},
      {stage2_23[8]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5]}
   );
   gpc606_5 gpc526 (
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[3],stage3_25[4],stage3_24[4],stage3_23[4]}
   );
   gpc606_5 gpc527 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[1],stage3_26[4],stage3_25[5]}
   );
   gpc1415_5 gpc528 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4]},
      {stage2_27[6]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[1],stage3_28[1],stage3_27[2],stage3_26[5]}
   );
   gpc615_5 gpc529 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[1]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[2],stage3_28[2]}
   );
   gpc615_5 gpc530 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[2]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], 1'b0},
      {stage3_32[1],stage3_31[1],stage3_30[2],stage3_29[3],stage3_28[3]}
   );
   gpc606_5 gpc531 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[2],stage3_31[2]}
   );
   gpc117_4 gpc532 (
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5], stage2_32[6]},
      {stage2_33[6]},
      {stage2_34[0]},
      {stage3_35[1],stage3_34[1],stage3_33[1],stage3_32[3]}
   );
   gpc1_1 gpc533 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc534 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc535 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc536 (
      {stage2_1[5]},
      {stage3_1[5]}
   );
   gpc1_1 gpc537 (
      {stage2_1[6]},
      {stage3_1[6]}
   );
   gpc1_1 gpc538 (
      {stage2_1[7]},
      {stage3_1[7]}
   );
   gpc1_1 gpc539 (
      {stage2_1[8]},
      {stage3_1[8]}
   );
   gpc1_1 gpc540 (
      {stage2_1[9]},
      {stage3_1[9]}
   );
   gpc1_1 gpc541 (
      {stage2_1[10]},
      {stage3_1[10]}
   );
   gpc1_1 gpc542 (
      {stage2_1[11]},
      {stage3_1[11]}
   );
   gpc1_1 gpc543 (
      {stage2_3[1]},
      {stage3_3[3]}
   );
   gpc1_1 gpc544 (
      {stage2_3[2]},
      {stage3_3[4]}
   );
   gpc1_1 gpc545 (
      {stage2_3[3]},
      {stage3_3[5]}
   );
   gpc1_1 gpc546 (
      {stage2_3[4]},
      {stage3_3[6]}
   );
   gpc1_1 gpc547 (
      {stage2_3[5]},
      {stage3_3[7]}
   );
   gpc1_1 gpc548 (
      {stage2_3[6]},
      {stage3_3[8]}
   );
   gpc1_1 gpc549 (
      {stage2_3[7]},
      {stage3_3[9]}
   );
   gpc1_1 gpc550 (
      {stage2_3[8]},
      {stage3_3[10]}
   );
   gpc1_1 gpc551 (
      {stage2_3[9]},
      {stage3_3[11]}
   );
   gpc1_1 gpc552 (
      {stage2_3[10]},
      {stage3_3[12]}
   );
   gpc1_1 gpc553 (
      {stage2_4[9]},
      {stage3_4[4]}
   );
   gpc1_1 gpc554 (
      {stage2_7[12]},
      {stage3_7[5]}
   );
   gpc1_1 gpc555 (
      {stage2_7[13]},
      {stage3_7[6]}
   );
   gpc1_1 gpc556 (
      {stage2_7[14]},
      {stage3_7[7]}
   );
   gpc1_1 gpc557 (
      {stage2_7[15]},
      {stage3_7[8]}
   );
   gpc1_1 gpc558 (
      {stage2_8[13]},
      {stage3_8[5]}
   );
   gpc1_1 gpc559 (
      {stage2_8[14]},
      {stage3_8[6]}
   );
   gpc1_1 gpc560 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc561 (
      {stage2_8[16]},
      {stage3_8[8]}
   );
   gpc1_1 gpc562 (
      {stage2_9[6]},
      {stage3_9[4]}
   );
   gpc1_1 gpc563 (
      {stage2_9[7]},
      {stage3_9[5]}
   );
   gpc1_1 gpc564 (
      {stage2_9[8]},
      {stage3_9[6]}
   );
   gpc1_1 gpc565 (
      {stage2_9[9]},
      {stage3_9[7]}
   );
   gpc1_1 gpc566 (
      {stage2_10[6]},
      {stage3_10[4]}
   );
   gpc1_1 gpc567 (
      {stage2_10[7]},
      {stage3_10[5]}
   );
   gpc1_1 gpc568 (
      {stage2_10[8]},
      {stage3_10[6]}
   );
   gpc1_1 gpc569 (
      {stage2_12[14]},
      {stage3_12[4]}
   );
   gpc1_1 gpc570 (
      {stage2_12[15]},
      {stage3_12[5]}
   );
   gpc1_1 gpc571 (
      {stage2_13[17]},
      {stage3_13[5]}
   );
   gpc1_1 gpc572 (
      {stage2_13[18]},
      {stage3_13[6]}
   );
   gpc1_1 gpc573 (
      {stage2_14[9]},
      {stage3_14[5]}
   );
   gpc1_1 gpc574 (
      {stage2_16[7]},
      {stage3_16[5]}
   );
   gpc1_1 gpc575 (
      {stage2_16[8]},
      {stage3_16[6]}
   );
   gpc1_1 gpc576 (
      {stage2_16[9]},
      {stage3_16[7]}
   );
   gpc1_1 gpc577 (
      {stage2_16[10]},
      {stage3_16[8]}
   );
   gpc1_1 gpc578 (
      {stage2_18[12]},
      {stage3_18[5]}
   );
   gpc1_1 gpc579 (
      {stage2_18[13]},
      {stage3_18[6]}
   );
   gpc1_1 gpc580 (
      {stage2_19[8]},
      {stage3_19[5]}
   );
   gpc1_1 gpc581 (
      {stage2_19[9]},
      {stage3_19[6]}
   );
   gpc1_1 gpc582 (
      {stage2_20[6]},
      {stage3_20[3]}
   );
   gpc1_1 gpc583 (
      {stage2_20[7]},
      {stage3_20[4]}
   );
   gpc1_1 gpc584 (
      {stage2_20[8]},
      {stage3_20[5]}
   );
   gpc1_1 gpc585 (
      {stage2_20[9]},
      {stage3_20[6]}
   );
   gpc1_1 gpc586 (
      {stage2_20[10]},
      {stage3_20[7]}
   );
   gpc1_1 gpc587 (
      {stage2_21[8]},
      {stage3_21[3]}
   );
   gpc1_1 gpc588 (
      {stage2_21[9]},
      {stage3_21[4]}
   );
   gpc1_1 gpc589 (
      {stage2_21[10]},
      {stage3_21[5]}
   );
   gpc1_1 gpc590 (
      {stage2_21[11]},
      {stage3_21[6]}
   );
   gpc1_1 gpc591 (
      {stage2_22[15]},
      {stage3_22[6]}
   );
   gpc1_1 gpc592 (
      {stage2_22[16]},
      {stage3_22[7]}
   );
   gpc1_1 gpc593 (
      {stage2_23[15]},
      {stage3_23[5]}
   );
   gpc1_1 gpc594 (
      {stage2_23[16]},
      {stage3_23[6]}
   );
   gpc1_1 gpc595 (
      {stage2_26[5]},
      {stage3_26[6]}
   );
   gpc1_1 gpc596 (
      {stage2_26[6]},
      {stage3_26[7]}
   );
   gpc1_1 gpc597 (
      {stage2_26[7]},
      {stage3_26[8]}
   );
   gpc1_1 gpc598 (
      {stage2_26[8]},
      {stage3_26[9]}
   );
   gpc1_1 gpc599 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc600 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc601 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc602 (
      {stage2_29[6]},
      {stage3_29[7]}
   );
   gpc1_1 gpc603 (
      {stage2_29[7]},
      {stage3_29[8]}
   );
   gpc1_1 gpc604 (
      {stage2_29[8]},
      {stage3_29[9]}
   );
   gpc1_1 gpc605 (
      {stage2_29[9]},
      {stage3_29[10]}
   );
   gpc1_1 gpc606 (
      {stage2_29[10]},
      {stage3_29[11]}
   );
   gpc1_1 gpc607 (
      {stage2_29[11]},
      {stage3_29[12]}
   );
   gpc1_1 gpc608 (
      {stage2_29[12]},
      {stage3_29[13]}
   );
   gpc1_1 gpc609 (
      {stage2_29[13]},
      {stage3_29[14]}
   );
   gpc1_1 gpc610 (
      {stage2_29[14]},
      {stage3_29[15]}
   );
   gpc1_1 gpc611 (
      {stage2_29[15]},
      {stage3_29[16]}
   );
   gpc1_1 gpc612 (
      {stage2_29[16]},
      {stage3_29[17]}
   );
   gpc1_1 gpc613 (
      {stage2_29[17]},
      {stage3_29[18]}
   );
   gpc1_1 gpc614 (
      {stage2_31[6]},
      {stage3_31[3]}
   );
   gpc1_1 gpc615 (
      {stage2_31[7]},
      {stage3_31[4]}
   );
   gpc1_1 gpc616 (
      {stage2_31[8]},
      {stage3_31[5]}
   );
   gpc1_1 gpc617 (
      {stage2_31[9]},
      {stage3_31[6]}
   );
   gpc1_1 gpc618 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1_1 gpc619 (
      {stage2_34[2]},
      {stage3_34[3]}
   );
   gpc1_1 gpc620 (
      {stage2_34[3]},
      {stage3_34[4]}
   );
   gpc1_1 gpc621 (
      {stage2_35[0]},
      {stage3_35[2]}
   );
   gpc1_1 gpc622 (
      {stage2_35[1]},
      {stage3_35[3]}
   );
   gpc615_5 gpc623 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4]},
      {stage3_2[0]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc624 (
      {stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9]},
      {stage3_2[1]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc2135_5 gpc625 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[2]}
   );
   gpc623_5 gpc626 (
      {stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1]}
   );
   gpc615_5 gpc627 (
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[2]}
   );
   gpc615_5 gpc628 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[2]}
   );
   gpc623_5 gpc629 (
      {stage3_11[1], stage3_11[2], stage3_11[3]},
      {1'b0, 1'b0},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1],stage4_11[2]}
   );
   gpc1406_5 gpc630 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[2]}
   );
   gpc215_4 gpc631 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[4]},
      {stage3_17[1], stage3_17[2]},
      {stage4_18[1],stage4_17[1],stage4_16[1],stage4_15[2]}
   );
   gpc606_5 gpc632 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[2]}
   );
   gpc117_4 gpc633 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_20[6]},
      {stage3_21[0]},
      {stage4_22[1],stage4_21[1],stage4_20[1],stage4_19[1]}
   );
   gpc606_5 gpc634 (
      {stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[0],stage4_23[0],stage4_22[2],stage4_21[2]}
   );
   gpc606_5 gpc635 (
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], 1'b0},
      {stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[1],stage4_22[3]}
   );
   gpc1343_5 gpc636 (
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3]},
      {stage3_27[0], stage3_27[1], stage3_27[2]},
      {stage3_28[0]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[1],stage4_25[2]}
   );
   gpc135_4 gpc637 (
      {stage3_28[1], stage3_28[2], stage3_28[3], 1'b0, 1'b0},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[1]}
   );
   gpc207_4 gpc638 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[2]}
   );
   gpc207_4 gpc639 (
      {stage3_29[10], stage3_29[11], stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc623_5 gpc640 (
      {stage3_32[0], stage3_32[1], stage3_32[2]},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], 1'b0},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[2]}
   );
   gpc215_4 gpc641 (
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], 1'b0},
      {1'b0},
      {1'b0, 1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[1]}
   );
   gpc1_1 gpc642 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc643 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc644 (
      {stage3_1[10]},
      {stage4_1[2]}
   );
   gpc1_1 gpc645 (
      {stage3_1[11]},
      {stage4_1[3]}
   );
   gpc1_1 gpc646 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc647 (
      {stage3_3[12]},
      {stage4_3[2]}
   );
   gpc1_1 gpc648 (
      {stage3_6[4]},
      {stage4_6[2]}
   );
   gpc1_1 gpc649 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc650 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc651 (
      {stage3_9[6]},
      {stage4_9[2]}
   );
   gpc1_1 gpc652 (
      {stage3_9[7]},
      {stage4_9[3]}
   );
   gpc1_1 gpc653 (
      {stage3_10[5]},
      {stage4_10[3]}
   );
   gpc1_1 gpc654 (
      {stage3_10[6]},
      {stage4_10[4]}
   );
   gpc1_1 gpc655 (
      {stage3_13[6]},
      {stage4_13[2]}
   );
   gpc1_1 gpc656 (
      {stage3_15[5]},
      {stage4_15[3]}
   );
   gpc1_1 gpc657 (
      {stage3_16[5]},
      {stage4_16[2]}
   );
   gpc1_1 gpc658 (
      {stage3_16[6]},
      {stage4_16[3]}
   );
   gpc1_1 gpc659 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc660 (
      {stage3_16[8]},
      {stage4_16[5]}
   );
   gpc1_1 gpc661 (
      {stage3_18[6]},
      {stage4_18[3]}
   );
   gpc1_1 gpc662 (
      {stage3_20[7]},
      {stage4_20[2]}
   );
   gpc1_1 gpc663 (
      {stage3_22[6]},
      {stage4_22[4]}
   );
   gpc1_1 gpc664 (
      {stage3_22[7]},
      {stage4_22[5]}
   );
   gpc1_1 gpc665 (
      {stage3_23[6]},
      {stage4_23[2]}
   );
   gpc1_1 gpc666 (
      {stage3_25[3]},
      {stage4_25[3]}
   );
   gpc1_1 gpc667 (
      {stage3_25[4]},
      {stage4_25[4]}
   );
   gpc1_1 gpc668 (
      {stage3_25[5]},
      {stage4_25[5]}
   );
   gpc1_1 gpc669 (
      {stage3_26[4]},
      {stage4_26[2]}
   );
   gpc1_1 gpc670 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc671 (
      {stage3_26[6]},
      {stage4_26[4]}
   );
   gpc1_1 gpc672 (
      {stage3_26[7]},
      {stage4_26[5]}
   );
   gpc1_1 gpc673 (
      {stage3_26[8]},
      {stage4_26[6]}
   );
   gpc1_1 gpc674 (
      {stage3_26[9]},
      {stage4_26[7]}
   );
   gpc1_1 gpc675 (
      {stage3_29[17]},
      {stage4_29[4]}
   );
   gpc1_1 gpc676 (
      {stage3_29[18]},
      {stage4_29[5]}
   );
   gpc1_1 gpc677 (
      {stage3_30[1]},
      {stage4_30[3]}
   );
   gpc1_1 gpc678 (
      {stage3_30[2]},
      {stage4_30[4]}
   );
   gpc1_1 gpc679 (
      {stage3_31[4]},
      {stage4_31[3]}
   );
   gpc1_1 gpc680 (
      {stage3_31[5]},
      {stage4_31[4]}
   );
   gpc1_1 gpc681 (
      {stage3_31[6]},
      {stage4_31[5]}
   );
   gpc1_1 gpc682 (
      {stage3_32[3]},
      {stage4_32[3]}
   );
   gpc23_3 gpc683 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc2223_5 gpc684 (
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1]},
      {stage4_5[0], stage4_5[1]},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[1]}
   );
   gpc1343_5 gpc685 (
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1]}
   );
   gpc135_4 gpc686 (
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], 1'b0},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1423_5 gpc687 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc1325_5 gpc688 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0], stage4_17[1]},
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc689 (
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0], stage4_21[1], stage4_21[2], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1]}
   );
   gpc223_4 gpc690 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[1],stage5_23[1],stage5_22[1]}
   );
   gpc2116_5 gpc691 (
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage4_26[0]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1]}
   );
   gpc7_3 gpc692 (
      {stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage5_28[1],stage5_27[1],stage5_26[1]}
   );
   gpc606_5 gpc693 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[0],stage5_29[1]}
   );
   gpc1415_5 gpc694 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4]},
      {1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[1]}
   );
   gpc1_1 gpc695 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc696 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc697 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc698 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc699 (
      {stage4_4[2]},
      {stage5_4[1]}
   );
   gpc1_1 gpc700 (
      {stage4_5[2]},
      {stage5_5[1]}
   );
   gpc1_1 gpc701 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc702 (
      {stage4_8[4]},
      {stage5_8[1]}
   );
   gpc1_1 gpc703 (
      {stage4_9[3]},
      {stage5_9[1]}
   );
   gpc1_1 gpc704 (
      {stage4_12[1]},
      {stage5_12[1]}
   );
   gpc1_1 gpc705 (
      {stage4_14[2]},
      {stage5_14[1]}
   );
   gpc1_1 gpc706 (
      {stage4_18[3]},
      {stage5_18[1]}
   );
   gpc1_1 gpc707 (
      {stage4_19[1]},
      {stage5_19[1]}
   );
   gpc1_1 gpc708 (
      {stage4_34[0]},
      {stage5_34[1]}
   );
   gpc1_1 gpc709 (
      {stage4_35[0]},
      {stage5_35[0]}
   );
   gpc1_1 gpc710 (
      {stage4_35[1]},
      {stage5_35[1]}
   );
   gpc1_1 gpc711 (
      {stage4_36[0]},
      {stage5_36[0]}
   );
   gpc1_1 gpc712 (
      {stage4_36[1]},
      {stage5_36[1]}
   );
   gpc1_1 gpc713 (
      {stage4_37[0]},
      {stage5_37[0]}
   );
endmodule
module rowadder2_1_38(input [37:0] src0, input [37:0] src1, output [38:0] dst0);
    wire [37:0] gene;
    wire [37:0] prop;
    wire [39:0] out;
    wire [39:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[37:36]}),
        .S({2'h0, prop[37:36]})
    );
    assign dst0 = {carryout[37], out[37:0]};
endmodule


module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor2_1_54_32 compressor2_1_54_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h13d9c604479a9e69ad028fbcc64665f48c878a572ad38f57a94fde36fb07634498578cd687fdf960e244f3e5b446040bc5457658748769e6e13fd5d989aa28b4082fc44d0ea416528715ad29add9419013865a034d320535f924f95757f293cf411789c785f048e2c23615b292bb8cd89c1d6976f9610754dc6dbb488be9ae62d726a83f8897e4a29cc5db986fb329c5377912fe939c04d9770c747924853a444c74be241cc4d6961ee937e11705f96ea53d4ded96cd8d20b8722e795d62157b44cfe5b2b784187639b8097f845d5429c67475d651b3275f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h761ab1430226f954b04b49cc519de8d2550594a52844ee00898becabfd34f31712aa6bd455892387a1d01aceedee17e773ee38f41c4b5684bccc19b6084f5cfb30038e153bd6fcf6613f22695d78db3edb15b38d5718820105c02c58dd473ec137b0a8fd1155a7c12d264dbcde17db52b6d08b98ae533c8e86fd30206840d454a5b827e69c8d6340c2984de4c1cbc726c06b792fd7613b94fd4f5680cf7a0bfac06a6b307b2d97a348e09468842afa25ec506646cec34fbb99ddacd533b45cbe5abb093a74c0acfe2ae9fd56f897a7aec52c924b2623c08e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf12a0f1af1b2072413050d7f1b440c5004b8b59caa99050618318cbd5026792fbb8a8c081f8a38d7676c59d721fa795b86a8249742d078fb80c834e9133c5be489ede4d9b4f256999b6e3bf122ff22fb114567c6f1e4c80d6751dfd5ae1df041228bac340f84ffba4f6a42c6148493495c334d5ef99b27fdb6cfc5445eae3d9408313bd75713f298f804b683ed6e7739b31e353b2e0bb442f03ec6334049539c6b79e11d8bc8fe0f2fd1bbea3ee7efddeec5df23131094cabbedb22e5238cf3bf30bcb3537faa27aa0f8fc0677401e194af4a5cecb6fc059;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h13933751f7f23a684eab61a3b81d74805f5940b918a8efbd2f76f959f70cc87f66d4194dd4a5c229df1213494c86b0f85ad5a41a3781dd7d22d941f87bf091528daf0ea3e44e2aa5816f787ddaff637ecdf113e015378b02ff9ebb626967bf68b7a0b22fd76d75e8ddeeafa3a07abdf19fe81aa6b3e2199c58d82c92b140af6cacccb1b4aff0af37e347dcd87dea3d6981f0fa81237b8326524f0809f8ed6c0340e8553f5ea57b77ae86dd173efe80ea22add52462709ebc464a5c156668efc0333fdb1265829481b53be7824a0f6f296a78c264584b40f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd13e5c6c8f671f01c21a1345e7de66698caf97e9413013fc0b3d027863d37ecefc9ec8c655e60e40abcf09f0640f27a6e51f0649a8b126becafd4358bc17b05e52234779b9b5a60befe5015dd72ee255dd28938a684e08261e0f1067ce94ffdecfb21d651a8c5c041704cf2ed19e9fc7bd83d5fbccc5d4310ce513288950524364222facd0308bd6c62a7ff5235a36fd098f4682962beb8eaeabb816e7842f94f8483d0730e8520e6accd4bd7dd251b125829e03068a4a3c5165680f51fe40e11ac5bc48adb79ca13c381028eed59d9908ac353fc0fd0e35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h522b43f9079c8faf44dfbb4d64ed01d608089fa7597124c72dc26743e2eac254024939b0ed665c81652dff54de817129d09fbcaee17a395ad01620459036d5ca426fa57432c449b50e9f73565e394b13d3e4770c66b4bc77b0affe7bc2553b346e873e6a5f4e47c4239f63c7df7b933c3816f9bfdfacfd294cd2f65e43002f9a55078a05a7a0974c9d1d850aaf29d21b616ad7d701fb34d88149b0f6bacec9b43beff08951c8f83eb66ec714ceb4e9ce808162c1a73d8f00da56f27a39b3fc39b702eee15e5ee9a0d899c355dfec88e7dbd0665653a97120;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h37cfb995855a5f9ed10f51e70cdf3d99f464c0542c5f8c39fcfa0c22c16ecddfe0d689a15ae40d939a90ba4ddd1d7525417b5dd9b4ea7b8491d18d7f9607eebc83ee3ea28b6fc6ff2a4056302a55046b6e236e4e63d630bb310d5c3232f37fe5f58b3c3fdc32a9dc708ee2c1f47392998fc93979fbf12da139996f548b7617205a90c66a31f61034171b7898f2f3ba406066f183f10d3c358de976147fc9e8424cc2f618af04a06e24b4cbb426350033efa07c89a69934fd4ceaac57bcf1b0a6e790d36adc0ebc2317a6ac298ad0999f80d63e5cdb1dc511;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3e4b14efec34082c71db327b607497956522dc5a130f73260905fbb4960b01af1dd8226f13b9f2110666c1bba6d2a72bed24c61823cb074b9d566f65c83776744580123e0971dd2b5555434b6fe1ee0dd5c0dd785cc71132ab16cc8118b2bfd2d6b615fd9c03f1975b03d2578b9db04be478b58eb6d0d62367819948b06f9c37f17d774698189ed3ba3b792c6f1263d753f631a3755e2515d06297266c40f70862f73795f8eed98d868b2e2f98eb466d3d5868a83a3b06776ed6112389eabb524223a7704ad9f4280d3b4b7a116fabfde12717214e02068c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h94f3bb36ec06da7aa23098bc47b0eda103936067594f6d12a00d14e40ea1e2e273c8ac82eda0ce532739d6437157ac5567d9f3f3762acdc2b96dd13bbc4dd001565df0ff5ea488cc6764ffb3b9c5b825b6f1d413e010ed2c25add76d7c9ce21ce8e891d699f9aea52bc4197c8bf9c9b599153a2960c526081a79f0dea46cd79d6e17ff8ae3cb0dd3e0f92d2fb35b98e4a3b87308a8d767b5b6dcfb15e679e5fd4768948840f2726a2d6ac3aa0d19aeb4abab83f5c7c0d9109814919fd23086b52ec6ef3341ea382c982294e4e99980008bfadb01e98934a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h22382755f7dbf23439feaa3a385847fd0d5526a9dc19ac8cf4fbc87189dc2d7d7776afc8efe09f7a36e3bf34dcf9a94857fdc15a7a93ef348bb2ff9e751acc599b02e9f4a84cd0671b24ae9bbe9d73105ad4425234ab6371ac37e33b136a81ab105fc23f34c4e14e47bbee31ea0eb31742eadf8007f529682fb8f2cc480584621137b9338326a2133a1943782a34e7d50f9e7ef33e076ea6df937819e151835f72e118ab7584baabc41029feee29d23f7b1cf96f1939fa1017f9e7a5a936d5944348aab33b2e849fced62057887174b62a783342c2296ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'haf14e7f9a1675405fd8f20d9be407558d23056b2bf43a8e3814f550c7b4a254f1b2aa3351dea789bacf76a5b6e6adb16f549ffa4e0d3276e8b13b3d0e46f619b6479a4c7fe05f4abcc4f824188e0da0ddf7fa3dd95c0b2a965bd00c8fc74623d40e197cc5e8e0478fe5f26d6591d195d1fd014867087abf5fc01aff9342a9a17a6522fc3523530d98b5354270881de8fad52f238c9c71136745bcbdd893cc9204cd2d338a0a3f23435b771a318483e833bea9164936fbd73de1bcfecf5078b8e6d28e38006f13f449082bc81b350363499681c1539932a38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcc7fac28817fff1d07bc62970406ff7011885fcf898994d1033d499008386f2a94453e7a4753a002010a76ae8962579cced21689738bb5a02b99f37f91e1196e052a127857cf9d4e1160c3e3c324a756f4b85fe214a097d40926a8baaf0abc62d4e26be29a6c29206c6c031e688a885c81edb8728a645dc4b8e6ea8b4cb2f2416cab523d5dda2d08a224f94c187d4a4dcf4e00d4528f5ca590b6faa3ece9f0d6d900307a3ba69e72febb001078ad51b5a24d5683b51a883f412e5b41802ddc17b1be3ae8ed65b2f8ff565572e5c43f1e3bd43330a20b870;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hab2a6a912058df1a7b38152b9344c6766e50b93acfcfd07a8c0c387141cf6feccf338cc78931aa8af3b840c5ea70b3c592a7e1816776898032ef8fe7042984cef91e757f2aae9596bf27ae74543a00eeb256ead9e7c6588fba7e46df3bb3804ebf53ab06aee2a8047ffc75d47277271b038a29cf5f05ca39a1dd79858c72231862a98f961629ae9c0d25c3a831373b0542e0956239e34ad16886109355f47ecff55fbd4e6c67af1823b456cf998053b632c87f0ba938e3f40e31a98d37312991d55b6048e871128fbc0428f6335300d8040049414eff27f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6b79fad14706d5e7681dd45f20d1217a529e94ff944277382e1b2f3dc8f23483fff3fd4ecb5319e3541fa1fe256e95922081d8e8a0687336eb3879cb922e14732e85d45eb6413651cd83eb61abce13329dbfb60f6c8a1d7979a06124f4f0f50aa459e0c678b79ad9edb577c7e5d8debcf95a3f8906a8b39732bd47e2340f6c1a48ebcf62ff1f0c9a116369f736a9c543a2eef855c523e5da912fba16540692668c86e0b0200d03940295c2880f6320847072eedf059c2dedb2cb3e7d362ef19dfb55cc2766f0a1ebfa199b9d497a927af6d645a02272b400;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he4c441226f50392c30743107697c2e7ca28ea144ba1344a788d352d230e67baef88454164755ad75d23026d7fb96c706301872c3ebf30c92a8d9262e1c2e31700b666aba6d53dbd4bcdd9f5943dd1d780de838b44b7d3eca1dcf8b09af9ab8b2ed034fe9b3793e6dcb622ad126e5b568cc0002b8fba6b7b9946ae6df5573672ca101b1d48d0afe3ee94db6847993256b661067d3e43f2524fa28e9551e0edbe689ae11bff17243e16bcbc204548a787846f119f429f1c7eaac7fae1d2b532d6951fb80d0251e51789f3d4017632f496f82dc9d03bceabca4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h974bbbcaf487c5f4c5d147f05ac9151511f13d75f40ebbbff04c2ad6d0ed069b9536ad29f7ebf5b0c639cb04dfb5d314e9a24ac1164481981e3fe3d69f74f9841ec7703bf81fe65a6aa663c4a89d5960cfa50b7e11734fc391b4f3e5767f249b02174a1c862e49f1f605cd8ed0f0ce7577854c7c14cb10a7a7469fa3d20084dc6dac6bcfbfe55bfd65ffe579270742a467a580f275191a1fdd9571c79e991bd803e95f40e18877058a91fd98f99cd14b0a9f27650e5f86015d3c591c6eb57a7bdb71c2be1feb89bb24fecc10aa22ad9ab7b44851e6338dc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7b536f515bccec85320a244a4d069f54df5ab43cd1ddd86a6910be6a347bc0302020b2c18922ac87ee0cd9c3d4e229051e9bccd23bcbb9e00e1dd447c4939ea92037b72548f42a1c45b4d327ab563045a5e64709ec1db395d3995530f10d8e135bea2078ff2b3bedad5369fe2c32abcfc43f65ec443bf337b9d53b97dbdb4bd87bb09d459d22b5f62d8fed74859df14862d70c05f0119f1214d500f3aab3499c945c2a819d5da2d691ad95763c842716bfc588b84b55c098b384f60ecc2f45969d58659c5742f826cf86f2a50028898616e8fb091e2b754f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3723c48f853b07f2245eb96c5667a3299759404a67340e79684294e4a7ea48d662f0ed8e48baef17f5f00decc8efc12b04ce3d2333931bfa32c20dbfbe1bdc17a3912d12dcc0c5d91333a99920b0905fad656db1cc32f2c95527189274d41b62aa9d7490c2db3c210b49806fda02dd635981a001ae3d2ebb7dc1144f4bfa30492ef46b75d9499171ea0ee40c8d05dbcf8fc25f3e178563261d13ffcd8f257781e6c1194eb866ed24727047dd5416989e3f999fa5e21250985b9b8575a4f18dbb29fac55e2a07208014c3839e4091208dc5797a6b5c457ba5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'habebc7f0d855d03a384651e25fbfb4143094efdcd7fd0fed6fc04228bab11a215bc3761383f26e74532e7b7d378b855ac08363516bd61596fa56c5bdca32e55cb64b5f5daff7626007ba221c6d47e214e6ae761188bc88ffd104cdfc0bb78df662c22d5f5cdc42288ef393fc868c87ffa516027b72a206f7c38813fd47eec7d995d3dc6f55801389d9682efb23a40e7c04efb14a04fccb5cf4c8b0d797dc19c8ff593bac84bc398d229363979b0bcd0362e29af4808051362b2abaeda3d34770ec8cbe6e9de1c8334d920a1198f9913847ee6e4e72d64f00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb4640a0c488b8e5dc993445d2857f4c77ea13279d5f2aa253305ff4a63356e5d0931e7384a81221cb42f3889748c4de6901a94f7c9f0bc1ac52c7b83859721dbbf4e97fb3b2b2200cef6815a5966c860f5129fc7b1430ee27cc255e1c50102be1f762f142fe2911fb6f7b2bd6950caf821b271b729fedf590c22012f3eacc4b02d35f0cbe8f39571a2b3da00d6394ecbdeab9745eda48f2fe3e759d53af5c3107af991bc498a7f4a8063186f2df51501d7587e15e1f2324b2f60a8ae4029681cd4ad0d14629bc571baf9c93b920d103f63058fe9ded2f9b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h55a3333054553be9fc00961acc90f9aaef76175efde202a76099225026e629768ee972c68a4e56721e9510ed5e102b5968b60370b010b0e90f89d52036b01ba01efac8a6d25357f6e85b2078b4e92a94cc67da9390283945da5095142daedc333c94d45baef4f164607d140bc797be99f63e7397cd636114c51a2d0295e055efc81c79e1dc77c44f770481486bd771b125e57b52f7b041f94f5dbd98c169adf347d1f8e53b4723cada7133aa68fb32883268be4907f3c4a394f40cc39783816aa7b8ebd92e8d3d4d7a7ca33ba3820e91c8fff499f2d4ef7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcae8c7246aa73651aff0ad61505c3329d7ce56c44dbfa32d4b1f9075252f1922f2e9358a1231c74e8791a5408776cb5062d3344d39808f9dcbfe1509f8174dab38b1b252ae8dcde4760b5c4de7abef6b5c747ff96fe16b76eaac176486476a752241c9440eb7d6578a4cf555aa0604b9e1438f0923dce63bd3d096ae677a6122a2ceac8b4cc2a9e8fdf9de332f9521fb6800750b088d049c7969c5f00691c4e90dc5217d5b1bda15ec00034f62f1a23ccbd57378f15a7f304c2879199bf3a275f54f10bae8a0bcc2e99b91d99dc6c949f52c1859ec0b8f69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h311d85a6bc20ba6e710ca22305bf50f498272a420f2d2d1bba8c732f4d9dfda1a657c9dbd7f9dcb5285e14371d2f3526bb188afbf6af74f3cdb32351618c2123bd7d4c22c29845decfbf99aab461484f3e554b5d6fdc55e7f975bb4b4400720fa21db305c8502f4ade7a0ee376a756704e55ebacbaa2d812a92e61b1ba1e6962b7e9d2c87ec82f90552c21749b7c0446fa28a13b298c75c8d29aa7599f4c2165530fd9c60f7015d2efa3fc152ec5b1c486f5c6ee7dd5a67efc490caaef035d2696e7f4ce77ca3c2ddba4575cb2f09ff8202b817a9558122e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2a8b8aa8e98eea16ded26d64c5ccce3dd1684c62fa69b61c7e2ff8308b1aa92e9a97af1618a70476b0fbdb7fafc988052e55f2f39b04e91321225ab62c9c86bf1deffd7857049bf3d6113c7a04605399b9d71b4280c66762147bb86282f6a33721405a20a0686bfded89b10bbf25a9ab09bb24b71823005bbca35cc5cd96f9e18b9d09ae3d9ca1c929fd7db20ca7748a663cd0a5c35a2c4e78a4c9da197032669b7538dc9f3b45e316437c83d2f07be3599cbcf2c6502b5558ee69918aa832efd3bef9064df2115d8edcc8786c47a8eea7785ef459caa895;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc0acdc103998a4712462b630d354d5cc12a58851bb7ba121fbe7f856b14d6a0660265a2f7c60432eef7fca81852263e7308649508d21acf89dc2566ad331f23b7272ee6d47b0bae121102f0ebba305abb9359978785949c22ca5fc6c7234ab32c792f131428527ae42652e25287a40f13a556eaa782b1cf77fdcd961c04decc6982ec28b274c92a4dd7795a1d2c3427da2ec1f5902140d8af2290e8477ce75f9132bcc6ebbe49c279422018e14ca97a3ddd57091f2b66592f4f39757e87a6762ab43f88693a714ac2b35e21a433a28859554a37444f1db50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2bbef07760feded212b9533c814726a3e1435de204597aae2376385050cce70b72d1ffd8f70848176678bdbdc4b6af84087043d68d35b8f42a4fa93fda102edc4dbb3d08dd03de86df7d0f1da5a85e89673633900af05ab84f8dcad252a4410578220e6b65dcfdea19432b5546e717bd494c09c32b4910da2d0c20842359e1e3a0a7be58e166b06fa2699e0ab95bcb85f5780ddf75fbb7741fd898199eca7f752063ea01328bcb44069103d56347918fb6659fc8fbf1c7e6e4c5ad24047dd4063635948915be056fd834acc00c8f922dbcfe3a2e03c843f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfafc246ee3789ec468263d26be1d59b9a120a6ea251bf27913b18cc62700928567257954f48be966b0966d3e4f86d6f0db22055e6d1ade6bfcec250d803f5c8d83dd7d41549d11f136a0a1dae44a8c1a40c59920b8e462b684a15ba42f90d092760097667c6b68505806cbdcbd7b9aede328e76ca2d566aac9a7f7e3f3ec2dd30e4d02f71a8ab92acd7830b65b8804f80947a2c36c549b9d21941fc19ea26bc170953f50faee616fd323c201965aa31787192df9c7d0ef7cbd5b3ddea3073476f1c2ccff17e9fe7bdf70ba601e81eccd004b4981c7d76b4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb0b896fd2c80154b3a7db8550d49f3b6ac72d368d249517c6360ddf9d6150fba074eaa3ecbbcf4cc3ddff796d129a3c2bc6663cfeef259f8272297246805157162871bf018b85adb054b3225d7aa62be5930987f776fa265a6def6c4a8afbf9a38f4c1af57c95f589cd2573cb80305ea6223eaf45dac7e6d00ce573aca2421332802dc7776be6cd5b959a2a9e5a1ad5a28fd23407ed7ec09afd9bf0d4327aa343c61d697a63a6b909bb6a6436c57f2ca5976daea2e495080d94e912496ef8647b04f9815aed3a35ab52521c8b2a0262107211b59a17e747e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcba0b15fba69aea319730a349b813efa47f232c4f76cbf2128ce3cedc589892e194a9f2f1f3add081365d843d8be3f728e97999d843064eb4dc664b8d7f6ca0027dc638ef77db788e9543f3f530457c0c77641ab2c50ed7ada96757ee3becbc8b903c8c2f37d18b76715d42e59a1c2b412702843181a025da2d3e0d8ecc50142efce6e8fff0919fe32a4f2d4533340c60cb3b3c7a2e0df36cf319df2b5bc7cba76ac23928ad19defc6eaa57e3f467a605cd259e713c1ef4bd8593a95b43efd5f97bf983a28c1fef707dd7056dd30ac87e4fc9203a995c410;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h87466246b7eae5263fb0e9a13fbcda0c46c106e08f82f9a9a4acaed7f346007a63a83511eee26fa2a4b7c95980ed9e48cdd0f54add2cf5ebd61fa808c682a748f78f571aaa1296769bcaa11138cdabbe59ac2bb6b4b5e2f282399cc48bdd3ac4fbef4570a64e6ecbfcb0a33e2cdf3fc5c6f64ac5ccef9488f9799529628e8c584aa921385ecf473b8bd10e223852cf7aaaebe2e5238cedc6b9d5c6810d09d79ce75166835b4c66aa2b1edfd67eac4b5b5865a4caeb33097dbb431cfb205579af9c373d3d1b6ccdd6f0e030f2abb6e0ed1aec464dc615a04e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h934d1f388e237cbf63d7df0077fae925855ba8abd63f3d1727183f8231bf2e05364c347c4f27566d5da0d94b4760181094a39d9b0b6d718768ab93ddbe7887065d35defffe342c1a34c0bd2f909399254ade8d145be4fbd0254979f5c557507ade3aa2e8e4d7639fa8190d7821004c8761caa38605f70d00786bdd4c5fc987c3d3ac96117466b9634c0cf366ac39cef8e55be4b2901048344183e6445c381abea8bc08dbd68ef37d7f241bdbfd872dd69688ed3fcff3b4bb8116f71f4dded95e7dfe37f111d84a78b576cf42b0ff640db7eb18eb8fc81de6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3911d065abab541a80e45ccb1a5b156c8916535ebb0accbcdd9520c99b9460e54476a9505fcb1ec1b10ef6b68760441b4fcce42be7b793ad6b411dbdaa8e28d0cd153c65509b1ace3c47695eccb1bc931b246fbcab9c126029a1129755c45430b8767c32d90618f6fda842569cc493e35209d572c1fb6003a39df2fb0e0bc8f89aded3f3b458b5ad858634a910d20de5ee498ad10c2cb5b6ea1c077e7bc73e932d811dc587508f99e3df7b895ff0f057c8bc66322e7fc65d0c95ca3352c725512ddb1bfe40297f8d1c40a091b8ef7f99f1e659ed647df1e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h886289191d1cc33c8532ad235e6c76e55640179398657fb7e026c88093e23e4751769dfb59d588327f62b2d681fd5fbc652fd2de2415c22b7adff054069571e19fa3f82ee1f7b95a461b448949aee05aadaafa96a999f7198f07dabe9b9de8b6cdd89aa1d1cd3db0580c9a89108ebe9a1d500212c00ed59f27e20b8c7dfcf0c4699bab34504ec6d45810ce15e83ee156601c2108bdd0a00da313d5fbeff97442a6eb052f44ed7e18e1cc692c46788bf30a7a01e0be229ecc93482cd6061f8c732ef2282bedf74c8d7045af17038ae194abe007d1012072b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha59ad7a2443ee603b433d892979defff80e399cb44fc5c3234be10017fc6a98e7df3827575582fe5075b64cf2c01fe456949a3a7845340fc9dea79b7848cbc618d7e36b13d646017cc7b06ebdde22f2cf4b1846111d314452c6d4380a52a0fb15c69443f6c6f0b66ec2a8256e86a0b023364f9fb89feb78e8289a111c036e58cdfd62b009506d99928cc39510d6e811da6e080a39ef75548eaeb0a53e64d7b9e7d0f8009f528d9e8e91714b3391ea573349b96722dedab417fe08e99e9ba979faca505b3e5ef13a364c3a3aa12422e87277aebd334e009f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hdc85f9e1efa1d42755543af0065ea010dddf5a35cc16e0398d27a7a0a7af2da53aa2c8af7dd166051f819b22cb6896cd8f2ad7a6aa6f9d73a5ce8fd53478548f723c14bfade38352a1d3e4c590069bdf84bf329ada856e77232be80b61733061b56e861c390f2f49ea10628ea16deee2b7138789e9eb02299b92c327728d37de12025ff4dc4684bd966bb96bf71a189c8732360ed1c9552902493c5494b2a8c019f67c091d5767ea503a9fc6ccfe04bac5bbdd41032bf3415b7f54b648df5955d0d6f841312cfe3c8f8d68f5fa6d69d2d37f83ef68fc9bcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfd7c593ba088ebc10a6d3de8b37322001f9ba5df1e2554c18ca3d645396806d8794caaf230f1eeb3c0c88ec0dccb19832a4f3d5718a11cdcba4f681b132c266275da1d86d33b1daab0d5214dae8b96d5e9250c02c2d591df3dbb6946c2a3c1b49e9c37771baf9a8c6c47a4324bbccc90525cb3af80621f227bf7bc71df0208e1dfa1efd8fae0e505ffd901c2af1cf1a724bc01580a8282698fd249ad5c702d4929afd426b1c447b417518fb7b7bc163e35230ef6e3e828e18ea4afeb8d06f7eb5b70093d0b94def0f663a43204ea8b1b3c5b7797b88387a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h57018b3547f02a5fcc86938d8b224746733f7f1a18cdb91070f8918dfdb6fe86a56aaa5310447f39a548f91ae68a206b4c0e6401439dc1e2f404e546e1e2de51ec4749d3a024b8a961423089d40c020b308429e7b72bb4433825ab4aec5d510b06f6d9577f4ef88de92d851b6fb48775186f92cb0a57ea746478c3dd8772ee3d8368a0226878054de8d6146be458da58b1a0771b2bee4e8f49c3057094ace258b1af9c4e67d2af0265a57a6f3994b2ccb9d443ceced814d2e3361b991a882a9b5aa710d6a4c4fd68eb61cbd9d48d5baafcab7e4fcf8eae9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hdf4557a5f852186a810101c3bfe8a5e2908e8a98a0945135c922da3266067800066790552d73e2ecf08a69d133be935301593af08d805c06e9139ca4f83cdf3a368076034befe103820b3fcdbe786437e391f8cadc9a97381358e2829a814921e36a691f25d9040325bb13c23a2fcc7d9456bb113218da74c13da8fdde8e337537dcb4aa00675b840e1a16b0a855873a446907f61ee6584cb75cd9876e43dd40fd5fcdc32b9cf4edffa5f6858e4ad4f2b569febc460fe5bbd0a18d6f75116561aecacd8cdecba2528ba5624f34150555fc7f0bda92b4a40e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6f82a56a3a9bc3f7dad0449e85149704d88ee7f4a0ea7243537ca41abc11fc671126ecfd3db73676eccbc0bdebd2f6ca504755eb4126ef101ea644ec00b5b10156255125279efa700852d43ca9c5a34651c8a7bc9d427244f8b13a682938c8a53b1147de768a876116c953cfb91898cf0c6459517c2bbdba23d0b846b2bb1d6f6fc509c01c99b39eb497729afc55732ae1f216f2e61bd9c52c16288b12781f72f93979c7a6a412565fe25a6f86330788e6b97e21e2c6a239428bf89ad79f5efafe51a9721bd04bb98c1a097d015f6f5e708ec737cf1a83f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf34cc36229f886585504830b704f678bf95e23ef8ae77ad0a12b027318e690342729f668501159c50f1939b7cb4a62cd71ca6673fc9f7534109b503a109e3a3ca6b4d0444edd1a0589bb40ba4aa7c6ce295e618e0112331d9f700b592840ab86d1af9f146d6379d5adb0a9f28cab87b4a3fafc591a489ba291a0be4070cbaf88aac23688d5458e0bfc084668695f6367ec09f1243a88beed30ab4e8242da8bb1bbadbfacc059d9abb51376458b0c63d8e8985be0c52ae5a58190c90c0d4c3a181213cdbb669660862cae0ecb61a41531ffc20ffb15f0e170;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7ac273b4d1310707094f6f19e9dcd1c750c541d64456dc051af3f72709785d40fd2c47e7f33fb1ca65287211d4c25684440e605793168089dbc0837b998c5aa3c162bd2aa99ad5b902907b54193dfda5d04fdf6e06aa5e80e9fcb71fad461db688013d766851afbfd11b18eda67848c06edcdc57b8d277134c3f95f205b05a7d590c761c93ebe624af570c3af6968125b57ad6cda6d01a2b27e4ced82a730e7bd18cd53196a0b3bdddfce4946eda8af35f742bfa670f42069fa892ae41e32ca82ee0ff49371cc6d75cfc6299ba7f29d8d4e8c3823e09dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6c24b8a8a0fe5c67db154496b17631dbe1a8fc6dd617ca6f4ec7c7ed1cf92bec900f4aace2189d862324ddf97f7421f6a8aedc517ee5691800aa32ef860bd385f4223721f637121b15602214cbf11965a5a841cf7f93d0f04ff044ab39e9c466dee11b2e740eb3980c39f415981920816254acacbd32b26f570dd9f553bc0af65a81c6c8534602257909646dc134d25cedd65bba92fba2690eb953231f1dbfb6a90f50bad14697db9ca7f8777610803441d3e2e34733857274d7d57cd6b436e2c5ed10138ae2ec81988f25c5ac6215045dfb758b17989389;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h597d1f80639c532835ea4acdc55e97a4a8975d0fcca3cf5c2fc31d88198ab2d4f4fbee0aae9c3df48e0b1ac076ad989e58af6f5a97dbe1e8db335689b3d6082f8bdb72070c3aea6daa8389980e0005d942e8721609dca51cb5575183cf01e7d0d8f62f4478a290f88962aff6523f67fd4df2dcab192ebf59e6818e53fdf357b8b70447319069db8a61339fb33a78f64ab81dc0a79b5497bbe41f80deb91ec4de171437314d5d4904327e2e038f7355232e052e9ece37fe743bfcb181fe30d7533077a0a4cc969fe290d42f6a8bc7d0c2dc2c8f4badc65705;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'haae9bc9be12f9c6d83b5db06de915418ccbf1418caf3f8b318b9cd81f1569b2f7cb97fd48470b2b9097ef5859e02a96465c1b0b695757134cbba7dcbea85b804cbec91c2fe6d618a0af531494d4d7bbe245db340ac573582b7b994c5a494d5f6ff487c6bd19dab0230d9cd71d1fad2efff41024aef53cbaee191e39deaed267fdd423497a04edb193812eb027f6276256e57dda52da895d7f93ed3910e6fdcc3a0d57659acf5ca179394a46265c94a2dc0f5ccedf2fb8bec2e4eca515fb903b30e4926000a0d25300dbfc13f4a9327a14d30db8f50bb722f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h4ad79d4debf36b10c542de8aadc5641526d27cf41aa10b106408b68d5ab7daeb3bff38158f84601ef629e3f712dd383c60d1d01669fd9e76b8406368f16d0858786d18f6634e5e525b6de8988a1d64d14fabebaa29c331df329a1775e16fa9d1087be63a6253fd4dfc6e43aa9f1c8ffcb1dd1928c63ed7666fa1534deeda67412006119fd142e310749fef9a27cf92f1448467def94f71dc30fd68f5c4da341c38a6409b7404335f45bc7dfc0c6ec0b70db9621c3dd9f044a30e7405bae11975063c77d3722febacff74f51cd02e1270c607776d2b24db41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8ac229b893f094d8fd21063d0fd4bd75aa5a819675379d88ed3f662df5fc9903762fde6c1acacfaf5304fb4d9513d511f688ce2170499cd5a0b9b6a8785897d42bdea5f7031f844921e2d04e380934ec5f5e8d490b393d9ed6169980929ca70c0bba9cea888777b6a1d182f1d700565aab672c83b2215e0ba203cf5e3bb2358076a541736357a263d8cb17f9dd6999b256bdfccf9c4f174ad5fe9ae814db30f8b885d96ec8bca3bfb1ca0d95146961e5eed014651524f2d4cbf481db7115cc68a3c2718f492710fee6209294e65b6c4bc4e378057311b2b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1bd2dbe1724c0926886f0fe43e9fde752788051f0cfb1e5cb1324ac2c305d95901bd813699a4c894d7826dad8938f2251e7cda7d1e5fc46f1e53a641482673dbbff62538ea4e7e9d38d5d6c10a6c85e356c3cc27cc4ef7ba4890641de79fc5ba56c0ace0ad9af50cd96327e208de3bf9c75e006c3ed046f1268271b74b3cdf28c8e4038cc8dc72f99c9c75580d8ec088c3bd0ab68515d6e2a5beccaff92d7707c0412b0233a9b0f753862881108913ebf33a919425784868a798a55c4390b9d82f756abee9bacfbffe73ce257288b4e54e884485bf44fdd6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc34659d73119863ab78202bb8cb9eb1704fbfc41932cedeb656ea6589adfe823778628d082665452ab808e31b36c6b56fe841678aca21e084e530d7a657ba53eddafe273c37c8ea9234a8e105a5f09cdfd78aecfeb9eaf2e7a99f05a35332343642ab942b3cfc1ed6b5a6867984dbbd2506c106ba197c942f6dde7695f7a36496e46f4793e0ff91ee3b2e66f9efa835335f7b0ec5a3917c81de7a7acccd14116aa098d7b8ffe295d9bf084604def87b7efc0e898c6bc22d846088e69d20314124737207d7abc3c041431f998acf85b9cae03a74bfd3c1afb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha38bff43b4dab3256dc53cb090c2c69385743e0e6ca4e09849fd547ee6157910a28902161012379db5fbce536f22e47205ec77b68785bc9bb90a05cb99954c81560810fac56eee41f0299c80887150a9da7883c775e378a01bf9952d2c1f8f32ec977809060c66d13bc8f8733b83364f70990b14ef05ceb686df49941a18fbdd0d6a1f0ec9939848000e16212a84be26809df4c1ef60279114bbbd202f1ee3440c0bdfaa044ceff9bf416c5a782b0c4a389931bdf83de0630cbc8eb136e01ed587f891bc097c3b17c46007f822ea4b6b18ed223b9cd98872;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hffe04bfcf7365eb1a5f9dfd5231c7bfffdebb1b36dc0289a73257a843994dcd850db8ffae73dd63377606bfd24331cb80f6003998706a87d13e2c929053d39f76ac378d2e6641cea3d9e0e5d5e37d24933c068dbe8d0afca9cf09f4af4fd0988deb6ce0466375bce8f1c410fe88607aba117e991006d8ea494a80891ada95c40f487d14bca4efc58e70a1cb6c3fa2fa4702317d0fe288b40c90c8810a5c9fd68434703e7f75fca3e63736a782f32d012031ddf2035e33181e460f99fa4646cdca261c8e40400fa8e479200322a7a3db25dc35dccfa8d7942;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h715646683ada92a9d8ea3ccac9f90544b31e5f1d9183fae8b59e9e4685287926bb1c763bd6f8481bebd50a8017aece5546051b6ff4eabbd854171992e77f44e55acd66988f92edc922334961b0943ca3f59d872d99a3ae06f7b0c342050dbe860e2f19103bd41a77fd1b7953f79498de33e0a79c8053eb1d7e632dffe8dac522c8b6af8e9c570109d779940bf24ca294494dd2ca3bddd23c014b05ad16abf848ce1a297cf0eda76b52713c5ad6f07a029432bca9df4a4a6684775b826ddae87197dc32835c35ed5b3138b16198efa0d022b03dc148e6e6c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6d5fbdaa4deb91357a2dd66a16831010b79c36174a72fc7c0e543f85e4c29bccd4f8ff325cb281d49b9a08247a1d9da0fc64729cf039cb76ec62f05fec29e3403a3359783bf51baca0c5032302e9341f7cec84b90b0adee1f2b67f94bea3f5892519a8ae50fb8d1255c783a426fc2b6dc8969a09e0cd89303d909951f9ec2f213004f93f9f9a55303c097a1fc15867c154c1fbb995ca0280bb51d5a3a1b7d332a61b82c40a2efdbbe23ddcc68eb101252c04ae18a31b1124fdfc82aae8b29586a38f61c7c7c84370cf03f64560f48022249aacb4a2249c47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5ba0df6f59019fb441b6dab2b638a21d8a30e2f80310727e444371e1f2f7c315a13afefcebb0a7e4dec4bca36caf75e51b45b01142d81fe78ad10785bd0d5dc00152a2ba13c85edbd6147ffbac576ec5508c82cb1d81588bbb1da65fdcbc39a1a516caf3f46cc0e70b00c81a38249bcdf5be1ca0f44e645f6fa09d9917e83b78f73fdcb1bff8bf7b97c5fbc38932dc6f444bd3b9742305f764ad399a11f178bcf9526bfefdbfc64f5fbb34f6b2070f85ecd70b9e1d525aa7311c1fa67a6a3c622264e1aa9f6f571b54c4606dc0fe422aace0ea6af57d94d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha3ff580a4ab35dc3e562853d978969ddfc47d5f7a9f156f728cbf8f900ccc906a941d0b3e7bdac0a6d9f43701821d1dd568b934c2ddd7ddc47a1cba006d2c0f0ed044e9107f3143175c28dc8c3ebc5da5ee7c3b930b701502683f52c3533cfd33d1ffa4ee2af9a44d1335c2f10905ea92bdab5340092a439ccfa499f0eb4396375c521009c9d3dbeb0856116989dd76615492a41a9d7a67e1187a11d7e04f593decdb90f2e927cf836e109beaba09c4468a1118f89a90ad91672455feb8d94d28834014cc60870f54b8647fc45b0543f8ef4a96d9d2add88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6f2cc1efc1a08789b5b09e88d799781835802bce746891c94202f747bc836d384666cd533eefed8bcfc0aec0ac643355196d0a132be6967c84bb65ef2fe88a3d9f732ac36b1da2f241fceb399c3d06f8800dbd09167c8598f0c1a32802531c59bd20d08f07a279b6a74db7124e77eed0ba33f3e0622aaad75d28925d55117951b7f9724e6a0cefc8d05e8a7e22fcad05373a1d3665af5cc3356e5ddf8803528c6e18f1223e69b09f9854af0ce01ea75367897cf4c628534998217068e6bb65472cba299615d463d7504f81485a8131c2a67dc4b49bb6765b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha28f328a7f834ee20390e5cc5b7ab4cfdaf2a562a43cd06bfc44be21958b5d29c51f2b888a9d21a95c15644849731dc9e508ace9c7942bdda2a58c999c5435d28551060374850923160e5c91bc55edfb1a16add17a9fc8cf2b8bfdf1bcbe960516a84cef48bf1141449a41d2a1e32a7fafbf96d33a4e93fe00de3d737c0a64e7090eed4c33e0cacf47227bf729cab973450144fdf9f68171437a230036e63b2b4e6e48871c589b7bf1dc79a057acdb280874678ee55093fec8efee0e403833a382fffa65f5594bcdd78db848aa8825fc44d95d3007102dc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he6c91c14df614d64b798d8e9911c873db12ec64905eb6ec6b3e8bcdfaa8e32fb77889b11d98e53b14e9fcbd9f142c68f34b1a6be40b0164266a2aa974b561d7aff7b1d1f7501844e07cfde856cad0135108fa085abc52c7fcf4000dc52908dda0408448fe0dbbad3cd6e9e803debe56ca20830c2bdc5effd7cbe6e7808ffc54317923f5d9086871a095f787fe4915d458991ae04f8aeb403d5fc992b0c612272e6eeb79b29cec7bbc7d98927615dd42f2cc74e697676ca458362ea98928cb9ac2c09f406c0ca966ed1930d67a343b8f68269ec99a63c2983;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h55ce462179943abc926457abaa6d0d2b45d28969a6f39413bea339400d24d44b1f3c0a1cb91a01271c7b3cdc58c4d59bb23643eac80228e6be8621d971caf8c7e41fabf418538417c0cb15fd54f118f5f7f4cf757f393e10948b448ed83124bfb86aaab88522da09248523e99c91509fbae1a83a593799f8b6024681607ff3cc48f54eba5b4d86d342c823af1b319803bfb931fd63dffd1b02a744a425416f4f0217db28f84bca77d590156618820412db6717947495fe5a09bb72523484d5adc60ba5decad5022c34181b2ba1d58b426466e8775522ef5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h4623aa2633ca2cb2ffd4c529776d88151bf74866d17f63fcc180f0219e29498a3f77dd19325aea9d41cea4f45fe0bc3377d59cf11fdfa077bc7a7c41def8ebe1f37d70f1eeea7ff78d876a7ae3f158985fa0e0d312a45fb419d185d41b701a6387cd3d4c9671e53aaf090e5278cb26c87d300279293e02f469dbdc2d31946103bee468629430c15470b715972aaac4cda39dd2fb0511bdace1deb7779c7b2d8a695345101c53284040fc44885b85cd49ede2985dab8b64c19112bb1e86fb353e995640bb40d8fe07d2f1998486da3851e2177f3b3397bfe8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h707da72311aa6e9f8916a8256bfeb5a0b11ef7bfaf53510f8667fa485f0c7c48d45f50f06ac99ab73b4b987c40e3b9049b5dcb01afcb31716515871d2bb84e45d5d1cc2539d4068768b2af49e4540f9c7b05d6455268e8148da8139f7fcf65d2761b6d133a71e6e5a3d667e3b16b36cfb83499de22b4f853b40eecc423b416ee95a049fd3e79619fafed649e254a84302bde256b5bfe45907e14e85c44892b9e5236d64d807b3bca30ab228fdafbe2f7bcbc745508d9d718dafa5e7e8a12c83de47aecab772ed2727081c9b3d319edae122c2517a183fd38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h85ea88fc9749cadc2932dbc65be90b4f418898fd3157629c1b55b87d6cb51cde0bdb121e8f67d25aae4597b3ee584b532fd6d6307e6677833613d51286a556f592fb16f7ab99e5a2c113c4bc16d299df6265978abf635afee0762cced0b018edea038b3749602409282a27e8c68e9c2e5e8c9b97e4053a6b6f01b8fc3364a0327ea04ae36afc87a5b6c232b0081d88b02478e8c66df5d9f5611e15ef1a16b24eb677af112d78864f320ddbdc15d97a3f528c08c5f746bdf370a4674c3b85169b7d3ecf2d27755ffa4b0636c87a43f7812cad1d709cd81ed2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h621993b4cb90bd1a58db8406e761f3f3c4d0c49cdce6756b2f33d1845c0135bdb76924a125b28c0be642556a3cc6dd144212e9d7e3444e0426e27994c4e3ed9caa25232877b45e51bb5bbfaf88b86e94a55d0ed64985ab16861a143fb7ec2861261cb7c26f5bb8fb61223a47e15ed944331443268037bb46b9e7c4ffecac942623287174b7e50047fc0215dd47b9606ae66eca7fcbee8c04b623ccf8e6910ded4ef28ab9e6cbe7d1e1c45544b19a30538dac384d79754aeddbc5cf4be11c79944f2ef65c4325836af7ce5740942ad7a7cd99edc0ae9c661e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8fadd707477f69bc62783f8a0c22a1ef5f31c429de000f5ec8b1d1469bca56f56e4539562baaa16f3e24be0584775fa74a9a8e9a806c58f24be1d9c2eb87282d4dfaab9b5d04174344c97c02b3b1e6ad7c8957448da0a018fb3f51f2788c5d54dd330ea4f5962e7ea27c1873dbb402492eaaf817a5ebd515a2a203c2d9f293f882fbddcae4433dc3a1305308d2e8272ca51747bc87c0b63e93aa841bd63ca675f692dd16379fd0fe2a1eefd15a574a889af668c973da67d5e7e331148b182b1bcf915c782c20e2a8821e40bd0e886e8bf9eb6f6b63e1de0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9c42f1db503ca91f7bfa4b18dcbc52b5515df76b907708979b9469842d8b4d0dfbc7ba69d1f96decb93b606bb4b17af610b87d0598245f76a90cc08a14357b23849943d89a466fc43fc40016208e59b3332b7a306eb393b6e614a1f51a866559d8b08a4d4ab3dcd13ba0c3a96980fd993b0d95b2b6eb5ab0ffd0603f255b944ba49a48c615aa40cce144840644fffd5090d5a882238ee2c29809f09c8aacbfd00bb1332a1b5c3cfc8054bd057551eae45ac46ad5144aaf220bd7fffc9b1ce2aa08df25e5a10f655ce6abfff40cbba8b05376f3510ce27c9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h43a5a521405d5d39e46ee6027fde0112486eef11966e3c281f530c48f468e8f7c1dc450685f1e3bec900346d0ff03642e5d73d3c3230e8681493b457be56d3521b859f34b4dcc3b93c1d322f2f48be6dbc5fc1b09163b51047d85d8cfafb5e2fd78e512081388f39e89c84d8357d0db3001eff90c845fc8ef85597562e41955f9d0d6fc989a8b43c91b9baf72312de9d986a0d2f4051a926fa5756b60e5442640a8c6f91f992d26939cfa8afba9fd37fa04c4de7a95675e0bfdfd6146876eb46b36b556cd0665cf9d7456be473886da58ac234a29fa6bb59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8a065312afb6a4ba8b3668ccc23545885c0d471b06575034ca5fcd8cf5ea1d3fc2edb0cca95c9e0ec08678a83aa70c3acad1f50fca18a1fab97b7d8574a2921567b1e9abac9696b8bbb3b58f52d620b6af349a6b395d0c24b3c89744c92b2437768a5cd9e4f6a0c4accc7145656ed7b04364e135e1fbb74300e76aac51ae02febd09737355c36428a2632163fd3caddcd1e3d340850ee970e1b047359fad47c54cf36c3692daa0e904df7a7064d45a42e622f05f93441b3fda2f1ae867dbb592441fe0cef72b1162860fb55739daf0fe04bd5c6c66e58ef0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he9ee5f074ecf656a3c1d6c5c2cc23e9a85764cd3b510a1b9c29eab4053af572d6785427453e774f3dd009ad56b8bde54225010f8c5c67f183ca910fb6d0c3fd3fd00997018cac27db11b17f827f9649f691164f72b4e6898d7fe5ce68f29a5be44327df8681176820ad2ab87481df9dc8f1588c0896696a06faa7d8146bd9785d1b2a49ed3c051d62deae3a7d30caffdb0689a2e45ee25e75d8816d48ca0338142fe9e2a4ed2e18264f8102ab1b380db014c88471a2bf54a75f22d130db0fc1b9f3520269d927fca6263d06636a165495dfe3a12bae612a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3c7b811531be4f30ca327121da8f658233f609ee5ee2eae75570b91b6b9f3e1854aea23563cf8835eef8146a2e8fb679a579a9d91868ee708a2729d96b009f2eae1269b256c08b3ae3991281ac40fb37012acc82f97e6a402fd7ff6f98a41e9d4c78cee03726d3e495febebf25ed3da5e14bcc0ef3156c924a864d0c70d2a1f33aea407fb6a331f53f9a217081867133a9ea641016c71f620df164ec4449a031a957c3aab7051fdca2fbf8dbdaef87ddf31fee534d995d74102894566352339839d3974bb30527c1e52e7df006783fb7a53c2349d5571af2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h77beead5e1b7692510fe62fc1bb50a03d52aa76019d2785512fb24b5f2b59baaeedbfaa8604baa6bd1a55a5e5af29067d95e5abc7074546816b536b9dfe470f619185555f5585d29a8a7465d6aeaf13623b84f8d01d2d45ce33b74bc29b26ebfa0cf208a4ce8a0928dc2d70c827c4e1afb3fe0e5ed9af97b0ba4017e8d52a3f3a9b9035e037afe5d6f5d2f32ea178c448df382ba92fd4ca1fffc7a387834f36ec16b0cb7d121a765908bdba8d84cdcf0b99799bd13ab99f3381a5f526646d8a2178c881bc2ce8046ffdb457a1cf3bbf2af4295661abafe6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha2edf6dc9454476b3a47f6adc004026d6c9f7c23d8ed3f8ec24b3c0ceeaf88ff380faa9ba0668c34ac08811689101a9d6144500a854ade58d9b4c1c8ad8d9c1981b8a1310779b06b9a8c86fb7947bff63ebc77498896364d7e0fc644a6e7fcd810289ee6acd93bf4f3471ab6972a8b44c25309f92ad6c038df28ffd734eb767a5b9a9b58921993ad6974e4880b460c4f00af55a1dbe2b83c900e506e127e84922c1f38d7e6b3b247ec3dd0ef129a6870b5558f62fe4918a093e0e56518aaadebb22c09a55a206838621580bd4cbdc2da8c135c91ecbfae0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8439431c185bf48d88d553a1b3fb5108abcb0169d2404b9e671b63531931bccfb08a7a06cfb2fe2b8891dabb80ced1586aaf09f824a4ac97be11df91ac7df59552dd1a8fe01547002b9a127fcee67f1cb4b286fb8b934969076cd461b506d91a0bae8bb9e7a2a885754aad981d672d5d2e39801834bf2e64622e4cf9ba73baff1414cb02ee7c2636a256d047e76ab79d488518cf252bb3c57af31e53b64346ddd6aa3b4bfe35fad18d8e2fe62290f1b227b792c262ce34d05a051b95d246842a9f39ef51aacbffba9d3e40d61f01fdfc661b71ba3f94b788;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h291a05b442397c6b5be63f24cf6376be4ae206c139307e28daba1a2467e4f950764cf3a279b06fe1f5ae4398134763df942ad9a54bc8b72f0011e9d17286f0fe88d10e526674dd461c78fca6a12bd05999b9478639be3c6e381cd24976be3e32264084d9cf33a1b08c25dac2b41066e80aaf221d2ec3ce6ce7bc2bc49ddc99cc544e547d6c5a9ffa00211b3580c497502810df5dbeafa96853f8bac3ad6c038e16081918568a6e082a235891ba33e92ee96dd95380cdf4a00a567d5903c4bc921570ef00413315e472b5189fa115cfa33c0088cc72845d48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7226c5f4d57cc1afd0aa5068751eb43ac6c974da660b72b5768530e751963230a2ad9e16d5e9ce080f37432465e4712a90477b81db164339b5b733bf7ad3ad79da3550be259eb6f38eaa3dd6256cd4dcdc6ba431865a99439fb258d6a18cf4e7a95bf549898b13a580c9734dccc09599187dc4a2df20863780439c7351c176b7a7778891f4bb083270037e37295f24a86a2252f9cfb4d32b25e48b5294df1c373ca81e90813ae66f7d8a00ba101a991e27f213351d7d9c4c9dd21a89517657778bdb470a1c18312ad4e0331ead034b829f6ebc3121819ea4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8d331e53e2a50146acfe059322c1b347039475109c747777afc7ff7c639cb271460a5e54f18b31fef19ac4724714d4670b51151fad4847d106df68bda86a33c6dd6e798fcf4a367ddd237d4facbea98f4590f82789f84b8a1cdf1efcf037b10368c09f538e9e48781ef43e7afbb28a6a60c1d8407a577e280ae9cfaa1eb74a33c7bb698ee76eb252cca15490ab0fc5afc57d3cc865717a84b0cbf1996b3a50f14a53425633b69b3e19c01282ffec093f8712622ed0ab2f80ac952cb018604f64dc1f331f14073455faf565fa74dd86d8706bde4f7135975c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfeecdc7799e5702f26d24cba6fa89ab5edee7d38a32965cb67d71dc2317daef38b4fb0af1d4217139ef793f1bcc039ca47f83c1247e66fb97715aa80cd0b8aace6ddb7415c1a2a654d838cba99f4384dbfac9255d46cfe4c28d7d51dfe40900b88908fb075a91c2b3d78f7fe560358860563af642a1017a31494665a010c3ec38b572b670ce34d5857048d4b0cabb554d063a43c564d94af847c81b8704e043e05a31fc5b9f7e4d84a123e819255945812d73d678063d7536c073f17946faeb0be98eac1d92cfda7a2d2bfaa24cef1abeaf22f6e408c87a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hab3144cfc979a54126e8199bda4a228ffcfe50738cab606f78cd911deee3868c77bd7d5f29451873ab7747e0f1c7e198a7a75fd5c2388a507199d9ece36b5a671238695edd9a91f5dd2597339e6bcdfcf2e62728f250fdce632552b94b4e8a96a0bd3db4c2f536c54777fe99a50c753b23187c056e72a5b3adf6288b5975f46b5724d16fc70f3e3bea304af0caba5ee845a0d128195e4580b649e39bf05bc3b1e4630d6c7e829daa45150a8c9cf6ce4eb9e5592cd73f6ace9ee7a6c28bb83ad42485d2d7a0233adbc3e4dad7d85fe1eeed557e462ffb64cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcd6d9f62226107749c2962ea6562dcac25fe052424f85d31d6045a26503951dc11235cb049a17b0db52afd08181fb12a656cd646652f0881d39f3398a8877760c8aa859ceb0bac7ed75ce14fb8266bcd7382e580a1d1c94c5c0e388e44484bb54e54e363019c2c293a678ea94102a207196c9b169b7c1c49a3087bf00f8fdd08c0efdad44585aa5080b6d64d6759ebcad561f53f53e68ebd03bf3452b9d68cf73f9f844037eb8b1c87d15f2ef2bf1ff5bbfd22f2dd5dbc8fd8b96e4bdf62632852de0ee69cf4bc0cd680c9eb3f41c0c46d302d56cb5fed0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6b4f3ae0de4f4efecbfb05d24b3ce035dedf3da89ea86f7b482df80e1884aa74a70cd35538aaf6a4192a1df3b5eac6ad971daa9fe7b9567ebd33aaf1e3018e4e64e3720695b9440aba8082b1e3faa4b8da3c567ea44fa492cb65bcf5d9d94d8f065651f81630bf4c5c12348fe22c3225e5be3c22e5fc49c431c8e7cc69a4cb205a885e00b8c3208e6bb5b5edb7fe2c33ac4d9d3daf355ab9ca2dabb329851473b2bd029504e0fc6ba2682cb19ae3e46773d2fe565ad27d2a1fa9873a492e288a34cf3b5f1ff74f2a976bf263298d30d5899139c829e00de9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7cd10df023560d86237b17d427057045c77d76f2ab210a6ae91ff6bf7fd1aab24923353ebc24f3802211b03ba7a8841ae8f4bdada81ecbc34a8e7a96703af8e263e5bbc699c0c56600223bce5bb8d6db24a7897e1544223b2fae4c3288ed3d6364a09cabe343011643684583583b54c44927e03510c1caa0ffac208d57a883b2b14308e976b321578258826faf303991e9ae0fa4161918d40af714a7380bd300088557ecc95cd15ed009027c126e533288680b3ef8862a2a099e7843cc3912e0d112cb6f4a1865874625102467811f1f5ecab10ad227bb7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7a82e8045fc8752377712d0df11651c9688274f5ff8c0f1c3c0a84f4ba5f52e09781516cafc914a2d503c052211228981e2ec2d9c14e3216f5e86dcb8af79ff3ba0399ab2d2b0e20b0f5292509f42797523f69292fc59c82d47ab435ca15a292553f45cc0d1ace4cf1d55e1b64f197699f123af8bfeea17be907aaaa7cc3ad6ec3f8e174c1d265caf04dfd7feead4dc37c4654bff4e6466378b776b05f226916b1979c0cd75fc1572af9331988e621a8c9933163b42e5d3bd6b50f349a12299d9a05fb960d56b83efef36b77f43577364bcf706d1607b08d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7f658198208435e9da1f9a7fbadc47d99c2913387495dffa7194c815503a540eaac9621e985ba0c49081e6db836bd81ca1c7605c3b2a66ab14ec1085dab5e20233edd449b17f81f383c6c6177bbe706c945eb24b7ac1c1cae61289eb33c49a77882cae01f9363d972b2adf6123fde2db87d4e1c9c62d5a0181e99bcccdfcf592a50490c3dfd9181736538370e712ea77679fbd302351fcf2d4a2176829b570db651c0b19b6678c05f2e5aac61d4b6434195e8af1b5402be418325652789033a2d78a45918f36567564a632f7cd686c1e9d5bd4ad922d4be5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8be2de9e40d6072ba0a9a4167bb1b79db69285938033b6e914ba689de57e9fd2d8501b1edd35a154c909337185b4fb38628082bc97c3a09950a8872206041227b7dafc5f67290c90daaf244be5f81a9e52834cf85567640c56418873fb178838069c5dd8d429ff025e67637eab65cc20cf4b2a4c2317390de7a1464da4d8bbb2cb58b191605aa945d979bf6eaab08792c0be3a8bbe51f988c16d505a1fec67dcef70570d00f2f4867a00b98000b65bb2348f025e8d00cc1ef4f115e23da8fea2f143b38e8684a7eff2bf86c855df9a4c396dbe81b2017c06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h273fb96060ea05e0ac02fc0e152e93ec89b1c1919aba5699c718323b79c973cc63acc33bf0a315752d21d0dbd7cf91bfa609bb4562db72020e8c3e72352fed599065a29e2a6946d0792e1d1f03835750549d486981ca5ba455a869cac80ceb5fab9f652e8d0dba046c95f467f7fd9831c6f80345cb3349bdb77c7ae8824c082052992adf412ca433280f0240a388f5cc66af08e80b29ec9ab479095c8f26848f681330008fe9bb2885b50bc0b288d702f5f9eb210a7eb802d52d07e3655775966af87899312d4555c438310757dcd5942f84e1b9840b9ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h115618fe6a695893b4e194c19af612b89637ff88cd51047cb5ff01c5f6b8bbe41c32c2e0cb625736aa59a51c3dab5507d194866e86145c72727f609e9a48b6329c2ef35986cfec6ebf68d0a72e00c2304c21ce0cae75d97843fff144a236c456b77cc1d253df19a747f3f73dff1df85f7508fe05d668ce4bf1d3483ae232def0ce23c2415ea20115a2a216355a0d15cf103e93148e8c0fb1b1b277e38e1e16a7102e14e82bb3305f5e6ba736c51dced68ada6badcdf8c19c85dc5989c83b906224f87c658e50f140138336c6da806412adb4b2a0cd3ef0ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8b6764182084bb1eddedaa81840ec6afa0824d5dd3e6b4bbc437863a56fb4c14978a2e9ca35035a17e5e9d194c808909c627e91e1250af9ad94c2640b5f2cff8639e6c4ec364641a23daa44c958932747b166b0ec1f771b84b395ea68029082544c9f82d52782e9ab0d04b2927cfcfb8bb0dbdb369b5d2fb3f441754845748554acabfe621ff9199e84720d28b3764f14957465c5afca51bbb3bd12f50123b0526e568c5b16cd603be714cb34c827d055faafbbb20a4e038e29735e421ce48e75047aa7bbcbb5403c4e54e0911c0e2808c6f38a72a3b304e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf6e4a9420ae918aab198d7d72835b60e5324261f2c23825f833cb0af75644f92dcc2cc4191ade04ec85f7dd8a6cafb377fce085ef7f4d98cec5a6276575d4ccf04d5c836c82d014b1e8be8c8566161c70c47e625b73c81fcdfcb4b1f2ae1721dd9c9bd8e5b1862bfbf790cc8826e9eac420f80c15d25d6c51a9f82d6850dc1e5dca2a31011e499547813e83ed664366eeab982921a049cfab207f426d5f2117e64075c35b417755b1bb45a1b52bf923ecc742cfc7024808d07df71d54c99e3f380b2639933ff01ee5fc65b94c52342c2206b5b22abeec098;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8a9d415aabc836399578d3bbe2b11b67323ef2ccac276ccd4bc8e55a81631cb5a2d2cfe1a3a60c6bb7ec255fe383be41a7b089c0c41c8e340c3bc820889f18834f12ca10bcaac67f342a4db6712bd0e5f4c24b5637db4363dc51cd24de91978c2d2a7e178dd21cb79ea9be2b89a5bd735f3474515f03f4ecc1986f41c4f43e2696337939855466bd05c3794be786b54b344b8ece27366cc41c9b4a67cdd0b395be5362664137c6abaf50db2b03b1b66209d16066529409302cdce869d1f22a958801b8a26a62472af737d98f9440094c68e2acfd9ad1d6f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5fe28ae4357f4cfa34f6cd2927f2d093cc0d3883e8fd674756343e13491e5487bea9c1873c1b06695826532477f2e6fcaaf10f1ace145498fd0f816236596c83bea7b74693267c548ec85b9ed78e02cbe6a2c1aad56ebba67074661fba064dd1b18a70e3385f487fde8001261e902e2957e7cbb8e10370601af0639a0d06b6756701872bbc9961e564f05766b8e13868b2c3023012d46b94f411445ad79fa0f186418a0877424bf64b9d105836b82ff9c2499409c45d3badeae9e0832612270e9b66757fd35d9a942faeb6acbc9381c8e2d82c40efb7d86a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7cdc38be8ab156b7f7d9df3b8b0445ff0f1dd5369cc9a0b057928208c52b173f325917f88ce6a7c2ad13a28950d7511348a9b6fa5339560dc8ea4b79f17d5cab697b65920b269fcdf0c92f479f64a15be2db9a116d797b020ec1ae1cebfb65f3d6efef191718ba2d19288ccd33ea7035811620d4470610ac440ba19a70d99e25468376f6aefb830ec26e76aee54c370651180d30313f6dd7e3c40e4e83d9c96e30bc8ebfe6118fd244296f7880df6f35faf9a63cc1729b52d157479c37b726dd921daf6ad0d98d9b5d813eb5b53fa6661518e92e7b6389f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfee6df823fc812bb50edd03669b02f94eea8fc8107b2336de590a9bd296086f05761c36c6c02edcc28a32862671c382c8575694db478b68e3538b26cf03648f07a65b1cd755e52738a0f9647120be427a2cc90f81c8d5f798c212ffec1e2d6005eab95f4f17c490a3a0cc4a8a7542cbdd7301daee92ea6c8b1764ad5b47d83de7083ffcf1c7d951e5032a0fdbf5391213621fcd9ac8e0a94cc2c8db4b04fc33c59e42aa15110c04df799107b396475b6d59774e94e23d129f56ee5ec9d3c0a7d8e49458cc2e65445067d67d1dc58a81be9a214766ffa090c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h11783d948dcb22e083a098dbc4a75d58a44fdaeb1cab81c197dd1c10ca946b66ad504ed7016e13bc2ee911229824641cf0edd3b4c6b845e9d8dd5e27236dc3fd27f9fcd583d722f70b79d98016edfe48d0556382fde25c7349a3463f3c0acd726bfaba6fb8b5957fcb9bd0e474de94b7f8d9cd7697ad07a6dfa82d9af67f61d7d4ddd40e24a867de049faee286922f1d09a81be8b6e4808b53a5c8ed53547b195904fa5643b43912c7cb52a5589963bc1c4a1f299e6e0f6f5946e32b3062d0da9dbd1d7b7d9d77bded85ddd8877999a1c3561813a0bd4ea3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hbe424f917d0f150012fa3068e9c71a441b71cc606c15f9c882d53539c9b7fdf5dab06a7b82d7f6f8d55716d5801c2965605c0846f54bf8dc1c84449e1f2b25d8398365d3f5048fc7a5f5498102e5f978a6c7ec77e46bea87639109749b2f9b4ec310c405f16f9cd0b7f66187ed80870b57ce883fcdb04753cc2c74af56da8c0a52346c8f241054bc04637eef22e00c82aaeb94d2af1e33ac1ebfaffc87bbc84870b9cdcd3d44b7c6d3624eaf29479f3ff11432cf1bce156a1b8fd97de0359145ba0d4190f253d6e8bbed9a9366365278d85b4ef8c03651c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hcdf1b35c7c0de1c1c6412c07add5d4d62f74ada8d1d7c0b0266a7d650726e6ccbf03e25dfb2e0eb950d2d3f9dbc167f5fb0b3d1bf23382c7a0ac91ab5eaec9033c0b0e2cacdee5af1781943e7f4be03b7f6cdaf6632f4dcad075a584a685ab158ef6b5c50889a765304ce7401359c3aaac7a7dda5f6738c48d212faf625d31a5f97ba126c382cb35104e23d4417b50f712b3d23e3ad9141e9418ce6c45c217266c7bca7756ddbda981d4f97114632a17f027eff79ab94ebdaf8271ab2b75f62630a91a207c7c339f723d3b83c3a1a62c8682c1f74a4d33ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2655384e2d841e4128cfeca03f50ac4568a4a616041c14ca9de401add2df92ac4cbcd4a49ad5b38f7cb897670124acaaccbf41fc80f0300f7bf61340c15373ce4f27f49ef937633739e07e2d65a69189b1256277b95e403df9ccb5fbb41ea9eca4cbf8889f1f3282176255b42e2e2dad501a4a48134bc7243de175633767840c7fc13bd73622c1d4d6be9479f0ace978167b34d59c37347fceb8c0d981ea52e8318df98227efd23c3b60754c17e541033df3a5ffc67c99b3db57298d065bb2ccfd60b27269c45961f45e03ddf3c50e91f6bb3ede871aeee8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb6b222924065cc371d64d507e6c4989cceabe9ec70d90c8286848177a8db0970965be1265cbeca3a1bc5b1ba30b2bab8b0e6348b67c6044c394474cc53bdf3e548737cc76b68151d70d531f643250dbbf43aa6411da77852dca714679b395f11029dc334ebe5d620d0303b57dbe34540dcf213337500d9f4c16e9ea2c9a6217bfbcc841e92461201f01f1da6c153939054fc5db2590f6e1c21dc736e16616022130d6328c27921667e3fa755c33925f311444cf208c2c3446ff941e50395a5b49dee7c5ef29de7d2fa6a7dafd4c069c48be7c31fe6cf2ce6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5ad5d8888583415f454a8fbe4630864cb78dd8c5307747dde3b0aaaaa75452420384975b5729996a33a34bf09753720686cae3a83e4599b6b945d387c70547aaa1473bd0ef519733ac1d24c232ab2cdbeecfe5e916a99806cad661b70be8a96e91b6803a37b40ac49a6babf002ac31b4fdaff7dd549fc6d1452389bfc023207612fda4ab74dbc7fc4cdc585294d8425d8f2e6c292a5ab0553229114794df15846b2d14cb1e4097addfd794c35705c0cdb0909d88e80bd7908cd0367c47574da925d2c7e4c85a092ace3476d4ae35600773a1a00e7b20f28d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd3f52c9094989d12fc90c10e276b52cceee2b3ccd0a9a0224fdcc0232b4fc6f701b0326f4a6ac470ce73a638a3b10d068ef75ac7381e4e0632dc733d8893599b131dedd02773bf15b6cd19b0deb76087f5235f333739ce6a0b030fbde9389b62921445ea952bd34ba00b5a900a3d61b52a30d5d0b567323cb0fbd8a55cc0503fa76d2c665a8edb5a7fa0e250df779a0a36cbfaef8c75f734b2415e461a197fb5b894b796b470910443b13294cae909b1a7936afe6ae56dc9663fd2eacb92267adabd0ded748512f55ad1864f293ddc39ad514df7f9888569;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc754e43119a707b834047f217c37c4338d49799670b6b88dea4767687f97a850f26db0bf9a8fe3b1fdef58501af6f3dc88ae9918a2fa8ea214dbf1ad2c13de19a4b310230f3db5ecabe93fbd94fed2ee1a0a8699286e68d206ad3be345d94668987934fac437ced71984d406ba306b59b372eaff70514bb1228fb65c2d71861e4098137e2b67924cbf7c3e44de026605d7f276bbe0de69b494c2686a6a3f62f0e8504ea850d1d6df6b6c2be62f8c4282eb9de11ea232275e24373538937b94564f80a340c5b704f3be23ad4f7a8592693952dd40b9c4d20b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha39f5973432e9b9f8861db6dc8fa86485064215f19da812306e802af763f0b38ea559ce5b6eec168bc95aac16bfb95aab3c7901c9f1dead5568b335dc632348c8476ae939c4195167972c48066cc423b3b4fc783852e393519a7baf9ee8771a241b075c33e8e3e6c31bfb86b2d37f225d12739480f9b33003235cc95d1abe9caf18f08c66788ab6da6e36220239ec6301782b3c0a64ceb0e51f0593e93133a319c40575934adce54fb9050dcb3ec8856cf1e48c2b954de443c5da0391fd840f2bfb2ac79353318d1aabcf05c7f370f457daf52527e48d8b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9cfd346d11a738d7337a09bee5a20e5be999d8f7ab9da98494acd9e7eef72ab73091c45720dece1c5ec0336edaa62161466c18c4e064772e3978063ac753305545d6d6fe1b5949f325a536eb04baf16c3f345040ec2212d71db554d0e0a8bdb3e28b06ea2e905cb58f58e2b7911192dcf30e3c4aab882938a8321f038b8ab638bdc0d27000fbbae4c3954114648e3cf03f2fa0be4453d8f2948071a981504fa22e700ff1fd1f9b836026926581031384e3e0f2ba3fc23e65a5ffaa55472360bd0f51a43dbdfb2e604029aeb9aacd5a9eefce7a46711691;
        #1
        $finish();
    end
endmodule
